magic
tech sky130A
magscale 1 2
timestamp 1669428148
<< metal1 >>
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 201494 702992 201500 703044
rect 201552 703032 201558 703044
rect 202782 703032 202788 703044
rect 201552 703004 202788 703032
rect 201552 702992 201558 703004
rect 202782 702992 202788 703004
rect 202840 702992 202846 703044
rect 413278 700408 413284 700460
rect 413336 700448 413342 700460
rect 429838 700448 429844 700460
rect 413336 700420 429844 700448
rect 413336 700408 413342 700420
rect 429838 700408 429844 700420
rect 429896 700408 429902 700460
rect 410518 700340 410524 700392
rect 410576 700380 410582 700392
rect 494790 700380 494796 700392
rect 410576 700352 494796 700380
rect 410576 700340 410582 700352
rect 494790 700340 494796 700352
rect 494848 700340 494854 700392
rect 409138 700272 409144 700324
rect 409196 700312 409202 700324
rect 559650 700312 559656 700324
rect 409196 700284 559656 700312
rect 409196 700272 409202 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 348786 699796 348792 699848
rect 348844 699836 348850 699848
rect 351178 699836 351184 699848
rect 348844 699808 351184 699836
rect 348844 699796 348850 699808
rect 351178 699796 351184 699808
rect 351236 699796 351242 699848
rect 153010 699660 153016 699712
rect 153068 699700 153074 699712
rect 154114 699700 154120 699712
rect 153068 699672 154120 699700
rect 153068 699660 153074 699672
rect 154114 699660 154120 699672
rect 154172 699660 154178 699712
rect 218974 699700 218980 699712
rect 215312 699672 218980 699700
rect 215202 699592 215208 699644
rect 215260 699632 215266 699644
rect 215312 699632 215340 699672
rect 218974 699660 218980 699672
rect 219032 699660 219038 699712
rect 267642 699700 267648 699712
rect 263612 699672 267648 699700
rect 215260 699604 215340 699632
rect 215260 699592 215266 699604
rect 262858 699592 262864 699644
rect 262916 699632 262922 699644
rect 263612 699632 263640 699672
rect 267642 699660 267648 699672
rect 267700 699660 267706 699712
rect 282178 699660 282184 699712
rect 282236 699700 282242 699712
rect 283834 699700 283840 699712
rect 282236 699672 283840 699700
rect 282236 699660 282242 699672
rect 283834 699660 283840 699672
rect 283892 699660 283898 699712
rect 332502 699660 332508 699712
rect 332560 699700 332566 699712
rect 335998 699700 336004 699712
rect 332560 699672 336004 699700
rect 332560 699660 332566 699672
rect 335998 699660 336004 699672
rect 336056 699660 336062 699712
rect 262916 699604 263640 699632
rect 262916 699592 262922 699604
rect 364978 698096 364984 698148
rect 365036 698136 365042 698148
rect 369118 698136 369124 698148
rect 365036 698108 369124 698136
rect 365036 698096 365042 698108
rect 369118 698096 369124 698108
rect 369176 698096 369182 698148
rect 153010 696980 153016 696992
rect 151786 696952 153016 696980
rect 146938 696872 146944 696924
rect 146996 696912 147002 696924
rect 151786 696912 151814 696952
rect 153010 696940 153016 696952
rect 153068 696940 153074 696992
rect 146996 696884 151814 696912
rect 146996 696872 147002 696884
rect 211798 693608 211804 693660
rect 211856 693648 211862 693660
rect 215202 693648 215208 693660
rect 211856 693620 215208 693648
rect 211856 693608 211862 693620
rect 215202 693608 215208 693620
rect 215260 693608 215266 693660
rect 226978 693404 226984 693456
rect 227036 693444 227042 693456
rect 234614 693444 234620 693456
rect 227036 693416 234620 693444
rect 227036 693404 227042 693416
rect 234614 693404 234620 693416
rect 234672 693404 234678 693456
rect 351178 690616 351184 690668
rect 351236 690656 351242 690668
rect 359458 690656 359464 690668
rect 351236 690628 359464 690656
rect 351236 690616 351242 690628
rect 359458 690616 359464 690628
rect 359516 690616 359522 690668
rect 369118 690344 369124 690396
rect 369176 690384 369182 690396
rect 371234 690384 371240 690396
rect 369176 690356 371240 690384
rect 369176 690344 369182 690356
rect 371234 690344 371240 690356
rect 371292 690344 371298 690396
rect 145650 688644 145656 688696
rect 145708 688684 145714 688696
rect 146938 688684 146944 688696
rect 145708 688656 146944 688684
rect 145708 688644 145714 688656
rect 146938 688644 146944 688656
rect 146996 688644 147002 688696
rect 191098 687896 191104 687948
rect 191156 687936 191162 687948
rect 201494 687936 201500 687948
rect 191156 687908 201500 687936
rect 191156 687896 191162 687908
rect 201494 687896 201500 687908
rect 201552 687896 201558 687948
rect 371234 687896 371240 687948
rect 371292 687936 371298 687948
rect 377398 687936 377404 687948
rect 371292 687908 377404 687936
rect 371292 687896 371298 687908
rect 377398 687896 377404 687908
rect 377456 687896 377462 687948
rect 335998 684428 336004 684480
rect 336056 684468 336062 684480
rect 341242 684468 341248 684480
rect 336056 684440 341248 684468
rect 336056 684428 336062 684440
rect 341242 684428 341248 684440
rect 341300 684428 341306 684480
rect 144178 683952 144184 684004
rect 144236 683992 144242 684004
rect 145650 683992 145656 684004
rect 144236 683964 145656 683992
rect 144236 683952 144242 683964
rect 145650 683952 145656 683964
rect 145708 683952 145714 684004
rect 299474 681164 299480 681216
rect 299532 681204 299538 681216
rect 304994 681204 305000 681216
rect 299532 681176 305000 681204
rect 299532 681164 299538 681176
rect 304994 681164 305000 681176
rect 305052 681164 305058 681216
rect 187970 680552 187976 680604
rect 188028 680592 188034 680604
rect 191098 680592 191104 680604
rect 188028 680564 191104 680592
rect 188028 680552 188034 680564
rect 191098 680552 191104 680564
rect 191156 680552 191162 680604
rect 359458 679260 359464 679312
rect 359516 679300 359522 679312
rect 362218 679300 362224 679312
rect 359516 679272 362224 679300
rect 359516 679260 359522 679272
rect 362218 679260 362224 679272
rect 362276 679260 362282 679312
rect 341242 679124 341248 679176
rect 341300 679164 341306 679176
rect 344278 679164 344284 679176
rect 341300 679136 344284 679164
rect 341300 679124 341306 679136
rect 344278 679124 344284 679136
rect 344336 679124 344342 679176
rect 280890 678988 280896 679040
rect 280948 679028 280954 679040
rect 282178 679028 282184 679040
rect 280948 679000 282184 679028
rect 280948 678988 280954 679000
rect 282178 678988 282184 679000
rect 282236 678988 282242 679040
rect 377398 678920 377404 678972
rect 377456 678960 377462 678972
rect 385678 678960 385684 678972
rect 377456 678932 385684 678960
rect 377456 678920 377462 678932
rect 385678 678920 385684 678932
rect 385736 678920 385742 678972
rect 185578 677560 185584 677612
rect 185636 677600 185642 677612
rect 187970 677600 187976 677612
rect 185636 677572 187976 677600
rect 185636 677560 185642 677572
rect 187970 677560 187976 677572
rect 188028 677560 188034 677612
rect 279418 677016 279424 677068
rect 279476 677056 279482 677068
rect 280890 677056 280896 677068
rect 279476 677028 280896 677056
rect 279476 677016 279482 677028
rect 280890 677016 280896 677028
rect 280948 677016 280954 677068
rect 221458 676744 221464 676796
rect 221516 676784 221522 676796
rect 226978 676784 226984 676796
rect 221516 676756 226984 676784
rect 221516 676744 221522 676756
rect 226978 676744 226984 676756
rect 227036 676744 227042 676796
rect 304994 675588 305000 675640
rect 305052 675628 305058 675640
rect 307754 675628 307760 675640
rect 305052 675600 307760 675628
rect 305052 675588 305058 675600
rect 307754 675588 307760 675600
rect 307812 675588 307818 675640
rect 259454 674976 259460 675028
rect 259512 675016 259518 675028
rect 262858 675016 262864 675028
rect 259512 674988 262864 675016
rect 259512 674976 259518 674988
rect 262858 674976 262864 674988
rect 262916 674976 262922 675028
rect 307754 672732 307760 672784
rect 307812 672772 307818 672784
rect 319898 672772 319904 672784
rect 307812 672744 319904 672772
rect 307812 672732 307818 672744
rect 319898 672732 319904 672744
rect 319956 672732 319962 672784
rect 215294 672052 215300 672104
rect 215352 672092 215358 672104
rect 221458 672092 221464 672104
rect 215352 672064 221464 672092
rect 215352 672052 215358 672064
rect 221458 672052 221464 672064
rect 221516 672052 221522 672104
rect 259454 672092 259460 672104
rect 258046 672064 259460 672092
rect 255682 671984 255688 672036
rect 255740 672024 255746 672036
rect 258046 672024 258074 672064
rect 259454 672052 259460 672064
rect 259512 672052 259518 672104
rect 255740 671996 258074 672024
rect 255740 671984 255746 671996
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 15838 670732 15844 670744
rect 3568 670704 15844 670732
rect 3568 670692 3574 670704
rect 15838 670692 15844 670704
rect 15896 670692 15902 670744
rect 144178 670732 144184 670744
rect 142126 670704 144184 670732
rect 140314 670624 140320 670676
rect 140372 670664 140378 670676
rect 142126 670664 142154 670704
rect 144178 670692 144184 670704
rect 144236 670692 144242 670744
rect 407758 670692 407764 670744
rect 407816 670732 407822 670744
rect 580166 670732 580172 670744
rect 407816 670704 580172 670732
rect 407816 670692 407822 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 140372 670636 142154 670664
rect 140372 670624 140378 670636
rect 362218 669944 362224 669996
rect 362276 669984 362282 669996
rect 383930 669984 383936 669996
rect 362276 669956 383936 669984
rect 362276 669944 362282 669956
rect 383930 669944 383936 669956
rect 383988 669944 383994 669996
rect 253198 669332 253204 669384
rect 253256 669372 253262 669384
rect 255682 669372 255688 669384
rect 253256 669344 255688 669372
rect 253256 669332 253262 669344
rect 255682 669332 255688 669344
rect 255740 669332 255746 669384
rect 344278 669264 344284 669316
rect 344336 669304 344342 669316
rect 346670 669304 346676 669316
rect 344336 669276 346676 669304
rect 344336 669264 344342 669276
rect 346670 669264 346676 669276
rect 346728 669264 346734 669316
rect 138658 667904 138664 667956
rect 138716 667944 138722 667956
rect 140314 667944 140320 667956
rect 138716 667916 140320 667944
rect 138716 667904 138722 667916
rect 140314 667904 140320 667916
rect 140372 667904 140378 667956
rect 204898 667156 204904 667208
rect 204956 667196 204962 667208
rect 215294 667196 215300 667208
rect 204956 667168 215300 667196
rect 204956 667156 204962 667168
rect 215294 667156 215300 667168
rect 215352 667156 215358 667208
rect 383930 665796 383936 665848
rect 383988 665836 383994 665848
rect 395338 665836 395344 665848
rect 383988 665808 395344 665836
rect 383988 665796 383994 665808
rect 395338 665796 395344 665808
rect 395396 665796 395402 665848
rect 210418 665116 210424 665168
rect 210476 665156 210482 665168
rect 211798 665156 211804 665168
rect 210476 665128 211804 665156
rect 210476 665116 210482 665128
rect 211798 665116 211804 665128
rect 211856 665116 211862 665168
rect 319898 665116 319904 665168
rect 319956 665156 319962 665168
rect 324958 665156 324964 665168
rect 319956 665128 324964 665156
rect 319956 665116 319962 665128
rect 324958 665116 324964 665128
rect 325016 665116 325022 665168
rect 385678 665116 385684 665168
rect 385736 665156 385742 665168
rect 389818 665156 389824 665168
rect 385736 665128 389824 665156
rect 385736 665116 385742 665128
rect 389818 665116 389824 665128
rect 389876 665116 389882 665168
rect 197262 664436 197268 664488
rect 197320 664476 197326 664488
rect 204898 664476 204904 664488
rect 197320 664448 204904 664476
rect 197320 664436 197326 664448
rect 204898 664436 204904 664448
rect 204956 664436 204962 664488
rect 346670 664436 346676 664488
rect 346728 664476 346734 664488
rect 364978 664476 364984 664488
rect 346728 664448 364984 664476
rect 346728 664436 346734 664448
rect 364978 664436 364984 664448
rect 365036 664436 365042 664488
rect 277486 662396 277492 662448
rect 277544 662436 277550 662448
rect 279418 662436 279424 662448
rect 277544 662408 279424 662436
rect 277544 662396 277550 662408
rect 279418 662396 279424 662408
rect 279476 662396 279482 662448
rect 191098 661036 191104 661088
rect 191156 661076 191162 661088
rect 197262 661076 197268 661088
rect 191156 661048 197268 661076
rect 191156 661036 191162 661048
rect 197262 661036 197268 661048
rect 197320 661036 197326 661088
rect 276658 660560 276664 660612
rect 276716 660600 276722 660612
rect 277486 660600 277492 660612
rect 276716 660572 277492 660600
rect 276716 660560 276722 660572
rect 277486 660560 277492 660572
rect 277544 660560 277550 660612
rect 389818 656820 389824 656872
rect 389876 656860 389882 656872
rect 392578 656860 392584 656872
rect 389876 656832 392584 656860
rect 389876 656820 389882 656832
rect 392578 656820 392584 656832
rect 392636 656820 392642 656872
rect 136726 651380 136732 651432
rect 136784 651420 136790 651432
rect 138658 651420 138664 651432
rect 136784 651392 138664 651420
rect 136784 651380 136790 651392
rect 138658 651380 138664 651392
rect 138716 651380 138722 651432
rect 178034 650632 178040 650684
rect 178092 650672 178098 650684
rect 191098 650672 191104 650684
rect 178092 650644 191104 650672
rect 178092 650632 178098 650644
rect 191098 650632 191104 650644
rect 191156 650632 191162 650684
rect 170398 647844 170404 647896
rect 170456 647884 170462 647896
rect 178034 647884 178040 647896
rect 170456 647856 178040 647884
rect 170456 647844 170462 647856
rect 178034 647844 178040 647856
rect 178092 647844 178098 647896
rect 133690 646824 133696 646876
rect 133748 646864 133754 646876
rect 136726 646864 136732 646876
rect 133748 646836 136732 646864
rect 133748 646824 133754 646836
rect 136726 646824 136732 646836
rect 136784 646824 136790 646876
rect 392578 646144 392584 646196
rect 392636 646184 392642 646196
rect 395522 646184 395528 646196
rect 392636 646156 395528 646184
rect 392636 646144 392642 646156
rect 395522 646144 395528 646156
rect 395580 646144 395586 646196
rect 131758 644444 131764 644496
rect 131816 644484 131822 644496
rect 133690 644484 133696 644496
rect 131816 644456 133696 644484
rect 131816 644444 131822 644456
rect 133690 644444 133696 644456
rect 133748 644444 133754 644496
rect 181438 640296 181444 640348
rect 181496 640336 181502 640348
rect 185578 640336 185584 640348
rect 181496 640308 185584 640336
rect 181496 640296 181502 640308
rect 185578 640296 185584 640308
rect 185636 640296 185642 640348
rect 276658 640336 276664 640348
rect 274652 640308 276664 640336
rect 272518 640228 272524 640280
rect 272576 640268 272582 640280
rect 274652 640268 274680 640308
rect 276658 640296 276664 640308
rect 276716 640296 276722 640348
rect 272576 640240 274680 640268
rect 272576 640228 272582 640240
rect 207658 636216 207664 636268
rect 207716 636256 207722 636268
rect 210418 636256 210424 636268
rect 207716 636228 210424 636256
rect 207716 636216 207722 636228
rect 210418 636216 210424 636228
rect 210476 636216 210482 636268
rect 324958 635468 324964 635520
rect 325016 635508 325022 635520
rect 329190 635508 329196 635520
rect 325016 635480 329196 635508
rect 325016 635468 325022 635480
rect 329190 635468 329196 635480
rect 329248 635468 329254 635520
rect 155218 632680 155224 632732
rect 155276 632720 155282 632732
rect 170398 632720 170404 632732
rect 155276 632692 170404 632720
rect 155276 632680 155282 632692
rect 170398 632680 170404 632692
rect 170456 632680 170462 632732
rect 128354 632068 128360 632120
rect 128412 632108 128418 632120
rect 131758 632108 131764 632120
rect 128412 632080 131764 632108
rect 128412 632068 128418 632080
rect 131758 632068 131764 632080
rect 131816 632068 131822 632120
rect 127618 629688 127624 629740
rect 127676 629728 127682 629740
rect 128354 629728 128360 629740
rect 127676 629700 128360 629728
rect 127676 629688 127682 629700
rect 128354 629688 128360 629700
rect 128412 629688 128418 629740
rect 329190 629212 329196 629264
rect 329248 629252 329254 629264
rect 331858 629252 331864 629264
rect 329248 629224 331864 629252
rect 329248 629212 329254 629224
rect 331858 629212 331864 629224
rect 331916 629212 331922 629264
rect 364978 626492 364984 626544
rect 365036 626532 365042 626544
rect 369118 626532 369124 626544
rect 365036 626504 369124 626532
rect 365036 626492 365042 626504
rect 369118 626492 369124 626504
rect 369176 626492 369182 626544
rect 204898 625200 204904 625252
rect 204956 625240 204962 625252
rect 207658 625240 207664 625252
rect 204956 625212 207664 625240
rect 204956 625200 204962 625212
rect 207658 625200 207664 625212
rect 207716 625200 207722 625252
rect 127618 623812 127624 623824
rect 125612 623784 127624 623812
rect 124214 623704 124220 623756
rect 124272 623744 124278 623756
rect 125612 623744 125640 623784
rect 127618 623772 127624 623784
rect 127676 623772 127682 623824
rect 124272 623716 125640 623744
rect 124272 623704 124278 623716
rect 175918 622684 175924 622736
rect 175976 622724 175982 622736
rect 181438 622724 181444 622736
rect 175976 622696 181444 622724
rect 175976 622684 175982 622696
rect 181438 622684 181444 622696
rect 181496 622684 181502 622736
rect 123478 620984 123484 621036
rect 123536 621024 123542 621036
rect 124214 621024 124220 621036
rect 123536 620996 124220 621024
rect 123536 620984 123542 620996
rect 124214 620984 124220 620996
rect 124272 620984 124278 621036
rect 3510 618264 3516 618316
rect 3568 618304 3574 618316
rect 37918 618304 37924 618316
rect 3568 618276 37924 618304
rect 3568 618264 3574 618276
rect 37918 618264 37924 618276
rect 37976 618264 37982 618316
rect 406378 616836 406384 616888
rect 406436 616876 406442 616888
rect 579982 616876 579988 616888
rect 406436 616848 579988 616876
rect 406436 616836 406442 616848
rect 579982 616836 579988 616848
rect 580040 616836 580046 616888
rect 169018 616088 169024 616140
rect 169076 616128 169082 616140
rect 175918 616128 175924 616140
rect 169076 616100 175924 616128
rect 169076 616088 169082 616100
rect 175918 616088 175924 616100
rect 175976 616088 175982 616140
rect 270494 614116 270500 614168
rect 270552 614156 270558 614168
rect 272518 614156 272524 614168
rect 270552 614128 272524 614156
rect 270552 614116 270558 614128
rect 272518 614116 272524 614128
rect 272576 614116 272582 614168
rect 331858 611260 331864 611312
rect 331916 611300 331922 611312
rect 337378 611300 337384 611312
rect 331916 611272 337384 611300
rect 331916 611260 331922 611272
rect 337378 611260 337384 611272
rect 337436 611260 337442 611312
rect 203518 609220 203524 609272
rect 203576 609260 203582 609272
rect 204898 609260 204904 609272
rect 203576 609232 204904 609260
rect 203576 609220 203582 609232
rect 204898 609220 204904 609232
rect 204956 609220 204962 609272
rect 263594 609220 263600 609272
rect 263652 609260 263658 609272
rect 270494 609260 270500 609272
rect 263652 609232 270500 609260
rect 263652 609220 263658 609232
rect 270494 609220 270500 609232
rect 270552 609220 270558 609272
rect 262858 606568 262864 606620
rect 262916 606608 262922 606620
rect 263594 606608 263600 606620
rect 262916 606580 263600 606608
rect 262916 606568 262922 606580
rect 263594 606568 263600 606580
rect 263652 606568 263658 606620
rect 251910 601672 251916 601724
rect 251968 601712 251974 601724
rect 253198 601712 253204 601724
rect 251968 601684 253204 601712
rect 251968 601672 251974 601684
rect 253198 601672 253204 601684
rect 253256 601672 253262 601724
rect 123478 600352 123484 600364
rect 122806 600324 123484 600352
rect 120718 600244 120724 600296
rect 120776 600284 120782 600296
rect 122806 600284 122834 600324
rect 123478 600312 123484 600324
rect 123536 600312 123542 600364
rect 120776 600256 122834 600284
rect 120776 600244 120782 600256
rect 261478 598612 261484 598664
rect 261536 598652 261542 598664
rect 262858 598652 262864 598664
rect 261536 598624 262864 598652
rect 261536 598612 261542 598624
rect 262858 598612 262864 598624
rect 262916 598612 262922 598664
rect 250438 596912 250444 596964
rect 250496 596952 250502 596964
rect 251910 596952 251916 596964
rect 250496 596924 251916 596952
rect 250496 596912 250502 596924
rect 251910 596912 251916 596924
rect 251968 596912 251974 596964
rect 337378 592220 337384 592272
rect 337436 592260 337442 592272
rect 339494 592260 339500 592272
rect 337436 592232 339500 592260
rect 337436 592220 337442 592232
rect 339494 592220 339500 592232
rect 339552 592220 339558 592272
rect 112438 591268 112444 591320
rect 112496 591308 112502 591320
rect 120718 591308 120724 591320
rect 112496 591280 120724 591308
rect 112496 591268 112502 591280
rect 120718 591268 120724 591280
rect 120776 591268 120782 591320
rect 339494 590588 339500 590640
rect 339552 590628 339558 590640
rect 343634 590628 343640 590640
rect 339552 590600 343640 590628
rect 339552 590588 339558 590600
rect 343634 590588 343640 590600
rect 343692 590588 343698 590640
rect 343634 587596 343640 587648
rect 343692 587636 343698 587648
rect 347038 587636 347044 587648
rect 343692 587608 347044 587636
rect 343692 587596 343698 587608
rect 347038 587596 347044 587608
rect 347096 587596 347102 587648
rect 250438 586548 250444 586560
rect 247052 586520 250444 586548
rect 246298 586440 246304 586492
rect 246356 586480 246362 586492
rect 247052 586480 247080 586520
rect 250438 586508 250444 586520
rect 250496 586508 250502 586560
rect 246356 586452 247080 586480
rect 246356 586440 246362 586452
rect 369118 582224 369124 582276
rect 369176 582264 369182 582276
rect 373258 582264 373264 582276
rect 369176 582236 373264 582264
rect 369176 582224 369182 582236
rect 373258 582224 373264 582236
rect 373316 582224 373322 582276
rect 144178 571956 144184 572008
rect 144236 571996 144242 572008
rect 155218 571996 155224 572008
rect 144236 571968 155224 571996
rect 144236 571956 144242 571968
rect 155218 571956 155224 571968
rect 155276 571956 155282 572008
rect 3326 565836 3332 565888
rect 3384 565876 3390 565888
rect 19978 565876 19984 565888
rect 3384 565848 19984 565876
rect 3384 565836 3390 565848
rect 19978 565836 19984 565848
rect 20036 565836 20042 565888
rect 111058 565836 111064 565888
rect 111116 565876 111122 565888
rect 112438 565876 112444 565888
rect 111116 565848 112444 565876
rect 111116 565836 111122 565848
rect 112438 565836 112444 565848
rect 112496 565836 112502 565888
rect 243538 564408 243544 564460
rect 243596 564448 243602 564460
rect 246298 564448 246304 564460
rect 243596 564420 246304 564448
rect 243596 564408 243602 564420
rect 246298 564408 246304 564420
rect 246356 564408 246362 564460
rect 140774 563048 140780 563100
rect 140832 563088 140838 563100
rect 144178 563088 144184 563100
rect 140832 563060 144184 563088
rect 140832 563048 140838 563060
rect 144178 563048 144184 563060
rect 144236 563048 144242 563100
rect 260098 563048 260104 563100
rect 260156 563088 260162 563100
rect 261478 563088 261484 563100
rect 260156 563060 261484 563088
rect 260156 563048 260162 563060
rect 261478 563048 261484 563060
rect 261536 563048 261542 563100
rect 404998 563048 405004 563100
rect 405056 563088 405062 563100
rect 580166 563088 580172 563100
rect 405056 563060 580172 563088
rect 405056 563048 405062 563060
rect 580166 563048 580172 563060
rect 580224 563048 580230 563100
rect 373258 562980 373264 563032
rect 373316 563020 373322 563032
rect 376662 563020 376668 563032
rect 373316 562992 376668 563020
rect 373316 562980 373322 562992
rect 376662 562980 376668 562992
rect 376720 562980 376726 563032
rect 347038 562300 347044 562352
rect 347096 562340 347102 562352
rect 349798 562340 349804 562352
rect 347096 562312 349804 562340
rect 347096 562300 347102 562312
rect 349798 562300 349804 562312
rect 349856 562300 349862 562352
rect 127618 560940 127624 560992
rect 127676 560980 127682 560992
rect 140774 560980 140780 560992
rect 127676 560952 140780 560980
rect 127676 560940 127682 560952
rect 140774 560940 140780 560952
rect 140832 560940 140838 560992
rect 376662 559512 376668 559564
rect 376720 559552 376726 559564
rect 383654 559552 383660 559564
rect 376720 559524 383660 559552
rect 376720 559512 376726 559524
rect 383654 559512 383660 559524
rect 383712 559512 383718 559564
rect 202138 558832 202144 558884
rect 202196 558872 202202 558884
rect 203518 558872 203524 558884
rect 202196 558844 203524 558872
rect 202196 558832 202202 558844
rect 203518 558832 203524 558844
rect 203576 558832 203582 558884
rect 383654 556724 383660 556776
rect 383712 556764 383718 556776
rect 389818 556764 389824 556776
rect 383712 556736 389824 556764
rect 383712 556724 383718 556736
rect 389818 556724 389824 556736
rect 389876 556724 389882 556776
rect 349798 555432 349804 555484
rect 349856 555472 349862 555484
rect 368382 555472 368388 555484
rect 349856 555444 368388 555472
rect 349856 555432 349862 555444
rect 368382 555432 368388 555444
rect 368440 555432 368446 555484
rect 117222 554004 117228 554056
rect 117280 554044 117286 554056
rect 127618 554044 127624 554056
rect 117280 554016 127624 554044
rect 117280 554004 117286 554016
rect 127618 554004 127624 554016
rect 127676 554004 127682 554056
rect 2774 553800 2780 553852
rect 2832 553840 2838 553852
rect 4798 553840 4804 553852
rect 2832 553812 4804 553840
rect 2832 553800 2838 553812
rect 4798 553800 4804 553812
rect 4856 553800 4862 553852
rect 109678 551284 109684 551336
rect 109736 551324 109742 551336
rect 111058 551324 111064 551336
rect 109736 551296 111064 551324
rect 109736 551284 109742 551296
rect 111058 551284 111064 551296
rect 111116 551284 111122 551336
rect 104986 549856 104992 549908
rect 105044 549896 105050 549908
rect 117222 549896 117228 549908
rect 105044 549868 117228 549896
rect 105044 549856 105050 549868
rect 117222 549856 117228 549868
rect 117280 549856 117286 549908
rect 368382 549856 368388 549908
rect 368440 549896 368446 549908
rect 382918 549896 382924 549908
rect 368440 549868 382924 549896
rect 368440 549856 368446 549868
rect 382918 549856 382924 549868
rect 382976 549856 382982 549908
rect 94498 542988 94504 543040
rect 94556 543028 94562 543040
rect 104986 543028 104992 543040
rect 94556 543000 104992 543028
rect 94556 542988 94562 543000
rect 104986 542988 104992 543000
rect 105044 542988 105050 543040
rect 389818 537956 389824 538008
rect 389876 537996 389882 538008
rect 395154 537996 395160 538008
rect 389876 537968 395160 537996
rect 389876 537956 389882 537968
rect 395154 537956 395160 537968
rect 395212 537956 395218 538008
rect 83458 537548 83464 537600
rect 83516 537588 83522 537600
rect 94498 537588 94504 537600
rect 83516 537560 94504 537588
rect 83516 537548 83522 537560
rect 94498 537548 94504 537560
rect 94556 537548 94562 537600
rect 62666 537480 62672 537532
rect 62724 537520 62730 537532
rect 169754 537520 169760 537532
rect 62724 537492 169760 537520
rect 62724 537480 62730 537492
rect 169754 537480 169760 537492
rect 169812 537480 169818 537532
rect 395154 534080 395160 534132
rect 395212 534120 395218 534132
rect 397546 534120 397552 534132
rect 395212 534092 397552 534120
rect 395212 534080 395218 534092
rect 397546 534080 397552 534092
rect 397604 534080 397610 534132
rect 61378 532992 61384 533044
rect 61436 533032 61442 533044
rect 62666 533032 62672 533044
rect 61436 533004 62672 533032
rect 61436 532992 61442 533004
rect 62666 532992 62672 533004
rect 62724 532992 62730 533044
rect 257062 528572 257068 528624
rect 257120 528612 257126 528624
rect 260098 528612 260104 528624
rect 257120 528584 260104 528612
rect 257120 528572 257126 528584
rect 260098 528572 260104 528584
rect 260156 528572 260162 528624
rect 382918 528028 382924 528080
rect 382976 528068 382982 528080
rect 386322 528068 386328 528080
rect 382976 528040 386328 528068
rect 382976 528028 382982 528040
rect 386322 528028 386328 528040
rect 386380 528028 386386 528080
rect 386322 522928 386328 522980
rect 386380 522968 386386 522980
rect 391198 522968 391204 522980
rect 386380 522940 391204 522968
rect 386380 522928 386386 522940
rect 391198 522928 391204 522940
rect 391256 522928 391262 522980
rect 255958 522112 255964 522164
rect 256016 522152 256022 522164
rect 257062 522152 257068 522164
rect 256016 522124 257068 522152
rect 256016 522112 256022 522124
rect 257062 522112 257068 522124
rect 257120 522112 257126 522164
rect 243538 520316 243544 520328
rect 240152 520288 243544 520316
rect 239398 520208 239404 520260
rect 239456 520248 239462 520260
rect 240152 520248 240180 520288
rect 243538 520276 243544 520288
rect 243596 520276 243602 520328
rect 239456 520220 240180 520248
rect 239456 520208 239462 520220
rect 109678 516168 109684 516180
rect 106384 516140 109684 516168
rect 105538 516060 105544 516112
rect 105596 516100 105602 516112
rect 106384 516100 106412 516140
rect 109678 516128 109684 516140
rect 109736 516128 109742 516180
rect 105596 516072 106412 516100
rect 105596 516060 105602 516072
rect 3326 514768 3332 514820
rect 3384 514808 3390 514820
rect 42058 514808 42064 514820
rect 3384 514780 42064 514808
rect 3384 514768 3390 514780
rect 42058 514768 42064 514780
rect 42116 514768 42122 514820
rect 80054 512932 80060 512984
rect 80112 512972 80118 512984
rect 83458 512972 83464 512984
rect 80112 512944 83464 512972
rect 80112 512932 80118 512944
rect 83458 512932 83464 512944
rect 83516 512932 83522 512984
rect 253198 511912 253204 511964
rect 253256 511952 253262 511964
rect 255958 511952 255964 511964
rect 253256 511924 255964 511952
rect 253256 511912 253262 511924
rect 255958 511912 255964 511924
rect 256016 511912 256022 511964
rect 403618 510620 403624 510672
rect 403676 510660 403682 510672
rect 579798 510660 579804 510672
rect 403676 510632 579804 510660
rect 403676 510620 403682 510632
rect 579798 510620 579804 510632
rect 579856 510620 579862 510672
rect 69474 509872 69480 509924
rect 69532 509912 69538 509924
rect 80054 509912 80060 509924
rect 69532 509884 80060 509912
rect 69532 509872 69538 509884
rect 80054 509872 80060 509884
rect 80112 509872 80118 509924
rect 117958 508512 117964 508564
rect 118016 508552 118022 508564
rect 136634 508552 136640 508564
rect 118016 508524 136640 508552
rect 118016 508512 118022 508524
rect 136634 508512 136640 508524
rect 136692 508512 136698 508564
rect 61470 504364 61476 504416
rect 61528 504404 61534 504416
rect 69474 504404 69480 504416
rect 61528 504376 69480 504404
rect 61528 504364 61534 504376
rect 69474 504364 69480 504376
rect 69532 504364 69538 504416
rect 200758 502936 200764 502988
rect 200816 502976 200822 502988
rect 202138 502976 202144 502988
rect 200816 502948 202144 502976
rect 200816 502936 200822 502948
rect 202138 502936 202144 502948
rect 202196 502936 202202 502988
rect 2774 501032 2780 501084
rect 2832 501072 2838 501084
rect 4890 501072 4896 501084
rect 2832 501044 4896 501072
rect 2832 501032 2838 501044
rect 4890 501032 4896 501044
rect 4948 501032 4954 501084
rect 158714 498788 158720 498840
rect 158772 498828 158778 498840
rect 169018 498828 169024 498840
rect 158772 498800 169024 498828
rect 158772 498788 158778 498800
rect 169018 498788 169024 498800
rect 169076 498788 169082 498840
rect 391198 498380 391204 498432
rect 391256 498420 391262 498432
rect 393958 498420 393964 498432
rect 391256 498392 393964 498420
rect 391256 498380 391262 498392
rect 393958 498380 393964 498392
rect 394016 498380 394022 498432
rect 253198 494068 253204 494080
rect 251192 494040 253204 494068
rect 250438 493960 250444 494012
rect 250496 494000 250502 494012
rect 251192 494000 251220 494040
rect 253198 494028 253204 494040
rect 253256 494028 253262 494080
rect 250496 493972 251220 494000
rect 250496 493960 250502 493972
rect 150434 490560 150440 490612
rect 150492 490600 150498 490612
rect 158714 490600 158720 490612
rect 150492 490572 158720 490600
rect 150492 490560 150498 490572
rect 158714 490560 158720 490572
rect 158772 490560 158778 490612
rect 116578 487160 116584 487212
rect 116636 487200 116642 487212
rect 117958 487200 117964 487212
rect 116636 487172 117964 487200
rect 116636 487160 116642 487172
rect 117958 487160 117964 487172
rect 118016 487160 118022 487212
rect 146018 487160 146024 487212
rect 146076 487200 146082 487212
rect 150434 487200 150440 487212
rect 146076 487172 150440 487200
rect 146076 487160 146082 487172
rect 150434 487160 150440 487172
rect 150492 487160 150498 487212
rect 237374 486480 237380 486532
rect 237432 486520 237438 486532
rect 239398 486520 239404 486532
rect 237432 486492 239404 486520
rect 237432 486480 237438 486492
rect 239398 486480 239404 486492
rect 239456 486480 239462 486532
rect 142798 484304 142804 484356
rect 142856 484344 142862 484356
rect 146018 484344 146024 484356
rect 142856 484316 146024 484344
rect 142856 484304 142862 484316
rect 146018 484304 146024 484316
rect 146076 484304 146082 484356
rect 236638 482536 236644 482588
rect 236696 482576 236702 482588
rect 237374 482576 237380 482588
rect 236696 482548 237380 482576
rect 236696 482536 236702 482548
rect 237374 482536 237380 482548
rect 237432 482536 237438 482588
rect 135162 479476 135168 479528
rect 135220 479516 135226 479528
rect 142798 479516 142804 479528
rect 135220 479488 142804 479516
rect 135220 479476 135226 479488
rect 142798 479476 142804 479488
rect 142856 479476 142862 479528
rect 249426 478864 249432 478916
rect 249484 478904 249490 478916
rect 250438 478904 250444 478916
rect 249484 478876 250444 478904
rect 249484 478864 249490 478876
rect 250438 478864 250444 478876
rect 250496 478864 250502 478916
rect 129734 476280 129740 476332
rect 129792 476320 129798 476332
rect 135162 476320 135168 476332
rect 129792 476292 135168 476320
rect 129792 476280 129798 476292
rect 135162 476280 135168 476292
rect 135220 476280 135226 476332
rect 393958 475396 393964 475448
rect 394016 475436 394022 475448
rect 395430 475436 395436 475448
rect 394016 475408 395436 475436
rect 394016 475396 394022 475408
rect 395430 475396 395436 475408
rect 395488 475396 395494 475448
rect 58618 474648 58624 474700
rect 58676 474688 58682 474700
rect 61470 474688 61476 474700
rect 58676 474660 61476 474688
rect 58676 474648 58682 474660
rect 61470 474648 61476 474660
rect 61528 474648 61534 474700
rect 247678 474376 247684 474428
rect 247736 474416 247742 474428
rect 249426 474416 249432 474428
rect 247736 474388 249432 474416
rect 247736 474376 247742 474388
rect 249426 474376 249432 474388
rect 249484 474376 249490 474428
rect 115198 472948 115204 473000
rect 115256 472988 115262 473000
rect 116578 472988 116584 473000
rect 115256 472960 116584 472988
rect 115256 472948 115262 472960
rect 116578 472948 116584 472960
rect 116636 472948 116642 473000
rect 199378 471996 199384 472048
rect 199436 472036 199442 472048
rect 200758 472036 200764 472048
rect 199436 472008 200764 472036
rect 199436 471996 199442 472008
rect 200758 471996 200764 472008
rect 200816 471996 200822 472048
rect 120718 471248 120724 471300
rect 120776 471288 120782 471300
rect 129734 471288 129740 471300
rect 120776 471260 129740 471288
rect 120776 471248 120782 471260
rect 129734 471248 129740 471260
rect 129792 471248 129798 471300
rect 197998 469208 198004 469260
rect 198056 469248 198062 469260
rect 199378 469248 199384 469260
rect 198056 469220 199384 469248
rect 198056 469208 198062 469220
rect 199378 469208 199384 469220
rect 199436 469208 199442 469260
rect 55858 466420 55864 466472
rect 55916 466460 55922 466472
rect 58618 466460 58624 466472
rect 55916 466432 58624 466460
rect 55916 466420 55922 466432
rect 58618 466420 58624 466432
rect 58676 466420 58682 466472
rect 2774 462544 2780 462596
rect 2832 462584 2838 462596
rect 5074 462584 5080 462596
rect 2832 462556 5080 462584
rect 2832 462544 2838 462556
rect 5074 462544 5080 462556
rect 5132 462544 5138 462596
rect 197998 456804 198004 456816
rect 195992 456776 198004 456804
rect 193858 456696 193864 456748
rect 193916 456736 193922 456748
rect 195992 456736 196020 456776
rect 197998 456764 198004 456776
rect 198056 456764 198062 456816
rect 400858 456764 400864 456816
rect 400916 456804 400922 456816
rect 579982 456804 579988 456816
rect 400916 456776 579988 456804
rect 400916 456764 400922 456776
rect 579982 456764 579988 456776
rect 580040 456764 580046 456816
rect 193916 456708 196020 456736
rect 193916 456696 193922 456708
rect 46198 451868 46204 451920
rect 46256 451908 46262 451920
rect 55858 451908 55864 451920
rect 46256 451880 55864 451908
rect 46256 451868 46262 451880
rect 55858 451868 55864 451880
rect 55916 451868 55922 451920
rect 117958 449896 117964 449948
rect 118016 449936 118022 449948
rect 120718 449936 120724 449948
rect 118016 449908 120724 449936
rect 118016 449896 118022 449908
rect 120718 449896 120724 449908
rect 120776 449896 120782 449948
rect 2774 448808 2780 448860
rect 2832 448848 2838 448860
rect 4982 448848 4988 448860
rect 2832 448820 4988 448848
rect 2832 448808 2838 448820
rect 4982 448808 4988 448820
rect 5040 448808 5046 448860
rect 399570 444388 399576 444440
rect 399628 444428 399634 444440
rect 580074 444428 580080 444440
rect 399628 444400 580080 444428
rect 399628 444388 399634 444400
rect 580074 444388 580080 444400
rect 580132 444388 580138 444440
rect 45094 428272 45100 428324
rect 45152 428312 45158 428324
rect 46198 428312 46204 428324
rect 45152 428284 46204 428312
rect 45152 428272 45158 428284
rect 46198 428272 46204 428284
rect 46256 428272 46262 428324
rect 111058 427048 111064 427100
rect 111116 427088 111122 427100
rect 117958 427088 117964 427100
rect 111116 427060 117964 427088
rect 111116 427048 111122 427060
rect 117958 427048 117964 427060
rect 118016 427048 118022 427100
rect 192478 425688 192484 425740
rect 192536 425728 192542 425740
rect 193858 425728 193864 425740
rect 192536 425700 193864 425728
rect 192536 425688 192542 425700
rect 193858 425688 193864 425700
rect 193916 425688 193922 425740
rect 247678 419540 247684 419552
rect 245672 419512 247684 419540
rect 244918 419432 244924 419484
rect 244976 419472 244982 419484
rect 245672 419472 245700 419512
rect 247678 419500 247684 419512
rect 247736 419500 247742 419552
rect 244976 419444 245700 419472
rect 244976 419432 244982 419444
rect 398098 418140 398104 418192
rect 398156 418180 398162 418192
rect 580074 418180 580080 418192
rect 398156 418152 580080 418180
rect 398156 418140 398162 418152
rect 580074 418140 580080 418152
rect 580132 418140 580138 418192
rect 102778 412632 102784 412684
rect 102836 412672 102842 412684
rect 105538 412672 105544 412684
rect 102836 412644 105544 412672
rect 102836 412632 102842 412644
rect 105538 412632 105544 412644
rect 105596 412632 105602 412684
rect 3326 409912 3332 409964
rect 3384 409952 3390 409964
rect 8938 409952 8944 409964
rect 3384 409924 8944 409952
rect 3384 409912 3390 409924
rect 8938 409912 8944 409924
rect 8996 409912 9002 409964
rect 399478 404336 399484 404388
rect 399536 404376 399542 404388
rect 580074 404376 580080 404388
rect 399536 404348 580080 404376
rect 399536 404336 399542 404348
rect 580074 404336 580080 404348
rect 580132 404336 580138 404388
rect 243538 404268 243544 404320
rect 243596 404308 243602 404320
rect 244918 404308 244924 404320
rect 243596 404280 244924 404308
rect 243596 404268 243602 404280
rect 244918 404268 244924 404280
rect 244976 404268 244982 404320
rect 2774 397468 2780 397520
rect 2832 397508 2838 397520
rect 5166 397508 5172 397520
rect 2832 397480 5172 397508
rect 2832 397468 2838 397480
rect 5166 397468 5172 397480
rect 5224 397468 5230 397520
rect 235258 394612 235264 394664
rect 235316 394652 235322 394664
rect 236638 394652 236644 394664
rect 235316 394624 236644 394652
rect 235316 394612 235322 394624
rect 236638 394612 236644 394624
rect 236696 394612 236702 394664
rect 101398 391960 101404 392012
rect 101456 392000 101462 392012
rect 102778 392000 102784 392012
rect 101456 391972 102784 392000
rect 101456 391960 101462 391972
rect 102778 391960 102784 391972
rect 102836 391960 102842 392012
rect 189718 391960 189724 392012
rect 189776 392000 189782 392012
rect 192478 392000 192484 392012
rect 189776 391972 192484 392000
rect 189776 391960 189782 391972
rect 192478 391960 192484 391972
rect 192536 391960 192542 392012
rect 108298 390532 108304 390584
rect 108356 390572 108362 390584
rect 111058 390572 111064 390584
rect 108356 390544 111064 390572
rect 108356 390532 108362 390544
rect 111058 390532 111064 390544
rect 111116 390532 111122 390584
rect 396718 378156 396724 378208
rect 396776 378196 396782 378208
rect 580074 378196 580080 378208
rect 396776 378168 580080 378196
rect 396776 378156 396782 378168
rect 580074 378156 580080 378168
rect 580132 378156 580138 378208
rect 58618 376592 58624 376644
rect 58676 376632 58682 376644
rect 61378 376632 61384 376644
rect 58676 376604 61384 376632
rect 58676 376592 58682 376604
rect 61378 376592 61384 376604
rect 61436 376592 61442 376644
rect 239398 371220 239404 371272
rect 239456 371260 239462 371272
rect 243538 371260 243544 371272
rect 239456 371232 243544 371260
rect 239456 371220 239462 371232
rect 243538 371220 243544 371232
rect 243596 371220 243602 371272
rect 188430 369860 188436 369912
rect 188488 369900 188494 369912
rect 189718 369900 189724 369912
rect 188488 369872 189724 369900
rect 188488 369860 188494 369872
rect 189718 369860 189724 369872
rect 189776 369860 189782 369912
rect 101398 368540 101404 368552
rect 99392 368512 101404 368540
rect 98638 368432 98644 368484
rect 98696 368472 98702 368484
rect 99392 368472 99420 368512
rect 101398 368500 101404 368512
rect 101456 368500 101462 368552
rect 98696 368444 99420 368472
rect 98696 368432 98702 368444
rect 186958 365508 186964 365560
rect 187016 365548 187022 365560
rect 188430 365548 188436 365560
rect 187016 365520 188436 365548
rect 187016 365508 187022 365520
rect 188430 365508 188436 365520
rect 188488 365508 188494 365560
rect 396902 364352 396908 364404
rect 396960 364392 396966 364404
rect 579798 364392 579804 364404
rect 396960 364364 579804 364392
rect 396960 364352 396966 364364
rect 579798 364352 579804 364364
rect 579856 364352 579862 364404
rect 232498 360204 232504 360256
rect 232556 360244 232562 360256
rect 235258 360244 235264 360256
rect 232556 360216 235264 360244
rect 232556 360204 232562 360216
rect 235258 360204 235264 360216
rect 235316 360204 235322 360256
rect 3326 357416 3332 357468
rect 3384 357456 3390 357468
rect 10318 357456 10324 357468
rect 3384 357428 10324 357456
rect 3384 357416 3390 357428
rect 10318 357416 10324 357428
rect 10376 357416 10382 357468
rect 69658 356668 69664 356720
rect 69716 356708 69722 356720
rect 115198 356708 115204 356720
rect 69716 356680 115204 356708
rect 69716 356668 69722 356680
rect 115198 356668 115204 356680
rect 115256 356668 115262 356720
rect 99006 353948 99012 354000
rect 99064 353988 99070 354000
rect 108298 353988 108304 354000
rect 99064 353960 108304 353988
rect 99064 353948 99070 353960
rect 108298 353948 108304 353960
rect 108356 353948 108362 354000
rect 185578 353268 185584 353320
rect 185636 353308 185642 353320
rect 186958 353308 186964 353320
rect 185636 353280 186964 353308
rect 185636 353268 185642 353280
rect 186958 353268 186964 353280
rect 187016 353268 187022 353320
rect 235258 352044 235264 352096
rect 235316 352084 235322 352096
rect 239398 352084 239404 352096
rect 235316 352056 239404 352084
rect 235316 352044 235322 352056
rect 239398 352044 239404 352056
rect 239456 352044 239462 352096
rect 418798 351908 418804 351960
rect 418856 351948 418862 351960
rect 580074 351948 580080 351960
rect 418856 351920 580080 351948
rect 418856 351908 418862 351920
rect 580074 351908 580080 351920
rect 580132 351908 580138 351960
rect 94498 348848 94504 348900
rect 94556 348888 94562 348900
rect 99006 348888 99012 348900
rect 94556 348860 99012 348888
rect 94556 348848 94562 348860
rect 99006 348848 99012 348860
rect 99064 348848 99070 348900
rect 229738 348780 229744 348832
rect 229796 348820 229802 348832
rect 232498 348820 232504 348832
rect 229796 348792 232504 348820
rect 229796 348780 229802 348792
rect 232498 348780 232504 348792
rect 232556 348780 232562 348832
rect 56870 346332 56876 346384
rect 56928 346372 56934 346384
rect 58618 346372 58624 346384
rect 56928 346344 58624 346372
rect 56928 346332 56934 346344
rect 58618 346332 58624 346344
rect 58676 346332 58682 346384
rect 2774 345176 2780 345228
rect 2832 345216 2838 345228
rect 5258 345216 5264 345228
rect 2832 345188 5264 345216
rect 2832 345176 2838 345188
rect 5258 345176 5264 345188
rect 5316 345176 5322 345228
rect 233970 342252 233976 342304
rect 234028 342292 234034 342304
rect 235258 342292 235264 342304
rect 234028 342264 235264 342292
rect 234028 342252 234034 342264
rect 235258 342252 235264 342264
rect 235316 342252 235322 342304
rect 232498 340008 232504 340060
rect 232556 340048 232562 340060
rect 233970 340048 233976 340060
rect 232556 340020 233976 340048
rect 232556 340008 232562 340020
rect 233970 340008 233976 340020
rect 234028 340008 234034 340060
rect 68278 339668 68284 339720
rect 68336 339708 68342 339720
rect 69658 339708 69664 339720
rect 68336 339680 69664 339708
rect 68336 339668 68342 339680
rect 69658 339668 69664 339680
rect 69716 339668 69722 339720
rect 97258 338784 97264 338836
rect 97316 338824 97322 338836
rect 98638 338824 98644 338836
rect 97316 338796 98644 338824
rect 97316 338784 97322 338796
rect 98638 338784 98644 338796
rect 98696 338784 98702 338836
rect 55858 338240 55864 338292
rect 55916 338280 55922 338292
rect 56870 338280 56876 338292
rect 55916 338252 56876 338280
rect 55916 338240 55922 338252
rect 56870 338240 56876 338252
rect 56928 338240 56934 338292
rect 87598 336744 87604 336796
rect 87656 336784 87662 336796
rect 94498 336784 94504 336796
rect 87656 336756 94504 336784
rect 87656 336744 87662 336756
rect 94498 336744 94504 336756
rect 94556 336744 94562 336796
rect 229738 335356 229744 335368
rect 226352 335328 229744 335356
rect 225322 335248 225328 335300
rect 225380 335288 225386 335300
rect 226352 335288 226380 335328
rect 229738 335316 229744 335328
rect 229796 335316 229802 335368
rect 225380 335260 226380 335288
rect 225380 335248 225386 335260
rect 231210 333956 231216 334008
rect 231268 333996 231274 334008
rect 232498 333996 232504 334008
rect 231268 333968 232504 333996
rect 231268 333956 231274 333968
rect 232498 333956 232504 333968
rect 232556 333956 232562 334008
rect 95878 329060 95884 329112
rect 95936 329100 95942 329112
rect 97258 329100 97264 329112
rect 95936 329072 97264 329100
rect 95936 329060 95942 329072
rect 97258 329060 97264 329072
rect 97316 329060 97322 329112
rect 224218 328992 224224 329044
rect 224276 329032 224282 329044
rect 225322 329032 225328 329044
rect 224276 329004 225328 329032
rect 224276 328992 224282 329004
rect 225322 328992 225328 329004
rect 225380 328992 225386 329044
rect 229830 326272 229836 326324
rect 229888 326312 229894 326324
rect 231210 326312 231216 326324
rect 229888 326284 231216 326312
rect 229888 326272 229894 326284
rect 231210 326272 231216 326284
rect 231268 326272 231274 326324
rect 396810 324300 396816 324352
rect 396868 324340 396874 324352
rect 580074 324340 580080 324352
rect 396868 324312 580080 324340
rect 396868 324300 396874 324312
rect 580074 324300 580080 324312
rect 580132 324300 580138 324352
rect 81710 323552 81716 323604
rect 81768 323592 81774 323604
rect 87598 323592 87604 323604
rect 81768 323564 87604 323592
rect 81768 323552 81774 323564
rect 87598 323552 87604 323564
rect 87656 323552 87662 323604
rect 227714 323552 227720 323604
rect 227772 323592 227778 323604
rect 229830 323592 229836 323604
rect 227772 323564 229836 323592
rect 227772 323552 227778 323564
rect 229830 323552 229836 323564
rect 229888 323552 229894 323604
rect 53098 323348 53104 323400
rect 53156 323388 53162 323400
rect 55858 323388 55864 323400
rect 53156 323360 55864 323388
rect 53156 323348 53162 323360
rect 55858 323348 55864 323360
rect 55916 323348 55922 323400
rect 221458 322940 221464 322992
rect 221516 322980 221522 322992
rect 224218 322980 224224 322992
rect 221516 322952 224224 322980
rect 221516 322940 221522 322952
rect 224218 322940 224224 322952
rect 224276 322940 224282 322992
rect 94774 321716 94780 321768
rect 94832 321756 94838 321768
rect 95878 321756 95884 321768
rect 94832 321728 95884 321756
rect 94832 321716 94838 321728
rect 95878 321716 95884 321728
rect 95936 321716 95942 321768
rect 182450 320764 182456 320816
rect 182508 320804 182514 320816
rect 185578 320804 185584 320816
rect 182508 320776 185584 320804
rect 182508 320764 182514 320776
rect 185578 320764 185584 320776
rect 185636 320764 185642 320816
rect 91094 319744 91100 319796
rect 91152 319784 91158 319796
rect 94774 319784 94780 319796
rect 91152 319756 94780 319784
rect 91152 319744 91158 319756
rect 94774 319744 94780 319756
rect 94832 319744 94838 319796
rect 85574 318724 85580 318776
rect 85632 318764 85638 318776
rect 88334 318764 88340 318776
rect 85632 318736 88340 318764
rect 85632 318724 85638 318736
rect 88334 318724 88340 318736
rect 88392 318724 88398 318776
rect 180794 318656 180800 318708
rect 180852 318696 180858 318708
rect 182450 318696 182456 318708
rect 180852 318668 182456 318696
rect 180852 318656 180858 318668
rect 182450 318656 182456 318668
rect 182508 318656 182514 318708
rect 223114 318248 223120 318300
rect 223172 318288 223178 318300
rect 227714 318288 227720 318300
rect 223172 318260 227720 318288
rect 223172 318248 223178 318260
rect 227714 318248 227720 318260
rect 227772 318248 227778 318300
rect 91094 317472 91100 317484
rect 89732 317444 91100 317472
rect 88334 317364 88340 317416
rect 88392 317404 88398 317416
rect 89732 317404 89760 317444
rect 91094 317432 91100 317444
rect 91152 317432 91158 317484
rect 88392 317376 89760 317404
rect 88392 317364 88398 317376
rect 79226 316752 79232 316804
rect 79284 316792 79290 316804
rect 81710 316792 81716 316804
rect 79284 316764 81716 316792
rect 79284 316752 79290 316764
rect 81710 316752 81716 316764
rect 81768 316752 81774 316804
rect 62758 313896 62764 313948
rect 62816 313936 62822 313948
rect 104894 313936 104900 313948
rect 62816 313908 104900 313936
rect 62816 313896 62822 313908
rect 104894 313896 104900 313908
rect 104952 313896 104958 313948
rect 178678 313624 178684 313676
rect 178736 313664 178742 313676
rect 180794 313664 180800 313676
rect 178736 313636 180800 313664
rect 178736 313624 178742 313636
rect 180794 313624 180800 313636
rect 180852 313624 180858 313676
rect 79318 313352 79324 313404
rect 79376 313392 79382 313404
rect 85574 313392 85580 313404
rect 79376 313364 85580 313392
rect 79376 313352 79382 313364
rect 85574 313352 85580 313364
rect 85632 313352 85638 313404
rect 220078 313284 220084 313336
rect 220136 313324 220142 313336
rect 221458 313324 221464 313336
rect 220136 313296 221464 313324
rect 220136 313284 220142 313296
rect 221458 313284 221464 313296
rect 221516 313284 221522 313336
rect 220170 311856 220176 311908
rect 220228 311896 220234 311908
rect 223114 311896 223120 311908
rect 220228 311868 223120 311896
rect 220228 311856 220234 311868
rect 223114 311856 223120 311868
rect 223172 311856 223178 311908
rect 397086 311856 397092 311908
rect 397144 311896 397150 311908
rect 580074 311896 580080 311908
rect 397144 311868 580080 311896
rect 397144 311856 397150 311868
rect 580074 311856 580080 311868
rect 580132 311856 580138 311908
rect 69658 311108 69664 311160
rect 69716 311148 69722 311160
rect 79226 311148 79232 311160
rect 69716 311120 79232 311148
rect 69716 311108 69722 311120
rect 79226 311108 79232 311120
rect 79284 311108 79290 311160
rect 85390 309408 85396 309460
rect 85448 309448 85454 309460
rect 88242 309448 88248 309460
rect 85448 309420 88248 309448
rect 85448 309408 85454 309420
rect 88242 309408 88248 309420
rect 88300 309408 88306 309460
rect 81342 307776 81348 307828
rect 81400 307816 81406 307828
rect 85390 307816 85396 307828
rect 81400 307788 85396 307816
rect 81400 307776 81406 307788
rect 85390 307776 85396 307788
rect 85448 307776 85454 307828
rect 3234 304988 3240 305040
rect 3292 305028 3298 305040
rect 24118 305028 24124 305040
rect 3292 305000 24124 305028
rect 3292 304988 3298 305000
rect 24118 304988 24124 305000
rect 24176 304988 24182 305040
rect 51718 304988 51724 305040
rect 51776 305028 51782 305040
rect 53098 305028 53104 305040
rect 51776 305000 53104 305028
rect 51776 304988 51782 305000
rect 53098 304988 53104 305000
rect 53156 304988 53162 305040
rect 67174 303628 67180 303680
rect 67232 303668 67238 303680
rect 69658 303668 69664 303680
rect 67232 303640 69664 303668
rect 67232 303628 67238 303640
rect 69658 303628 69664 303640
rect 69716 303628 69722 303680
rect 57238 301452 57244 301504
rect 57296 301492 57302 301504
rect 79318 301492 79324 301504
rect 57296 301464 79324 301492
rect 57296 301452 57302 301464
rect 79318 301452 79324 301464
rect 79376 301452 79382 301504
rect 61378 301044 61384 301096
rect 61436 301084 61442 301096
rect 62758 301084 62764 301096
rect 61436 301056 62764 301084
rect 61436 301044 61442 301056
rect 62758 301044 62764 301056
rect 62816 301044 62822 301096
rect 79318 300296 79324 300348
rect 79376 300336 79382 300348
rect 81342 300336 81348 300348
rect 79376 300308 81348 300336
rect 79376 300296 79382 300308
rect 81342 300296 81348 300308
rect 81400 300296 81406 300348
rect 66898 300160 66904 300212
rect 66956 300200 66962 300212
rect 68278 300200 68284 300212
rect 66956 300172 68284 300200
rect 66956 300160 66962 300172
rect 68278 300160 68284 300172
rect 68336 300160 68342 300212
rect 51810 300092 51816 300144
rect 51868 300132 51874 300144
rect 67174 300132 67180 300144
rect 51868 300104 67180 300132
rect 51868 300092 51874 300104
rect 67174 300092 67180 300104
rect 67232 300092 67238 300144
rect 417418 298120 417424 298172
rect 417476 298160 417482 298172
rect 580074 298160 580080 298172
rect 417476 298132 580080 298160
rect 417476 298120 417482 298132
rect 580074 298120 580080 298132
rect 580132 298120 580138 298172
rect 3234 292544 3240 292596
rect 3292 292584 3298 292596
rect 43438 292584 43444 292596
rect 3292 292556 43444 292584
rect 3292 292544 3298 292556
rect 43438 292544 43444 292556
rect 43496 292544 43502 292596
rect 76558 292544 76564 292596
rect 76616 292584 76622 292596
rect 79318 292584 79324 292596
rect 76616 292556 79324 292584
rect 76616 292544 76622 292556
rect 79318 292544 79324 292556
rect 79376 292544 79382 292596
rect 218054 292544 218060 292596
rect 218112 292584 218118 292596
rect 220170 292584 220176 292596
rect 218112 292556 220176 292584
rect 218112 292544 218118 292556
rect 220170 292544 220176 292556
rect 220228 292544 220234 292596
rect 215938 289824 215944 289876
rect 215996 289864 216002 289876
rect 218054 289864 218060 289876
rect 215996 289836 218060 289864
rect 215996 289824 216002 289836
rect 218054 289824 218060 289836
rect 218112 289824 218118 289876
rect 55858 288328 55864 288380
rect 55916 288368 55922 288380
rect 57238 288368 57244 288380
rect 55916 288340 57244 288368
rect 55916 288328 55922 288340
rect 57238 288328 57244 288340
rect 57296 288328 57302 288380
rect 49602 287580 49608 287632
rect 49660 287620 49666 287632
rect 51810 287620 51816 287632
rect 49660 287592 51816 287620
rect 49660 287580 49666 287592
rect 51810 287580 51816 287592
rect 51868 287580 51874 287632
rect 46198 284316 46204 284368
rect 46256 284356 46262 284368
rect 49602 284356 49608 284368
rect 46256 284328 49608 284356
rect 46256 284316 46262 284328
rect 49602 284316 49608 284328
rect 49660 284316 49666 284368
rect 72050 281936 72056 281988
rect 72108 281976 72114 281988
rect 76558 281976 76564 281988
rect 72108 281948 76564 281976
rect 72108 281936 72114 281948
rect 76558 281936 76564 281948
rect 76616 281936 76622 281988
rect 59998 280780 60004 280832
rect 60056 280820 60062 280832
rect 61378 280820 61384 280832
rect 60056 280792 61384 280820
rect 60056 280780 60062 280792
rect 61378 280780 61384 280792
rect 61436 280780 61442 280832
rect 213914 279964 213920 280016
rect 213972 280004 213978 280016
rect 215938 280004 215944 280016
rect 213972 279976 215944 280004
rect 213972 279964 213978 279976
rect 215938 279964 215944 279976
rect 215996 279964 216002 280016
rect 69474 279692 69480 279744
rect 69532 279732 69538 279744
rect 72050 279732 72056 279744
rect 69532 279704 72056 279732
rect 69532 279692 69538 279704
rect 72050 279692 72056 279704
rect 72108 279692 72114 279744
rect 175918 276020 175924 276072
rect 175976 276060 175982 276072
rect 178678 276060 178684 276072
rect 175976 276032 178684 276060
rect 175976 276020 175982 276032
rect 178678 276020 178684 276032
rect 178736 276020 178742 276072
rect 218054 276020 218060 276072
rect 218112 276060 218118 276072
rect 220078 276060 220084 276072
rect 218112 276032 220084 276060
rect 218112 276020 218118 276032
rect 220078 276020 220084 276032
rect 220136 276020 220142 276072
rect 204162 275272 204168 275324
rect 204220 275312 204226 275324
rect 213914 275312 213920 275324
rect 204220 275284 213920 275312
rect 204220 275272 204226 275284
rect 213914 275272 213920 275284
rect 213972 275272 213978 275324
rect 45002 274728 45008 274780
rect 45060 274768 45066 274780
rect 46198 274768 46204 274780
rect 45060 274740 46204 274768
rect 45060 274728 45066 274740
rect 46198 274728 46204 274740
rect 46256 274728 46262 274780
rect 57974 274660 57980 274712
rect 58032 274700 58038 274712
rect 59998 274700 60004 274712
rect 58032 274672 60004 274700
rect 58032 274660 58038 274672
rect 59998 274660 60004 274672
rect 60056 274660 60062 274712
rect 54478 272892 54484 272944
rect 54536 272932 54542 272944
rect 55858 272932 55864 272944
rect 54536 272904 55864 272932
rect 54536 272892 54542 272904
rect 55858 272892 55864 272904
rect 55916 272892 55922 272944
rect 202138 271872 202144 271924
rect 202196 271912 202202 271924
rect 204162 271912 204168 271924
rect 202196 271884 204168 271912
rect 202196 271872 202202 271884
rect 204162 271872 204168 271884
rect 204220 271872 204226 271924
rect 396994 271872 397000 271924
rect 397052 271912 397058 271924
rect 579798 271912 579804 271924
rect 397052 271884 579804 271912
rect 397052 271872 397058 271884
rect 579798 271872 579804 271884
rect 579856 271872 579862 271924
rect 69474 270552 69480 270564
rect 67652 270524 69480 270552
rect 65518 270444 65524 270496
rect 65576 270484 65582 270496
rect 67652 270484 67680 270524
rect 69474 270512 69480 270524
rect 69532 270512 69538 270564
rect 217962 270552 217968 270564
rect 213932 270524 217968 270552
rect 65576 270456 67680 270484
rect 65576 270444 65582 270456
rect 213362 270444 213368 270496
rect 213420 270484 213426 270496
rect 213932 270484 213960 270524
rect 217962 270512 217968 270524
rect 218020 270512 218026 270564
rect 213420 270456 213960 270484
rect 213420 270444 213426 270456
rect 52362 269084 52368 269136
rect 52420 269124 52426 269136
rect 57882 269124 57888 269136
rect 52420 269096 57888 269124
rect 52420 269084 52426 269096
rect 57882 269084 57888 269096
rect 57940 269084 57946 269136
rect 63494 266500 63500 266552
rect 63552 266540 63558 266552
rect 66898 266540 66904 266552
rect 63552 266512 66904 266540
rect 63552 266500 63558 266512
rect 66898 266500 66904 266512
rect 66956 266500 66962 266552
rect 51074 266364 51080 266416
rect 51132 266404 51138 266416
rect 54478 266404 54484 266416
rect 51132 266376 54484 266404
rect 51132 266364 51138 266376
rect 54478 266364 54484 266376
rect 54536 266364 54542 266416
rect 202138 266404 202144 266416
rect 200086 266376 202144 266404
rect 197722 266296 197728 266348
rect 197780 266336 197786 266348
rect 200086 266336 200114 266376
rect 202138 266364 202144 266376
rect 202196 266364 202202 266416
rect 197780 266308 200114 266336
rect 197780 266296 197786 266308
rect 208394 264188 208400 264240
rect 208452 264228 208458 264240
rect 213362 264228 213368 264240
rect 208452 264200 213368 264228
rect 208452 264188 208458 264200
rect 213362 264188 213368 264200
rect 213420 264188 213426 264240
rect 50338 262828 50344 262880
rect 50396 262868 50402 262880
rect 63494 262868 63500 262880
rect 50396 262840 63500 262868
rect 50396 262828 50402 262840
rect 63494 262828 63500 262840
rect 63552 262828 63558 262880
rect 195238 261808 195244 261860
rect 195296 261848 195302 261860
rect 197722 261848 197728 261860
rect 195296 261820 197728 261848
rect 195296 261808 195302 261820
rect 197722 261808 197728 261820
rect 197780 261808 197786 261860
rect 189074 261468 189080 261520
rect 189132 261508 189138 261520
rect 208302 261508 208308 261520
rect 189132 261480 208308 261508
rect 189132 261468 189138 261480
rect 208302 261468 208308 261480
rect 208360 261468 208366 261520
rect 50890 261196 50896 261248
rect 50948 261236 50954 261248
rect 52362 261236 52368 261248
rect 50948 261208 52368 261236
rect 50948 261196 50954 261208
rect 52362 261196 52368 261208
rect 52420 261196 52426 261248
rect 174262 260788 174268 260840
rect 174320 260828 174326 260840
rect 175918 260828 175924 260840
rect 174320 260800 175924 260828
rect 174320 260788 174326 260800
rect 175918 260788 175924 260800
rect 175976 260788 175982 260840
rect 47578 260448 47584 260500
rect 47636 260488 47642 260500
rect 51074 260488 51080 260500
rect 47636 260460 51080 260488
rect 47636 260448 47642 260460
rect 51074 260448 51080 260460
rect 51132 260448 51138 260500
rect 65518 259468 65524 259480
rect 60752 259440 65524 259468
rect 60642 259360 60648 259412
rect 60700 259400 60706 259412
rect 60752 259400 60780 259440
rect 65518 259428 65524 259440
rect 65576 259428 65582 259480
rect 189074 259468 189080 259480
rect 187712 259440 189080 259468
rect 60700 259372 60780 259400
rect 60700 259360 60706 259372
rect 185578 259360 185584 259412
rect 185636 259400 185642 259412
rect 187712 259400 187740 259440
rect 189074 259428 189080 259440
rect 189132 259428 189138 259480
rect 185636 259372 187740 259400
rect 185636 259360 185642 259372
rect 49234 258952 49240 259004
rect 49292 258992 49298 259004
rect 50890 258992 50896 259004
rect 49292 258964 50896 258992
rect 49292 258952 49298 258964
rect 50890 258952 50896 258964
rect 50948 258952 50954 259004
rect 397178 258068 397184 258120
rect 397236 258108 397242 258120
rect 579982 258108 579988 258120
rect 397236 258080 579988 258108
rect 397236 258068 397242 258080
rect 579982 258068 579988 258080
rect 580040 258068 580046 258120
rect 47486 256708 47492 256760
rect 47544 256748 47550 256760
rect 49234 256748 49240 256760
rect 47544 256720 49240 256748
rect 47544 256708 47550 256720
rect 49234 256708 49240 256720
rect 49292 256708 49298 256760
rect 193858 256708 193864 256760
rect 193916 256748 193922 256760
rect 195238 256748 195244 256760
rect 193916 256720 195244 256748
rect 193916 256708 193922 256720
rect 195238 256708 195244 256720
rect 195296 256708 195302 256760
rect 3142 253920 3148 253972
rect 3200 253960 3206 253972
rect 22738 253960 22744 253972
rect 3200 253932 22744 253960
rect 3200 253920 3206 253932
rect 22738 253920 22744 253932
rect 22796 253920 22802 253972
rect 45830 253920 45836 253972
rect 45888 253960 45894 253972
rect 47486 253960 47492 253972
rect 45888 253932 47492 253960
rect 45888 253920 45894 253932
rect 47486 253920 47492 253932
rect 47544 253920 47550 253972
rect 48682 252560 48688 252612
rect 48740 252600 48746 252612
rect 50338 252600 50344 252612
rect 48740 252572 50344 252600
rect 48740 252560 48746 252572
rect 50338 252560 50344 252572
rect 50396 252560 50402 252612
rect 173158 252492 173164 252544
rect 173216 252532 173222 252544
rect 174262 252532 174268 252544
rect 173216 252504 174268 252532
rect 173216 252492 173222 252504
rect 174262 252492 174268 252504
rect 174320 252492 174326 252544
rect 57974 251880 57980 251932
rect 58032 251920 58038 251932
rect 60642 251920 60648 251932
rect 58032 251892 60648 251920
rect 58032 251880 58038 251892
rect 60642 251880 60648 251892
rect 60700 251880 60706 251932
rect 47670 251812 47676 251864
rect 47728 251852 47734 251864
rect 71774 251852 71780 251864
rect 47728 251824 71780 251852
rect 47728 251812 47734 251824
rect 71774 251812 71780 251824
rect 71832 251812 71838 251864
rect 46934 249432 46940 249484
rect 46992 249472 46998 249484
rect 48682 249472 48688 249484
rect 46992 249444 48688 249472
rect 46992 249432 46998 249444
rect 48682 249432 48688 249444
rect 48740 249432 48746 249484
rect 52454 249024 52460 249076
rect 52512 249064 52518 249076
rect 57974 249064 57980 249076
rect 52512 249036 57980 249064
rect 52512 249024 52518 249036
rect 57974 249024 57980 249036
rect 58032 249024 58038 249076
rect 49694 247052 49700 247104
rect 49752 247092 49758 247104
rect 51718 247092 51724 247104
rect 49752 247064 51724 247092
rect 49752 247052 49758 247064
rect 51718 247052 51724 247064
rect 51776 247052 51782 247104
rect 173158 247092 173164 247104
rect 167012 247064 173164 247092
rect 166258 246984 166264 247036
rect 166316 247024 166322 247036
rect 167012 247024 167040 247064
rect 173158 247052 173164 247064
rect 173216 247052 173222 247104
rect 185578 247092 185584 247104
rect 183572 247064 185584 247092
rect 166316 246996 167040 247024
rect 166316 246984 166322 246996
rect 182910 246984 182916 247036
rect 182968 247024 182974 247036
rect 183572 247024 183600 247064
rect 185578 247052 185584 247064
rect 185636 247052 185642 247104
rect 182968 246996 183600 247024
rect 182968 246984 182974 246996
rect 414658 244264 414664 244316
rect 414716 244304 414722 244316
rect 579982 244304 579988 244316
rect 414716 244276 579988 244304
rect 414716 244264 414722 244276
rect 579982 244264 579988 244276
rect 580040 244264 580046 244316
rect 44818 243856 44824 243908
rect 44876 243896 44882 243908
rect 46842 243896 46848 243908
rect 44876 243868 46848 243896
rect 44876 243856 44882 243868
rect 46842 243856 46848 243868
rect 46900 243856 46906 243908
rect 45738 243516 45744 243568
rect 45796 243556 45802 243568
rect 49694 243556 49700 243568
rect 45796 243528 49700 243556
rect 45796 243516 45802 243528
rect 49694 243516 49700 243528
rect 49752 243516 49758 243568
rect 47118 241680 47124 241732
rect 47176 241720 47182 241732
rect 52362 241720 52368 241732
rect 47176 241692 52368 241720
rect 47176 241680 47182 241692
rect 52362 241680 52368 241692
rect 52420 241680 52426 241732
rect 45646 241408 45652 241460
rect 45704 241448 45710 241460
rect 47670 241448 47676 241460
rect 45704 241420 47676 241448
rect 45704 241408 45710 241420
rect 47670 241408 47676 241420
rect 47728 241408 47734 241460
rect 45554 241340 45560 241392
rect 45612 241380 45618 241392
rect 47578 241380 47584 241392
rect 45612 241352 47584 241380
rect 45612 241340 45618 241352
rect 47578 241340 47584 241352
rect 47636 241340 47642 241392
rect 45370 240864 45376 240916
rect 45428 240904 45434 240916
rect 166258 240904 166264 240916
rect 45428 240876 166264 240904
rect 45428 240864 45434 240876
rect 166258 240864 166264 240876
rect 166316 240864 166322 240916
rect 45278 240796 45284 240848
rect 45336 240836 45342 240848
rect 182910 240836 182916 240848
rect 45336 240808 182916 240836
rect 45336 240796 45342 240808
rect 182910 240796 182916 240808
rect 182968 240796 182974 240848
rect 44910 240728 44916 240780
rect 44968 240768 44974 240780
rect 193858 240768 193864 240780
rect 44968 240740 193864 240768
rect 44968 240728 44974 240740
rect 193858 240728 193864 240740
rect 193916 240728 193922 240780
rect 3050 240116 3056 240168
rect 3108 240156 3114 240168
rect 43530 240156 43536 240168
rect 3108 240128 43536 240156
rect 3108 240116 3114 240128
rect 43530 240116 43536 240128
rect 43588 240116 43594 240168
rect 47118 240156 47124 240168
rect 45526 240128 47124 240156
rect 45526 240100 45554 240128
rect 47118 240116 47124 240128
rect 47176 240116 47182 240168
rect 45462 240048 45468 240100
rect 45520 240060 45554 240100
rect 45520 240048 45526 240060
rect 395430 240048 395436 240100
rect 395488 240088 395494 240100
rect 396534 240088 396540 240100
rect 395488 240060 396540 240088
rect 395488 240048 395494 240060
rect 396534 240048 396540 240060
rect 396592 240048 396598 240100
rect 396534 238824 396540 238876
rect 396592 238824 396598 238876
rect 45186 238756 45192 238808
rect 45244 238796 45250 238808
rect 45830 238796 45836 238808
rect 45244 238768 45836 238796
rect 45244 238756 45250 238768
rect 45830 238756 45836 238768
rect 45888 238756 45894 238808
rect 396552 238796 396580 238824
rect 396046 238768 396580 238796
rect 396046 238728 396074 238768
rect 396534 238728 396540 238740
rect 396046 238700 396540 238728
rect 396534 238688 396540 238700
rect 396592 238688 396598 238740
rect 44818 233180 44824 233232
rect 44876 233220 44882 233232
rect 45830 233220 45836 233232
rect 44876 233192 45836 233220
rect 44876 233180 44882 233192
rect 45830 233180 45836 233192
rect 45888 233180 45894 233232
rect 45186 232908 45192 232960
rect 45244 232948 45250 232960
rect 45244 232920 64874 232948
rect 45244 232908 45250 232920
rect 45526 232444 46980 232472
rect 45526 232416 45554 232444
rect 45462 232364 45468 232416
rect 45520 232376 45554 232416
rect 45520 232364 45526 232376
rect 46952 232348 46980 232444
rect 64846 232404 64874 232920
rect 86310 232404 86316 232416
rect 64846 232376 86316 232404
rect 86310 232364 86316 232376
rect 86368 232364 86374 232416
rect 45370 232296 45376 232348
rect 45428 232336 45434 232348
rect 46842 232336 46848 232348
rect 45428 232308 46848 232336
rect 45428 232296 45434 232308
rect 46842 232296 46848 232308
rect 46900 232296 46906 232348
rect 46934 232296 46940 232348
rect 46992 232296 46998 232348
rect 45278 232228 45284 232280
rect 45336 232268 45342 232280
rect 46198 232268 46204 232280
rect 45336 232240 46204 232268
rect 45336 232228 45342 232240
rect 46198 232228 46204 232240
rect 46256 232228 46262 232280
rect 45738 232160 45744 232212
rect 45796 232200 45802 232212
rect 53190 232200 53196 232212
rect 45796 232172 53196 232200
rect 45796 232160 45802 232172
rect 53190 232160 53196 232172
rect 53248 232160 53254 232212
rect 394694 232092 394700 232144
rect 394752 232132 394758 232144
rect 396534 232132 396540 232144
rect 394752 232104 396540 232132
rect 394752 232092 394758 232104
rect 396534 232092 396540 232104
rect 396592 232092 396598 232144
rect 44910 231140 44916 231192
rect 44968 231180 44974 231192
rect 52362 231180 52368 231192
rect 44968 231152 52368 231180
rect 44968 231140 44974 231152
rect 52362 231140 52368 231152
rect 52420 231140 52426 231192
rect 86310 231140 86316 231192
rect 86368 231180 86374 231192
rect 153194 231180 153200 231192
rect 86368 231152 153200 231180
rect 86368 231140 86374 231152
rect 153194 231140 153200 231152
rect 153252 231140 153258 231192
rect 4062 231072 4068 231124
rect 4120 231112 4126 231124
rect 177850 231112 177856 231124
rect 4120 231084 177856 231112
rect 4120 231072 4126 231084
rect 177850 231072 177856 231084
rect 177908 231072 177914 231124
rect 394694 230500 394700 230512
rect 389192 230472 394700 230500
rect 46198 230392 46204 230444
rect 46256 230432 46262 230444
rect 48958 230432 48964 230444
rect 46256 230404 48964 230432
rect 46256 230392 46262 230404
rect 48958 230392 48964 230404
rect 49016 230392 49022 230444
rect 387794 230392 387800 230444
rect 387852 230432 387858 230444
rect 389192 230432 389220 230472
rect 394694 230460 394700 230472
rect 394752 230460 394758 230512
rect 387852 230404 389220 230432
rect 387852 230392 387858 230404
rect 45830 230324 45836 230376
rect 45888 230364 45894 230376
rect 47578 230364 47584 230376
rect 45888 230336 47584 230364
rect 45888 230324 45894 230336
rect 47578 230324 47584 230336
rect 47636 230324 47642 230376
rect 46934 230256 46940 230308
rect 46992 230296 46998 230308
rect 52454 230296 52460 230308
rect 46992 230268 52460 230296
rect 46992 230256 46998 230268
rect 52454 230256 52460 230268
rect 52512 230256 52518 230308
rect 166258 229712 166264 229764
rect 166316 229752 166322 229764
rect 176654 229752 176660 229764
rect 166316 229724 176660 229752
rect 166316 229712 166322 229724
rect 176654 229712 176660 229724
rect 176712 229712 176718 229764
rect 391934 229100 391940 229152
rect 391992 229140 391998 229152
rect 394602 229140 394608 229152
rect 391992 229112 394608 229140
rect 391992 229100 391998 229112
rect 394602 229100 394608 229112
rect 394660 229100 394666 229152
rect 157978 228420 157984 228472
rect 158036 228460 158042 228472
rect 266538 228460 266544 228472
rect 158036 228432 266544 228460
rect 158036 228420 158042 228432
rect 266538 228420 266544 228432
rect 266596 228420 266602 228472
rect 297358 228420 297364 228472
rect 297416 228460 297422 228472
rect 327074 228460 327080 228472
rect 297416 228432 327080 228460
rect 297416 228420 297422 228432
rect 327074 228420 327080 228432
rect 327132 228420 327138 228472
rect 117222 228352 117228 228404
rect 117280 228392 117286 228404
rect 138658 228392 138664 228404
rect 117280 228364 138664 228392
rect 117280 228352 117286 228364
rect 138658 228352 138664 228364
rect 138716 228352 138722 228404
rect 153194 228352 153200 228404
rect 153252 228392 153258 228404
rect 165062 228392 165068 228404
rect 153252 228364 165068 228392
rect 153252 228352 153258 228364
rect 165062 228352 165068 228364
rect 165120 228352 165126 228404
rect 236638 228352 236644 228404
rect 236696 228392 236702 228404
rect 386506 228392 386512 228404
rect 236696 228364 386512 228392
rect 236696 228352 236702 228364
rect 386506 228352 386512 228364
rect 386564 228352 386570 228404
rect 46934 228284 46940 228336
rect 46992 228324 46998 228336
rect 52546 228324 52552 228336
rect 46992 228296 52552 228324
rect 46992 228284 46998 228296
rect 52546 228284 52552 228296
rect 52604 228284 52610 228336
rect 52362 228080 52368 228132
rect 52420 228120 52426 228132
rect 53834 228120 53840 228132
rect 52420 228092 53840 228120
rect 52420 228080 52426 228092
rect 53834 228080 53840 228092
rect 53892 228080 53898 228132
rect 53190 227536 53196 227588
rect 53248 227576 53254 227588
rect 57238 227576 57244 227588
rect 53248 227548 57244 227576
rect 53248 227536 53254 227548
rect 57238 227536 57244 227548
rect 57296 227536 57302 227588
rect 165062 227196 165068 227248
rect 165120 227236 165126 227248
rect 170398 227236 170404 227248
rect 165120 227208 170404 227236
rect 165120 227196 165126 227208
rect 170398 227196 170404 227208
rect 170456 227196 170462 227248
rect 52546 226992 52552 227044
rect 52604 227032 52610 227044
rect 59262 227032 59268 227044
rect 52604 227004 59268 227032
rect 52604 226992 52610 227004
rect 59262 226992 59268 227004
rect 59320 226992 59326 227044
rect 53834 226312 53840 226364
rect 53892 226352 53898 226364
rect 53892 226324 55214 226352
rect 53892 226312 53898 226324
rect 55186 226284 55214 226324
rect 56962 226284 56968 226296
rect 55186 226256 56968 226284
rect 56962 226244 56968 226256
rect 57020 226244 57026 226296
rect 391842 224992 391848 225004
rect 389192 224964 391848 224992
rect 387794 224884 387800 224936
rect 387852 224924 387858 224936
rect 389192 224924 389220 224964
rect 391842 224952 391848 224964
rect 391900 224952 391906 225004
rect 387852 224896 389220 224924
rect 387852 224884 387858 224896
rect 384942 223660 384948 223712
rect 385000 223700 385006 223712
rect 387702 223700 387708 223712
rect 385000 223672 387708 223700
rect 385000 223660 385006 223672
rect 387702 223660 387708 223672
rect 387760 223660 387766 223712
rect 59262 223592 59268 223644
rect 59320 223632 59326 223644
rect 59320 223604 60780 223632
rect 59320 223592 59326 223604
rect 52454 223524 52460 223576
rect 52512 223564 52518 223576
rect 55766 223564 55772 223576
rect 52512 223536 55772 223564
rect 52512 223524 52518 223536
rect 55766 223524 55772 223536
rect 55824 223524 55830 223576
rect 60752 223564 60780 223604
rect 66990 223564 66996 223576
rect 60752 223536 66996 223564
rect 66990 223524 66996 223536
rect 67048 223524 67054 223576
rect 387058 223524 387064 223576
rect 387116 223564 387122 223576
rect 390370 223564 390376 223576
rect 387116 223536 390376 223564
rect 387116 223524 387122 223536
rect 390370 223524 390376 223536
rect 390428 223524 390434 223576
rect 56962 222844 56968 222896
rect 57020 222884 57026 222896
rect 58618 222884 58624 222896
rect 57020 222856 58624 222884
rect 57020 222844 57026 222856
rect 58618 222844 58624 222856
rect 58676 222844 58682 222896
rect 45002 220804 45008 220856
rect 45060 220844 45066 220856
rect 47670 220844 47676 220856
rect 45060 220816 47676 220844
rect 45060 220804 45066 220816
rect 47670 220804 47676 220816
rect 47728 220804 47734 220856
rect 48958 220804 48964 220856
rect 49016 220844 49022 220856
rect 49016 220816 52500 220844
rect 49016 220804 49022 220816
rect 52472 220776 52500 220816
rect 53926 220776 53932 220788
rect 52472 220748 53932 220776
rect 53926 220736 53932 220748
rect 53984 220736 53990 220788
rect 55766 220736 55772 220788
rect 55824 220776 55830 220788
rect 62758 220776 62764 220788
rect 55824 220748 62764 220776
rect 55824 220736 55830 220748
rect 62758 220736 62764 220748
rect 62816 220736 62822 220788
rect 66990 220736 66996 220788
rect 67048 220776 67054 220788
rect 69658 220776 69664 220788
rect 67048 220748 69664 220776
rect 67048 220736 67054 220748
rect 69658 220736 69664 220748
rect 69716 220736 69722 220788
rect 385034 220464 385040 220516
rect 385092 220504 385098 220516
rect 387702 220504 387708 220516
rect 385092 220476 387708 220504
rect 385092 220464 385098 220476
rect 387702 220464 387708 220476
rect 387760 220464 387766 220516
rect 381354 219444 381360 219496
rect 381412 219484 381418 219496
rect 384942 219484 384948 219496
rect 381412 219456 384948 219484
rect 381412 219444 381418 219456
rect 384942 219444 384948 219456
rect 385000 219444 385006 219496
rect 384298 218084 384304 218136
rect 384356 218124 384362 218136
rect 387058 218124 387064 218136
rect 384356 218096 387064 218124
rect 384356 218084 384362 218096
rect 387058 218084 387064 218096
rect 387116 218084 387122 218136
rect 115842 218016 115848 218068
rect 115900 218056 115906 218068
rect 579798 218056 579804 218068
rect 115900 218028 579804 218056
rect 115900 218016 115906 218028
rect 579798 218016 579804 218028
rect 579856 218016 579862 218068
rect 47578 217404 47584 217456
rect 47636 217444 47642 217456
rect 53834 217444 53840 217456
rect 47636 217416 53840 217444
rect 47636 217404 47642 217416
rect 53834 217404 53840 217416
rect 53892 217404 53898 217456
rect 58618 216656 58624 216708
rect 58676 216696 58682 216708
rect 58676 216668 60780 216696
rect 58676 216656 58682 216668
rect 60752 216628 60780 216668
rect 65518 216628 65524 216640
rect 60752 216600 65524 216628
rect 65518 216588 65524 216600
rect 65576 216588 65582 216640
rect 53926 215908 53932 215960
rect 53984 215948 53990 215960
rect 63402 215948 63408 215960
rect 53984 215920 63408 215948
rect 53984 215908 53990 215920
rect 63402 215908 63408 215920
rect 63460 215908 63466 215960
rect 53834 215296 53840 215348
rect 53892 215336 53898 215348
rect 53892 215308 55214 215336
rect 53892 215296 53898 215308
rect 55186 215268 55214 215308
rect 56686 215268 56692 215280
rect 55186 215240 56692 215268
rect 56686 215228 56692 215240
rect 56744 215228 56750 215280
rect 3142 213936 3148 213988
rect 3200 213976 3206 213988
rect 175366 213976 175372 213988
rect 3200 213948 175372 213976
rect 3200 213936 3206 213948
rect 175366 213936 175372 213948
rect 175424 213936 175430 213988
rect 385034 213976 385040 213988
rect 383626 213948 385040 213976
rect 380894 213868 380900 213920
rect 380952 213908 380958 213920
rect 383626 213908 383654 213948
rect 385034 213936 385040 213948
rect 385092 213936 385098 213988
rect 380952 213880 383654 213908
rect 380952 213868 380958 213880
rect 378778 213596 378784 213648
rect 378836 213636 378842 213648
rect 381354 213636 381360 213648
rect 378836 213608 381360 213636
rect 378836 213596 378842 213608
rect 381354 213596 381360 213608
rect 381412 213596 381418 213648
rect 57238 213188 57244 213240
rect 57296 213228 57302 213240
rect 71038 213228 71044 213240
rect 57296 213200 71044 213228
rect 57296 213188 57302 213200
rect 71038 213188 71044 213200
rect 71096 213188 71102 213240
rect 378134 211624 378140 211676
rect 378192 211664 378198 211676
rect 380894 211664 380900 211676
rect 378192 211636 380900 211664
rect 378192 211624 378198 211636
rect 380894 211624 380900 211636
rect 380952 211624 380958 211676
rect 56686 211148 56692 211200
rect 56744 211188 56750 211200
rect 56744 211160 60780 211188
rect 56744 211148 56750 211160
rect 47670 211080 47676 211132
rect 47728 211120 47734 211132
rect 51350 211120 51356 211132
rect 47728 211092 51356 211120
rect 47728 211080 47734 211092
rect 51350 211080 51356 211092
rect 51408 211080 51414 211132
rect 60752 211120 60780 211160
rect 62114 211120 62120 211132
rect 60752 211092 62120 211120
rect 62114 211080 62120 211092
rect 62172 211080 62178 211132
rect 63494 210196 63500 210248
rect 63552 210236 63558 210248
rect 65610 210236 65616 210248
rect 63552 210208 65616 210236
rect 63552 210196 63558 210208
rect 65610 210196 65616 210208
rect 65668 210196 65674 210248
rect 393314 209924 393320 209976
rect 393372 209964 393378 209976
rect 397546 209964 397552 209976
rect 393372 209936 397552 209964
rect 393372 209924 393378 209936
rect 397546 209924 397552 209936
rect 397604 209924 397610 209976
rect 45094 208360 45100 208412
rect 45152 208400 45158 208412
rect 46382 208400 46388 208412
rect 45152 208372 46388 208400
rect 45152 208360 45158 208372
rect 46382 208360 46388 208372
rect 46440 208360 46446 208412
rect 69658 208360 69664 208412
rect 69716 208400 69722 208412
rect 69716 208372 70440 208400
rect 69716 208360 69722 208372
rect 70412 208332 70440 208372
rect 72418 208332 72424 208344
rect 70412 208304 72424 208332
rect 72418 208292 72424 208304
rect 72476 208292 72482 208344
rect 62114 207612 62120 207664
rect 62172 207652 62178 207664
rect 63494 207652 63500 207664
rect 62172 207624 63500 207652
rect 62172 207612 62178 207624
rect 63494 207612 63500 207624
rect 63552 207612 63558 207664
rect 65518 207000 65524 207052
rect 65576 207040 65582 207052
rect 65576 207012 67680 207040
rect 65576 207000 65582 207012
rect 67652 206972 67680 207012
rect 69658 206972 69664 206984
rect 67652 206944 69664 206972
rect 69658 206932 69664 206944
rect 69716 206932 69722 206984
rect 382918 206252 382924 206304
rect 382976 206292 382982 206304
rect 393314 206292 393320 206304
rect 382976 206264 393320 206292
rect 382976 206252 382982 206264
rect 393314 206252 393320 206264
rect 393372 206252 393378 206304
rect 62758 205640 62764 205692
rect 62816 205680 62822 205692
rect 62816 205652 64874 205680
rect 62816 205640 62822 205652
rect 64846 205612 64874 205652
rect 188338 205640 188344 205692
rect 188396 205680 188402 205692
rect 579982 205680 579988 205692
rect 188396 205652 579988 205680
rect 188396 205640 188402 205652
rect 579982 205640 579988 205652
rect 580040 205640 580046 205692
rect 65518 205612 65524 205624
rect 64846 205584 65524 205612
rect 65518 205572 65524 205584
rect 65576 205572 65582 205624
rect 65610 205436 65616 205488
rect 65668 205476 65674 205488
rect 66898 205476 66904 205488
rect 65668 205448 66904 205476
rect 65668 205436 65674 205448
rect 66898 205436 66904 205448
rect 66956 205436 66962 205488
rect 51350 204892 51356 204944
rect 51408 204932 51414 204944
rect 58618 204932 58624 204944
rect 51408 204904 58624 204932
rect 51408 204892 51414 204904
rect 58618 204892 58624 204904
rect 58676 204892 58682 204944
rect 375742 204620 375748 204672
rect 375800 204660 375806 204672
rect 378042 204660 378048 204672
rect 375800 204632 378048 204660
rect 375800 204620 375806 204632
rect 378042 204620 378048 204632
rect 378100 204620 378106 204672
rect 71038 203532 71044 203584
rect 71096 203572 71102 203584
rect 95142 203572 95148 203584
rect 71096 203544 95148 203572
rect 71096 203532 71102 203544
rect 95142 203532 95148 203544
rect 95200 203532 95206 203584
rect 366358 203532 366364 203584
rect 366416 203572 366422 203584
rect 375742 203572 375748 203584
rect 366416 203544 375748 203572
rect 366416 203532 366422 203544
rect 375742 203532 375748 203544
rect 375800 203532 375806 203584
rect 377122 202988 377128 203040
rect 377180 203028 377186 203040
rect 378778 203028 378784 203040
rect 377180 203000 378784 203028
rect 377180 202988 377186 203000
rect 378778 202988 378784 203000
rect 378836 202988 378842 203040
rect 63494 202172 63500 202224
rect 63552 202212 63558 202224
rect 66254 202212 66260 202224
rect 63552 202184 66260 202212
rect 63552 202172 63558 202184
rect 66254 202172 66260 202184
rect 66312 202172 66318 202224
rect 3142 201492 3148 201544
rect 3200 201532 3206 201544
rect 22830 201532 22836 201544
rect 3200 201504 22836 201532
rect 3200 201492 3206 201504
rect 22830 201492 22836 201504
rect 22888 201492 22894 201544
rect 46382 201424 46388 201476
rect 46440 201464 46446 201476
rect 47578 201464 47584 201476
rect 46440 201436 47584 201464
rect 46440 201424 46446 201436
rect 47578 201424 47584 201436
rect 47636 201424 47642 201476
rect 95142 200744 95148 200796
rect 95200 200784 95206 200796
rect 104894 200784 104900 200796
rect 95200 200756 104900 200784
rect 95200 200744 95206 200756
rect 104894 200744 104900 200756
rect 104952 200744 104958 200796
rect 375374 200744 375380 200796
rect 375432 200784 375438 200796
rect 377122 200784 377128 200796
rect 375432 200756 377128 200784
rect 375432 200744 375438 200756
rect 377122 200744 377128 200756
rect 377180 200744 377186 200796
rect 155954 199384 155960 199436
rect 156012 199424 156018 199436
rect 296714 199424 296720 199436
rect 156012 199396 296720 199424
rect 156012 199384 156018 199396
rect 296714 199384 296720 199396
rect 296772 199384 296778 199436
rect 72418 199180 72424 199232
rect 72476 199220 72482 199232
rect 75270 199220 75276 199232
rect 72476 199192 75276 199220
rect 72476 199180 72482 199192
rect 75270 199180 75276 199192
rect 75328 199180 75334 199232
rect 66254 198704 66260 198756
rect 66312 198744 66318 198756
rect 68186 198744 68192 198756
rect 66312 198716 68192 198744
rect 66312 198704 66318 198716
rect 68186 198704 68192 198716
rect 68244 198704 68250 198756
rect 170398 198704 170404 198756
rect 170456 198744 170462 198756
rect 171778 198744 171784 198756
rect 170456 198716 171784 198744
rect 170456 198704 170462 198716
rect 171778 198704 171784 198716
rect 171836 198704 171842 198756
rect 104894 198500 104900 198552
rect 104952 198540 104958 198552
rect 108298 198540 108304 198552
rect 104952 198512 108304 198540
rect 104952 198500 104958 198512
rect 108298 198500 108304 198512
rect 108356 198500 108362 198552
rect 65518 198092 65524 198144
rect 65576 198132 65582 198144
rect 66254 198132 66260 198144
rect 65576 198104 66260 198132
rect 65576 198092 65582 198104
rect 66254 198092 66260 198104
rect 66312 198092 66318 198144
rect 148962 197956 148968 198008
rect 149020 197996 149026 198008
rect 207014 197996 207020 198008
rect 149020 197968 207020 197996
rect 149020 197956 149026 197968
rect 207014 197956 207020 197968
rect 207072 197956 207078 198008
rect 154482 197412 154488 197464
rect 154540 197452 154546 197464
rect 155954 197452 155960 197464
rect 154540 197424 155960 197452
rect 154540 197412 154546 197424
rect 155954 197412 155960 197424
rect 156012 197412 156018 197464
rect 364978 197344 364984 197396
rect 365036 197384 365042 197396
rect 366358 197384 366364 197396
rect 365036 197356 366364 197384
rect 365036 197344 365042 197356
rect 366358 197344 366364 197356
rect 366416 197344 366422 197396
rect 379514 197344 379520 197396
rect 379572 197384 379578 197396
rect 382918 197384 382924 197396
rect 379572 197356 382924 197384
rect 379572 197344 379578 197356
rect 382918 197344 382924 197356
rect 382976 197344 382982 197396
rect 152734 197276 152740 197328
rect 152792 197316 152798 197328
rect 157978 197316 157984 197328
rect 152792 197288 157984 197316
rect 152792 197276 152798 197288
rect 157978 197276 157984 197288
rect 158036 197276 158042 197328
rect 147950 196732 147956 196784
rect 148008 196772 148014 196784
rect 166258 196772 166264 196784
rect 148008 196744 166264 196772
rect 148008 196732 148014 196744
rect 166258 196732 166264 196744
rect 166316 196732 166322 196784
rect 160830 196664 160836 196716
rect 160888 196704 160894 196716
rect 236638 196704 236644 196716
rect 160888 196676 236644 196704
rect 160888 196664 160894 196676
rect 236638 196664 236644 196676
rect 236696 196664 236702 196716
rect 151170 196596 151176 196648
rect 151228 196636 151234 196648
rect 235994 196636 236000 196648
rect 151228 196608 236000 196636
rect 151228 196596 151234 196608
rect 235994 196596 236000 196608
rect 236052 196596 236058 196648
rect 66898 196460 66904 196512
rect 66956 196500 66962 196512
rect 68278 196500 68284 196512
rect 66956 196472 68284 196500
rect 66956 196460 66962 196472
rect 68278 196460 68284 196472
rect 68336 196460 68342 196512
rect 58618 196256 58624 196308
rect 58676 196296 58682 196308
rect 61378 196296 61384 196308
rect 58676 196268 61384 196296
rect 58676 196256 58682 196268
rect 61378 196256 61384 196268
rect 61436 196256 61442 196308
rect 68186 195984 68192 196036
rect 68244 196024 68250 196036
rect 68244 195996 69060 196024
rect 68244 195984 68250 195996
rect 69032 195956 69060 195996
rect 71038 195956 71044 195968
rect 69032 195928 71044 195956
rect 71038 195916 71044 195928
rect 71096 195916 71102 195968
rect 138658 195916 138664 195968
rect 138716 195956 138722 195968
rect 141418 195956 141424 195968
rect 138716 195928 141424 195956
rect 138716 195916 138722 195928
rect 141418 195916 141424 195928
rect 141476 195916 141482 195968
rect 157518 195916 157524 195968
rect 157576 195956 157582 195968
rect 356054 195956 356060 195968
rect 157576 195928 356060 195956
rect 157576 195916 157582 195928
rect 356054 195916 356060 195928
rect 356112 195916 356118 195968
rect 86954 195848 86960 195900
rect 87012 195888 87018 195900
rect 139394 195888 139400 195900
rect 87012 195860 139400 195888
rect 87012 195848 87018 195860
rect 139394 195848 139400 195860
rect 139452 195848 139458 195900
rect 157426 195848 157432 195900
rect 157484 195888 157490 195900
rect 297358 195888 297364 195900
rect 157484 195860 297364 195888
rect 157484 195848 157490 195860
rect 297358 195848 297364 195860
rect 297416 195848 297422 195900
rect 56594 195780 56600 195832
rect 56652 195820 56658 195832
rect 138106 195820 138112 195832
rect 56652 195792 138112 195820
rect 56652 195780 56658 195792
rect 138106 195780 138112 195792
rect 138164 195780 138170 195832
rect 66254 195440 66260 195492
rect 66312 195480 66318 195492
rect 68370 195480 68376 195492
rect 66312 195452 68376 195480
rect 66312 195440 66318 195452
rect 68370 195440 68376 195452
rect 68428 195440 68434 195492
rect 75270 195440 75276 195492
rect 75328 195480 75334 195492
rect 77938 195480 77944 195492
rect 75328 195452 77944 195480
rect 75328 195440 75334 195452
rect 77938 195440 77944 195452
rect 77996 195440 78002 195492
rect 376018 195168 376024 195220
rect 376076 195208 376082 195220
rect 379514 195208 379520 195220
rect 376076 195180 379520 195208
rect 376076 195168 376082 195180
rect 379514 195168 379520 195180
rect 379572 195168 379578 195220
rect 371234 194352 371240 194404
rect 371292 194392 371298 194404
rect 375282 194392 375288 194404
rect 371292 194364 375288 194392
rect 371292 194352 371298 194364
rect 375282 194352 375288 194364
rect 375340 194352 375346 194404
rect 217318 193808 217324 193860
rect 217376 193848 217382 193860
rect 580166 193848 580172 193860
rect 217376 193820 580172 193848
rect 217376 193808 217382 193820
rect 580166 193808 580172 193820
rect 580224 193808 580230 193860
rect 47578 193128 47584 193180
rect 47636 193168 47642 193180
rect 48958 193168 48964 193180
rect 47636 193140 48964 193168
rect 47636 193128 47642 193140
rect 48958 193128 48964 193140
rect 49016 193128 49022 193180
rect 371234 191876 371240 191888
rect 369872 191848 371240 191876
rect 365070 191768 365076 191820
rect 365128 191808 365134 191820
rect 369872 191808 369900 191848
rect 371234 191836 371240 191848
rect 371292 191836 371298 191888
rect 365128 191780 369900 191808
rect 365128 191768 365134 191780
rect 157334 189864 157340 189916
rect 157392 189864 157398 189916
rect 61378 188300 61384 188352
rect 61436 188340 61442 188352
rect 68922 188340 68928 188352
rect 61436 188312 68928 188340
rect 61436 188300 61442 188312
rect 68922 188300 68928 188312
rect 68980 188300 68986 188352
rect 71038 187892 71044 187944
rect 71096 187932 71102 187944
rect 73154 187932 73160 187944
rect 71096 187904 73160 187932
rect 71096 187892 71102 187904
rect 73154 187892 73160 187904
rect 73212 187892 73218 187944
rect 3142 187688 3148 187740
rect 3200 187728 3206 187740
rect 112438 187728 112444 187740
rect 3200 187700 112444 187728
rect 3200 187688 3206 187700
rect 112438 187688 112444 187700
rect 112496 187688 112502 187740
rect 166166 187620 166172 187672
rect 166224 187660 166230 187672
rect 399570 187660 399576 187672
rect 166224 187632 399576 187660
rect 166224 187620 166230 187632
rect 399570 187620 399576 187632
rect 399628 187620 399634 187672
rect 108298 186600 108304 186652
rect 108356 186640 108362 186652
rect 111058 186640 111064 186652
rect 108356 186612 111064 186640
rect 108356 186600 108362 186612
rect 111058 186600 111064 186612
rect 111116 186600 111122 186652
rect 45646 184832 45652 184884
rect 45704 184872 45710 184884
rect 53098 184872 53104 184884
rect 45704 184844 53104 184872
rect 45704 184832 45710 184844
rect 53098 184832 53104 184844
rect 53156 184832 53162 184884
rect 73154 184832 73160 184884
rect 73212 184872 73218 184884
rect 75178 184872 75184 184884
rect 73212 184844 75184 184872
rect 73212 184832 73218 184844
rect 75178 184832 75184 184844
rect 75236 184832 75242 184884
rect 142430 184260 142436 184272
rect 137986 184232 142436 184260
rect 135254 184152 135260 184204
rect 135312 184192 135318 184204
rect 137986 184192 138014 184232
rect 142430 184220 142436 184232
rect 142488 184220 142494 184272
rect 135312 184164 138014 184192
rect 135312 184152 135318 184164
rect 376110 182792 376116 182844
rect 376168 182832 376174 182844
rect 384298 182832 384304 182844
rect 376168 182804 384304 182832
rect 376168 182792 376174 182804
rect 384298 182792 384304 182804
rect 384356 182792 384362 182844
rect 68922 181432 68928 181484
rect 68980 181472 68986 181484
rect 83458 181472 83464 181484
rect 68980 181444 83464 181472
rect 68980 181432 68986 181444
rect 83458 181432 83464 181444
rect 83516 181432 83522 181484
rect 141234 180384 141240 180396
rect 137986 180356 141240 180384
rect 117314 180140 117320 180192
rect 117372 180180 117378 180192
rect 136358 180180 136364 180192
rect 117372 180152 136364 180180
rect 117372 180140 117378 180152
rect 136358 180140 136364 180152
rect 136416 180140 136422 180192
rect 53098 180072 53104 180124
rect 53156 180112 53162 180124
rect 63494 180112 63500 180124
rect 53156 180084 63500 180112
rect 53156 180072 53162 180084
rect 63494 180072 63500 180084
rect 63552 180072 63558 180124
rect 122098 180072 122104 180124
rect 122156 180112 122162 180124
rect 137986 180112 138014 180356
rect 141234 180344 141240 180356
rect 141292 180344 141298 180396
rect 122156 180084 138014 180112
rect 122156 180072 122162 180084
rect 77938 179392 77944 179444
rect 77996 179432 78002 179444
rect 79318 179432 79324 179444
rect 77996 179404 79324 179432
rect 77996 179392 78002 179404
rect 79318 179392 79324 179404
rect 79376 179392 79382 179444
rect 136358 178780 136364 178832
rect 136416 178820 136422 178832
rect 136726 178820 136732 178832
rect 136416 178792 136732 178820
rect 136416 178780 136422 178792
rect 136726 178780 136732 178792
rect 136784 178780 136790 178832
rect 120718 178644 120724 178696
rect 120776 178684 120782 178696
rect 136450 178684 136456 178696
rect 120776 178656 136456 178684
rect 120776 178644 120782 178656
rect 136450 178644 136456 178656
rect 136508 178644 136514 178696
rect 154390 178168 154396 178220
rect 154448 178208 154454 178220
rect 157794 178208 157800 178220
rect 154448 178180 157800 178208
rect 154448 178168 154454 178180
rect 157794 178168 157800 178180
rect 157852 178168 157858 178220
rect 75178 178100 75184 178152
rect 75236 178140 75242 178152
rect 77202 178140 77208 178152
rect 75236 178112 77208 178140
rect 75236 178100 75242 178112
rect 77202 178100 77208 178112
rect 77260 178100 77266 178152
rect 135990 178100 135996 178152
rect 136048 178140 136054 178152
rect 136542 178140 136548 178152
rect 136048 178112 136548 178140
rect 136048 178100 136054 178112
rect 136542 178100 136548 178112
rect 136600 178100 136606 178152
rect 48958 178032 48964 178084
rect 49016 178072 49022 178084
rect 49694 178072 49700 178084
rect 49016 178044 49700 178072
rect 49016 178032 49022 178044
rect 49694 178032 49700 178044
rect 49752 178032 49758 178084
rect 115750 178032 115756 178084
rect 115808 178072 115814 178084
rect 153930 178072 153936 178084
rect 115808 178044 153936 178072
rect 115808 178032 115814 178044
rect 153930 178032 153936 178044
rect 153988 178032 153994 178084
rect 158622 178032 158628 178084
rect 158680 178072 158686 178084
rect 579982 178072 579988 178084
rect 158680 178044 579988 178072
rect 158680 178032 158686 178044
rect 579982 178032 579988 178044
rect 580040 178032 580046 178084
rect 63494 177284 63500 177336
rect 63552 177324 63558 177336
rect 69750 177324 69756 177336
rect 63552 177296 69756 177324
rect 63552 177284 63558 177296
rect 69750 177284 69756 177296
rect 69808 177284 69814 177336
rect 120074 177284 120080 177336
rect 120132 177324 120138 177336
rect 135990 177324 135996 177336
rect 120132 177296 135996 177324
rect 120132 177284 120138 177296
rect 135990 177284 135996 177296
rect 136048 177284 136054 177336
rect 135714 176128 135720 176180
rect 135772 176168 135778 176180
rect 136542 176168 136548 176180
rect 135772 176140 136548 176168
rect 135772 176128 135778 176140
rect 136542 176128 136548 176140
rect 136600 176128 136606 176180
rect 122834 176060 122840 176112
rect 122892 176100 122898 176112
rect 136450 176100 136456 176112
rect 122892 176072 136456 176100
rect 122892 176060 122898 176072
rect 136450 176060 136456 176072
rect 136508 176060 136514 176112
rect 121454 175924 121460 175976
rect 121512 175964 121518 175976
rect 136358 175964 136364 175976
rect 121512 175936 136364 175964
rect 121512 175924 121518 175936
rect 136358 175924 136364 175936
rect 136416 175924 136422 175976
rect 149974 175516 149980 175568
rect 150032 175516 150038 175568
rect 144454 175448 144460 175500
rect 144512 175488 144518 175500
rect 149992 175488 150020 175516
rect 144512 175460 150020 175488
rect 144512 175448 144518 175460
rect 144086 175380 144092 175432
rect 144144 175420 144150 175432
rect 153930 175420 153936 175432
rect 144144 175392 153936 175420
rect 144144 175380 144150 175392
rect 153930 175380 153936 175392
rect 153988 175380 153994 175432
rect 77202 175244 77208 175296
rect 77260 175284 77266 175296
rect 77260 175256 77340 175284
rect 77260 175244 77266 175256
rect 77312 175216 77340 175256
rect 154390 175244 154396 175296
rect 154448 175284 154454 175296
rect 156506 175284 156512 175296
rect 154448 175256 156512 175284
rect 154448 175244 154454 175256
rect 156506 175244 156512 175256
rect 156564 175244 156570 175296
rect 78674 175216 78680 175228
rect 77312 175188 78680 175216
rect 78674 175176 78680 175188
rect 78732 175176 78738 175228
rect 141694 174700 141700 174752
rect 141752 174700 141758 174752
rect 141786 174700 141792 174752
rect 141844 174700 141850 174752
rect 125594 174496 125600 174548
rect 125652 174536 125658 174548
rect 135714 174536 135720 174548
rect 125652 174508 135720 174536
rect 125652 174496 125658 174508
rect 135714 174496 135720 174508
rect 135772 174496 135778 174548
rect 141712 174536 141740 174700
rect 141804 174604 141832 174700
rect 153470 174604 153476 174616
rect 141804 174576 153476 174604
rect 153470 174564 153476 174576
rect 153528 174564 153534 174616
rect 162486 174536 162492 174548
rect 141712 174508 162492 174536
rect 162486 174496 162492 174508
rect 162544 174496 162550 174548
rect 115658 174292 115664 174344
rect 115716 174332 115722 174344
rect 580442 174332 580448 174344
rect 115716 174304 580448 174332
rect 115716 174292 115722 174304
rect 580442 174292 580448 174304
rect 580500 174292 580506 174344
rect 129734 173884 129740 173936
rect 129792 173924 129798 173936
rect 137278 173924 137284 173936
rect 129792 173896 137284 173924
rect 129792 173884 129798 173896
rect 137278 173884 137284 173896
rect 137336 173884 137342 173936
rect 153470 173884 153476 173936
rect 153528 173924 153534 173936
rect 153528 173896 159496 173924
rect 153528 173884 153534 173896
rect 83458 173136 83464 173188
rect 83516 173176 83522 173188
rect 91554 173176 91560 173188
rect 83516 173148 91560 173176
rect 83516 173136 83522 173148
rect 91554 173136 91560 173148
rect 91612 173136 91618 173188
rect 126974 173136 126980 173188
rect 127032 173176 127038 173188
rect 136634 173176 136640 173188
rect 127032 173148 136640 173176
rect 127032 173136 127038 173148
rect 136634 173136 136640 173148
rect 136692 173136 136698 173188
rect 159468 173052 159496 173896
rect 161474 173136 161480 173188
rect 161532 173176 161538 173188
rect 166534 173176 166540 173188
rect 161532 173148 166540 173176
rect 161532 173136 161538 173148
rect 166534 173136 166540 173148
rect 166592 173136 166598 173188
rect 159450 173000 159456 173052
rect 159508 173000 159514 173052
rect 143442 172932 143448 172984
rect 143500 172972 143506 172984
rect 145650 172972 145656 172984
rect 143500 172944 145656 172972
rect 143500 172932 143506 172944
rect 145650 172932 145656 172944
rect 145708 172932 145714 172984
rect 146478 172932 146484 172984
rect 146536 172972 146542 172984
rect 148594 172972 148600 172984
rect 146536 172944 148600 172972
rect 146536 172932 146542 172944
rect 148594 172932 148600 172944
rect 148652 172932 148658 172984
rect 156506 172932 156512 172984
rect 156564 172972 156570 172984
rect 158438 172972 158444 172984
rect 156564 172944 158444 172972
rect 156564 172932 156570 172944
rect 158438 172932 158444 172944
rect 158496 172932 158502 172984
rect 143534 172864 143540 172916
rect 143592 172904 143598 172916
rect 146662 172904 146668 172916
rect 143592 172876 146668 172904
rect 143592 172864 143598 172876
rect 146662 172864 146668 172876
rect 146720 172864 146726 172916
rect 142430 172796 142436 172848
rect 142488 172836 142494 172848
rect 147582 172836 147588 172848
rect 142488 172808 147588 172836
rect 142488 172796 142494 172808
rect 147582 172796 147588 172808
rect 147640 172796 147646 172848
rect 49694 172456 49700 172508
rect 49752 172496 49758 172508
rect 53098 172496 53104 172508
rect 49752 172468 53104 172496
rect 49752 172456 49758 172468
rect 53098 172456 53104 172468
rect 53156 172456 53162 172508
rect 78674 172456 78680 172508
rect 78732 172496 78738 172508
rect 80606 172496 80612 172508
rect 78732 172468 80612 172496
rect 78732 172456 78738 172468
rect 80606 172456 80612 172468
rect 80664 172456 80670 172508
rect 133874 172116 133880 172168
rect 133932 172156 133938 172168
rect 140774 172156 140780 172168
rect 133932 172128 140780 172156
rect 133932 172116 133938 172128
rect 140774 172116 140780 172128
rect 140832 172116 140838 172168
rect 131114 171912 131120 171964
rect 131172 171952 131178 171964
rect 138658 171952 138664 171964
rect 131172 171924 138664 171952
rect 131172 171912 131178 171924
rect 138658 171912 138664 171924
rect 138716 171912 138722 171964
rect 140774 171776 140780 171828
rect 140832 171816 140838 171828
rect 144914 171816 144920 171828
rect 140832 171788 144920 171816
rect 140832 171776 140838 171788
rect 144914 171776 144920 171788
rect 144972 171776 144978 171828
rect 132494 171504 132500 171556
rect 132552 171544 132558 171556
rect 139670 171544 139676 171556
rect 132552 171516 139676 171544
rect 132552 171504 132558 171516
rect 139670 171504 139676 171516
rect 139728 171504 139734 171556
rect 128354 171096 128360 171148
rect 128412 171136 128418 171148
rect 136726 171136 136732 171148
rect 128412 171108 136732 171136
rect 128412 171096 128418 171108
rect 136726 171096 136732 171108
rect 136784 171096 136790 171148
rect 111058 170688 111064 170740
rect 111116 170728 111122 170740
rect 114462 170728 114468 170740
rect 111116 170700 114468 170728
rect 111116 170688 111122 170700
rect 114462 170688 114468 170700
rect 114520 170688 114526 170740
rect 45554 170348 45560 170400
rect 45612 170388 45618 170400
rect 63494 170388 63500 170400
rect 45612 170360 63500 170388
rect 45612 170348 45618 170360
rect 63494 170348 63500 170360
rect 63552 170348 63558 170400
rect 91554 170348 91560 170400
rect 91612 170388 91618 170400
rect 99374 170388 99380 170400
rect 91612 170360 99380 170388
rect 91612 170348 91618 170360
rect 99374 170348 99380 170360
rect 99432 170348 99438 170400
rect 358538 170348 358544 170400
rect 358596 170388 358602 170400
rect 376110 170388 376116 170400
rect 358596 170360 376116 170388
rect 358596 170348 358602 170360
rect 376110 170348 376116 170360
rect 376168 170348 376174 170400
rect 117406 169736 117412 169788
rect 117464 169776 117470 169788
rect 122098 169776 122104 169788
rect 117464 169748 122104 169776
rect 117464 169736 117470 169748
rect 122098 169736 122104 169748
rect 122156 169736 122162 169788
rect 362954 169056 362960 169108
rect 363012 169096 363018 169108
rect 364978 169096 364984 169108
rect 363012 169068 364984 169096
rect 363012 169056 363018 169068
rect 364978 169056 364984 169068
rect 365036 169056 365042 169108
rect 366358 168988 366364 169040
rect 366416 169028 366422 169040
rect 376018 169028 376024 169040
rect 366416 169000 376024 169028
rect 366416 168988 366422 169000
rect 376018 168988 376024 169000
rect 376076 168988 376082 169040
rect 79318 168716 79324 168768
rect 79376 168756 79382 168768
rect 81526 168756 81532 168768
rect 79376 168728 81532 168756
rect 79376 168716 79382 168728
rect 81526 168716 81532 168728
rect 81584 168716 81590 168768
rect 80606 168444 80612 168496
rect 80664 168484 80670 168496
rect 83458 168484 83464 168496
rect 80664 168456 83464 168484
rect 80664 168444 80670 168456
rect 83458 168444 83464 168456
rect 83516 168444 83522 168496
rect 114462 167628 114468 167680
rect 114520 167668 114526 167680
rect 138658 167668 138664 167680
rect 114520 167640 138664 167668
rect 114520 167628 114526 167640
rect 138658 167628 138664 167640
rect 138716 167628 138722 167680
rect 355318 167016 355324 167068
rect 355376 167056 355382 167068
rect 358538 167056 358544 167068
rect 355376 167028 358544 167056
rect 355376 167016 355382 167028
rect 358538 167016 358544 167028
rect 358596 167016 358602 167068
rect 68370 166404 68376 166456
rect 68428 166444 68434 166456
rect 69842 166444 69848 166456
rect 68428 166416 69848 166444
rect 68428 166404 68434 166416
rect 69842 166404 69848 166416
rect 69900 166404 69906 166456
rect 115106 166268 115112 166320
rect 115164 166308 115170 166320
rect 117406 166308 117412 166320
rect 115164 166280 117412 166308
rect 115164 166268 115170 166280
rect 117406 166268 117412 166280
rect 117464 166268 117470 166320
rect 185578 165588 185584 165640
rect 185636 165628 185642 165640
rect 579798 165628 579804 165640
rect 185636 165600 579804 165628
rect 185636 165588 185642 165600
rect 579798 165588 579804 165600
rect 579856 165588 579862 165640
rect 363598 165112 363604 165164
rect 363656 165152 363662 165164
rect 365070 165152 365076 165164
rect 363656 165124 365076 165152
rect 363656 165112 363662 165124
rect 365070 165112 365076 165124
rect 365128 165112 365134 165164
rect 81526 164160 81532 164212
rect 81584 164200 81590 164212
rect 83550 164200 83556 164212
rect 81584 164172 83556 164200
rect 81584 164160 81590 164172
rect 83550 164160 83556 164172
rect 83608 164160 83614 164212
rect 63494 163548 63500 163600
rect 63552 163588 63558 163600
rect 66254 163588 66260 163600
rect 63552 163560 66260 163588
rect 63552 163548 63558 163560
rect 66254 163548 66260 163560
rect 66312 163548 66318 163600
rect 99374 163480 99380 163532
rect 99432 163520 99438 163532
rect 113726 163520 113732 163532
rect 99432 163492 113732 163520
rect 99432 163480 99438 163492
rect 113726 163480 113732 163492
rect 113784 163480 113790 163532
rect 53098 162936 53104 162988
rect 53156 162976 53162 162988
rect 55858 162976 55864 162988
rect 53156 162948 55864 162976
rect 53156 162936 53162 162948
rect 55858 162936 55864 162948
rect 55916 162936 55922 162988
rect 3142 162868 3148 162920
rect 3200 162908 3206 162920
rect 175274 162908 175280 162920
rect 3200 162880 175280 162908
rect 3200 162868 3206 162880
rect 175274 162868 175280 162880
rect 175332 162868 175338 162920
rect 362954 162908 362960 162920
rect 361592 162880 362960 162908
rect 358446 162800 358452 162852
rect 358504 162840 358510 162852
rect 361592 162840 361620 162880
rect 362954 162868 362960 162880
rect 363012 162868 363018 162920
rect 358504 162812 361620 162840
rect 358504 162800 358510 162812
rect 66254 160692 66260 160744
rect 66312 160732 66318 160744
rect 79318 160732 79324 160744
rect 66312 160704 79324 160732
rect 66312 160692 66318 160704
rect 79318 160692 79324 160704
rect 79376 160692 79382 160744
rect 138658 160692 138664 160744
rect 138716 160732 138722 160744
rect 147674 160732 147680 160744
rect 138716 160704 147680 160732
rect 138716 160692 138722 160704
rect 147674 160692 147680 160704
rect 147732 160692 147738 160744
rect 69658 159196 69664 159248
rect 69716 159236 69722 159248
rect 71682 159236 71688 159248
rect 69716 159208 71688 159236
rect 69716 159196 69722 159208
rect 71682 159196 71688 159208
rect 71740 159196 71746 159248
rect 356054 157360 356060 157412
rect 356112 157400 356118 157412
rect 358446 157400 358452 157412
rect 356112 157372 358452 157400
rect 356112 157360 356118 157372
rect 358446 157360 358452 157372
rect 358504 157360 358510 157412
rect 79318 157292 79324 157344
rect 79376 157332 79382 157344
rect 85298 157332 85304 157344
rect 79376 157304 85304 157332
rect 79376 157292 79382 157304
rect 85298 157292 85304 157304
rect 85356 157292 85362 157344
rect 352558 157292 352564 157344
rect 352616 157332 352622 157344
rect 355318 157332 355324 157344
rect 352616 157304 355324 157332
rect 352616 157292 352622 157304
rect 355318 157292 355324 157304
rect 355376 157292 355382 157344
rect 69842 154504 69848 154556
rect 69900 154544 69906 154556
rect 71222 154544 71228 154556
rect 69900 154516 71228 154544
rect 69900 154504 69906 154516
rect 71222 154504 71228 154516
rect 71280 154504 71286 154556
rect 85298 154504 85304 154556
rect 85356 154544 85362 154556
rect 87598 154544 87604 154556
rect 85356 154516 87604 154544
rect 85356 154504 85362 154516
rect 87598 154504 87604 154516
rect 87656 154504 87662 154556
rect 147674 153824 147680 153876
rect 147732 153864 147738 153876
rect 159358 153864 159364 153876
rect 147732 153836 159364 153864
rect 147732 153824 147738 153836
rect 159358 153824 159364 153836
rect 159416 153824 159422 153876
rect 71774 153620 71780 153672
rect 71832 153660 71838 153672
rect 75914 153660 75920 153672
rect 71832 153632 75920 153660
rect 71832 153620 71838 153632
rect 75914 153620 75920 153632
rect 75972 153620 75978 153672
rect 356054 153252 356060 153264
rect 354646 153224 356060 153252
rect 147490 153144 147496 153196
rect 147548 153184 147554 153196
rect 149238 153184 149244 153196
rect 147548 153156 149244 153184
rect 147548 153144 147554 153156
rect 149238 153144 149244 153156
rect 149296 153144 149302 153196
rect 349798 153144 349804 153196
rect 349856 153184 349862 153196
rect 354646 153184 354674 153224
rect 356054 153212 356060 153224
rect 356112 153212 356118 153264
rect 349856 153156 354674 153184
rect 349856 153144 349862 153156
rect 343634 151036 343640 151088
rect 343692 151076 343698 151088
rect 349798 151076 349804 151088
rect 343692 151048 349804 151076
rect 343692 151036 343698 151048
rect 349798 151036 349804 151048
rect 349856 151036 349862 151088
rect 69750 150900 69756 150952
rect 69808 150940 69814 150952
rect 72142 150940 72148 150952
rect 69808 150912 72148 150940
rect 69808 150900 69814 150912
rect 72142 150900 72148 150912
rect 72200 150900 72206 150952
rect 71222 150424 71228 150476
rect 71280 150464 71286 150476
rect 72418 150464 72424 150476
rect 71280 150436 72424 150464
rect 71280 150424 71286 150436
rect 72418 150424 72424 150436
rect 72476 150424 72482 150476
rect 159358 149744 159364 149796
rect 159416 149784 159422 149796
rect 166258 149784 166264 149796
rect 159416 149756 166264 149784
rect 159416 149744 159422 149756
rect 166258 149744 166264 149756
rect 166316 149744 166322 149796
rect 115566 149676 115572 149728
rect 115624 149716 115630 149728
rect 580534 149716 580540 149728
rect 115624 149688 580540 149716
rect 115624 149676 115630 149688
rect 580534 149676 580540 149688
rect 580592 149676 580598 149728
rect 3142 149064 3148 149116
rect 3200 149104 3206 149116
rect 25498 149104 25504 149116
rect 3200 149076 25504 149104
rect 3200 149064 3206 149076
rect 25498 149064 25504 149076
rect 25556 149064 25562 149116
rect 363690 148792 363696 148844
rect 363748 148832 363754 148844
rect 366358 148832 366364 148844
rect 363748 148804 366364 148832
rect 363748 148792 363754 148804
rect 366358 148792 366364 148804
rect 366416 148792 366422 148844
rect 83458 148316 83464 148368
rect 83516 148356 83522 148368
rect 88242 148356 88248 148368
rect 83516 148328 88248 148356
rect 83516 148316 83522 148328
rect 88242 148316 88248 148328
rect 88300 148316 88306 148368
rect 149238 148316 149244 148368
rect 149296 148356 149302 148368
rect 155218 148356 155224 148368
rect 149296 148328 155224 148356
rect 149296 148316 149302 148328
rect 155218 148316 155224 148328
rect 155276 148316 155282 148368
rect 83550 147636 83556 147688
rect 83608 147676 83614 147688
rect 83608 147648 84194 147676
rect 83608 147636 83614 147648
rect 84166 147608 84194 147648
rect 171778 147636 171784 147688
rect 171836 147676 171842 147688
rect 173158 147676 173164 147688
rect 171836 147648 173164 147676
rect 171836 147636 171842 147648
rect 173158 147636 173164 147648
rect 173216 147636 173222 147688
rect 341518 147636 341524 147688
rect 341576 147676 341582 147688
rect 343634 147676 343640 147688
rect 341576 147648 343640 147676
rect 341576 147636 341582 147648
rect 343634 147636 343640 147648
rect 343692 147636 343698 147688
rect 86218 147608 86224 147620
rect 84166 147580 86224 147608
rect 86218 147568 86224 147580
rect 86276 147568 86282 147620
rect 351178 146888 351184 146940
rect 351236 146928 351242 146940
rect 363598 146928 363604 146940
rect 351236 146900 363604 146928
rect 351236 146888 351242 146900
rect 363598 146888 363604 146900
rect 363656 146888 363662 146940
rect 75914 146276 75920 146328
rect 75972 146316 75978 146328
rect 75972 146288 77340 146316
rect 75972 146276 75978 146288
rect 77312 146248 77340 146288
rect 80698 146248 80704 146260
rect 77312 146220 80704 146248
rect 80698 146208 80704 146220
rect 80756 146208 80762 146260
rect 88334 144848 88340 144900
rect 88392 144888 88398 144900
rect 89990 144888 89996 144900
rect 88392 144860 89996 144888
rect 88392 144848 88398 144860
rect 89990 144848 89996 144860
rect 90048 144848 90054 144900
rect 115474 144168 115480 144220
rect 115532 144208 115538 144220
rect 580626 144208 580632 144220
rect 115532 144180 580632 144208
rect 115532 144168 115538 144180
rect 580626 144168 580632 144180
rect 580684 144168 580690 144220
rect 72142 142808 72148 142860
rect 72200 142848 72206 142860
rect 91738 142848 91744 142860
rect 72200 142820 91744 142848
rect 72200 142808 72206 142820
rect 91738 142808 91744 142820
rect 91796 142808 91802 142860
rect 115934 142808 115940 142860
rect 115992 142848 115998 142860
rect 477494 142848 477500 142860
rect 115992 142820 477500 142848
rect 115992 142808 115998 142820
rect 477494 142808 477500 142820
rect 477552 142808 477558 142860
rect 89990 141380 89996 141432
rect 90048 141420 90054 141432
rect 97994 141420 98000 141432
rect 90048 141392 98000 141420
rect 90048 141380 90054 141392
rect 97994 141380 98000 141392
rect 98052 141380 98058 141432
rect 86218 141108 86224 141160
rect 86276 141148 86282 141160
rect 91094 141148 91100 141160
rect 86276 141120 91100 141148
rect 86276 141108 86282 141120
rect 91094 141108 91100 141120
rect 91152 141108 91158 141160
rect 166258 141108 166264 141160
rect 166316 141148 166322 141160
rect 169754 141148 169760 141160
rect 166316 141120 169760 141148
rect 166316 141108 166322 141120
rect 169754 141108 169760 141120
rect 169812 141108 169818 141160
rect 68278 140768 68284 140820
rect 68336 140808 68342 140820
rect 68336 140780 69060 140808
rect 68336 140768 68342 140780
rect 69032 140740 69060 140780
rect 71406 140740 71412 140752
rect 69032 140712 71412 140740
rect 71406 140700 71412 140712
rect 71464 140700 71470 140752
rect 173158 140292 173164 140344
rect 173216 140332 173222 140344
rect 177298 140332 177304 140344
rect 173216 140304 177304 140332
rect 173216 140292 173222 140304
rect 177298 140292 177304 140304
rect 177356 140292 177362 140344
rect 87598 139884 87604 139936
rect 87656 139924 87662 139936
rect 89898 139924 89904 139936
rect 87656 139896 89904 139924
rect 87656 139884 87662 139896
rect 89898 139884 89904 139896
rect 89956 139884 89962 139936
rect 347038 139408 347044 139460
rect 347096 139448 347102 139460
rect 351178 139448 351184 139460
rect 347096 139420 351184 139448
rect 347096 139408 347102 139420
rect 351178 139408 351184 139420
rect 351236 139408 351242 139460
rect 91738 138660 91744 138712
rect 91796 138700 91802 138712
rect 97166 138700 97172 138712
rect 91796 138672 97172 138700
rect 91796 138660 91802 138672
rect 97166 138660 97172 138672
rect 97224 138660 97230 138712
rect 55858 138524 55864 138576
rect 55916 138564 55922 138576
rect 57882 138564 57888 138576
rect 55916 138536 57888 138564
rect 55916 138524 55922 138536
rect 57882 138524 57888 138536
rect 57940 138524 57946 138576
rect 3418 138320 3424 138372
rect 3476 138360 3482 138372
rect 4062 138360 4068 138372
rect 3476 138332 4068 138360
rect 3476 138320 3482 138332
rect 4062 138320 4068 138332
rect 4120 138320 4126 138372
rect 71406 137980 71412 138032
rect 71464 138020 71470 138032
rect 71464 137992 71820 138020
rect 71464 137980 71470 137992
rect 71792 137952 71820 137992
rect 80698 137980 80704 138032
rect 80756 138020 80762 138032
rect 80756 137992 81480 138020
rect 80756 137980 80762 137992
rect 73154 137952 73160 137964
rect 71792 137924 73160 137952
rect 73154 137912 73160 137924
rect 73212 137912 73218 137964
rect 81452 137952 81480 137992
rect 114462 137980 114468 138032
rect 114520 138020 114526 138032
rect 579614 138020 579620 138032
rect 114520 137992 579620 138020
rect 114520 137980 114526 137992
rect 579614 137980 579620 137992
rect 579672 137980 579678 138032
rect 86218 137952 86224 137964
rect 81452 137924 86224 137952
rect 86218 137912 86224 137924
rect 86276 137912 86282 137964
rect 119338 137912 119344 137964
rect 119396 137952 119402 137964
rect 120718 137952 120724 137964
rect 119396 137924 120724 137952
rect 119396 137912 119402 137924
rect 120718 137912 120724 137924
rect 120776 137912 120782 137964
rect 150526 137912 150532 137964
rect 150584 137952 150590 137964
rect 152182 137952 152188 137964
rect 150584 137924 152188 137952
rect 150584 137912 150590 137924
rect 152182 137912 152188 137924
rect 152240 137912 152246 137964
rect 152458 137912 152464 137964
rect 152516 137952 152522 137964
rect 153746 137952 153752 137964
rect 152516 137924 153752 137952
rect 152516 137912 152522 137924
rect 153746 137912 153752 137924
rect 153804 137912 153810 137964
rect 164510 137912 164516 137964
rect 164568 137952 164574 137964
rect 172514 137952 172520 137964
rect 164568 137924 172520 137952
rect 164568 137912 164574 137924
rect 172514 137912 172520 137924
rect 172572 137912 172578 137964
rect 155218 137640 155224 137692
rect 155276 137680 155282 137692
rect 164694 137680 164700 137692
rect 155276 137652 164700 137680
rect 155276 137640 155282 137652
rect 164694 137640 164700 137652
rect 164752 137640 164758 137692
rect 144454 137572 144460 137624
rect 144512 137612 144518 137624
rect 156874 137612 156880 137624
rect 144512 137584 156880 137612
rect 144512 137572 144518 137584
rect 156874 137572 156880 137584
rect 156932 137572 156938 137624
rect 163498 137572 163504 137624
rect 163556 137612 163562 137624
rect 174078 137612 174084 137624
rect 163556 137584 174084 137612
rect 163556 137572 163562 137584
rect 174078 137572 174084 137584
rect 174136 137572 174142 137624
rect 342254 137572 342260 137624
rect 342312 137612 342318 137624
rect 352558 137612 352564 137624
rect 342312 137584 352564 137612
rect 342312 137572 342318 137584
rect 352558 137572 352564 137584
rect 352616 137572 352622 137624
rect 114186 137504 114192 137556
rect 114244 137544 114250 137556
rect 396902 137544 396908 137556
rect 114244 137516 396908 137544
rect 114244 137504 114250 137516
rect 396902 137504 396908 137516
rect 396960 137504 396966 137556
rect 114278 137436 114284 137488
rect 114336 137476 114342 137488
rect 397086 137476 397092 137488
rect 114336 137448 397092 137476
rect 114336 137436 114342 137448
rect 397086 137436 397092 137448
rect 397144 137436 397150 137488
rect 114370 137368 114376 137420
rect 114428 137408 114434 137420
rect 397178 137408 397184 137420
rect 114428 137380 397184 137408
rect 114428 137368 114434 137380
rect 397178 137368 397184 137380
rect 397236 137368 397242 137420
rect 114094 137300 114100 137352
rect 114152 137340 114158 137352
rect 398098 137340 398104 137352
rect 114152 137312 398104 137340
rect 114152 137300 114158 137312
rect 398098 137300 398104 137312
rect 398156 137300 398162 137352
rect 113910 137232 113916 137284
rect 113968 137272 113974 137284
rect 542354 137272 542360 137284
rect 113968 137244 542360 137272
rect 113968 137232 113974 137244
rect 542354 137232 542360 137244
rect 542412 137232 542418 137284
rect 142430 137028 142436 137080
rect 142488 137068 142494 137080
rect 145926 137068 145932 137080
rect 142488 137040 145932 137068
rect 142488 137028 142494 137040
rect 145926 137028 145932 137040
rect 145984 137028 145990 137080
rect 163590 136824 163596 136876
rect 163648 136864 163654 136876
rect 170950 136864 170956 136876
rect 163648 136836 170956 136864
rect 163648 136824 163654 136836
rect 170950 136824 170956 136836
rect 171008 136824 171014 136876
rect 138106 136756 138112 136808
rect 138164 136796 138170 136808
rect 142522 136796 142528 136808
rect 138164 136768 142528 136796
rect 138164 136756 138170 136768
rect 142522 136756 142528 136768
rect 142580 136756 142586 136808
rect 153470 136756 153476 136808
rect 153528 136796 153534 136808
rect 155310 136796 155316 136808
rect 153528 136768 155316 136796
rect 153528 136756 153534 136768
rect 155310 136756 155316 136768
rect 155368 136756 155374 136808
rect 3418 136620 3424 136672
rect 3476 136660 3482 136672
rect 115198 136660 115204 136672
rect 3476 136632 115204 136660
rect 3476 136620 3482 136632
rect 115198 136620 115204 136632
rect 115256 136620 115262 136672
rect 72418 136552 72424 136604
rect 72476 136592 72482 136604
rect 73798 136592 73804 136604
rect 72476 136564 73804 136592
rect 72476 136552 72482 136564
rect 73798 136552 73804 136564
rect 73856 136552 73862 136604
rect 89898 136552 89904 136604
rect 89956 136592 89962 136604
rect 95878 136592 95884 136604
rect 89956 136564 95884 136592
rect 89956 136552 89962 136564
rect 95878 136552 95884 136564
rect 95936 136552 95942 136604
rect 113726 136552 113732 136604
rect 113784 136592 113790 136604
rect 116578 136592 116584 136604
rect 113784 136564 116584 136592
rect 113784 136552 113790 136564
rect 116578 136552 116584 136564
rect 116636 136552 116642 136604
rect 73154 136484 73160 136536
rect 73212 136524 73218 136536
rect 75178 136524 75184 136536
rect 73212 136496 75184 136524
rect 73212 136484 73218 136496
rect 75178 136484 75184 136496
rect 75236 136484 75242 136536
rect 169754 136484 169760 136536
rect 169812 136524 169818 136536
rect 175918 136524 175924 136536
rect 169812 136496 175924 136524
rect 169812 136484 169818 136496
rect 175918 136484 175924 136496
rect 175976 136484 175982 136536
rect 40034 136416 40040 136468
rect 40092 136456 40098 136468
rect 175458 136456 175464 136468
rect 40092 136428 175464 136456
rect 40092 136416 40098 136428
rect 175458 136416 175464 136428
rect 175516 136416 175522 136468
rect 3970 136348 3976 136400
rect 4028 136388 4034 136400
rect 178770 136388 178776 136400
rect 4028 136360 178776 136388
rect 4028 136348 4034 136360
rect 178770 136348 178776 136360
rect 178828 136348 178834 136400
rect 3786 136280 3792 136332
rect 3844 136320 3850 136332
rect 178034 136320 178040 136332
rect 3844 136292 178040 136320
rect 3844 136280 3850 136292
rect 178034 136280 178040 136292
rect 178092 136280 178098 136332
rect 360838 136280 360844 136332
rect 360896 136320 360902 136332
rect 363690 136320 363696 136332
rect 360896 136292 363696 136320
rect 360896 136280 360902 136292
rect 363690 136280 363696 136292
rect 363748 136280 363754 136332
rect 3878 136212 3884 136264
rect 3936 136252 3942 136264
rect 178402 136252 178408 136264
rect 3936 136224 178408 136252
rect 3936 136212 3942 136224
rect 178402 136212 178408 136224
rect 178460 136212 178466 136264
rect 3694 136144 3700 136196
rect 3752 136184 3758 136196
rect 178678 136184 178684 136196
rect 3752 136156 178684 136184
rect 3752 136144 3758 136156
rect 178678 136144 178684 136156
rect 178736 136144 178742 136196
rect 3234 136076 3240 136128
rect 3292 136116 3298 136128
rect 178862 136116 178868 136128
rect 3292 136088 178868 136116
rect 3292 136076 3298 136088
rect 178862 136076 178868 136088
rect 178920 136076 178926 136128
rect 3326 136008 3332 136060
rect 3384 136048 3390 136060
rect 178494 136048 178500 136060
rect 3384 136020 178500 136048
rect 3384 136008 3390 136020
rect 178494 136008 178500 136020
rect 178552 136008 178558 136060
rect 113818 135940 113824 135992
rect 113876 135980 113882 135992
rect 412634 135980 412640 135992
rect 113876 135952 412640 135980
rect 113876 135940 113882 135952
rect 412634 135940 412640 135952
rect 412692 135940 412698 135992
rect 115382 135872 115388 135924
rect 115440 135912 115446 135924
rect 580810 135912 580816 135924
rect 115440 135884 580816 135912
rect 115440 135872 115446 135884
rect 580810 135872 580816 135884
rect 580868 135872 580874 135924
rect 97166 135192 97172 135244
rect 97224 135232 97230 135244
rect 102778 135232 102784 135244
rect 97224 135204 102784 135232
rect 97224 135192 97230 135204
rect 102778 135192 102784 135204
rect 102836 135192 102842 135244
rect 57882 134716 57888 134768
rect 57940 134756 57946 134768
rect 176562 134756 176568 134768
rect 57940 134728 176568 134756
rect 57940 134716 57946 134728
rect 176562 134716 176568 134728
rect 176620 134716 176626 134768
rect 3602 134648 3608 134700
rect 3660 134688 3666 134700
rect 178310 134688 178316 134700
rect 3660 134660 178316 134688
rect 3660 134648 3666 134660
rect 178310 134648 178316 134660
rect 178368 134648 178374 134700
rect 4062 134580 4068 134632
rect 4120 134620 4126 134632
rect 178126 134620 178132 134632
rect 4120 134592 178132 134620
rect 4120 134580 4126 134592
rect 178126 134580 178132 134592
rect 178184 134580 178190 134632
rect 115290 134512 115296 134564
rect 115348 134552 115354 134564
rect 342254 134552 342260 134564
rect 115348 134524 342260 134552
rect 115348 134512 115354 134524
rect 342254 134512 342260 134524
rect 342312 134512 342318 134564
rect 3786 133900 3792 133952
rect 3844 133940 3850 133952
rect 175366 133940 175372 133952
rect 3844 133912 175372 133940
rect 3844 133900 3850 133912
rect 175366 133900 175372 133912
rect 175424 133900 175430 133952
rect 97994 133832 98000 133884
rect 98052 133872 98058 133884
rect 101398 133872 101404 133884
rect 98052 133844 101404 133872
rect 98052 133832 98058 133844
rect 101398 133832 101404 133844
rect 101456 133832 101462 133884
rect 91094 133084 91100 133136
rect 91152 133124 91158 133136
rect 93854 133124 93860 133136
rect 91152 133096 93860 133124
rect 91152 133084 91158 133096
rect 93854 133084 93860 133096
rect 93912 133084 93918 133136
rect 3418 131112 3424 131164
rect 3476 131152 3482 131164
rect 113726 131152 113732 131164
rect 3476 131124 113732 131152
rect 3476 131112 3482 131124
rect 113726 131112 113732 131124
rect 113784 131112 113790 131164
rect 345658 131112 345664 131164
rect 345716 131152 345722 131164
rect 347038 131152 347044 131164
rect 345716 131124 347044 131152
rect 345716 131112 345722 131124
rect 347038 131112 347044 131124
rect 347096 131112 347102 131164
rect 95878 130364 95884 130416
rect 95936 130404 95942 130416
rect 108298 130404 108304 130416
rect 95936 130376 108304 130404
rect 95936 130364 95942 130376
rect 108298 130364 108304 130376
rect 108356 130364 108362 130416
rect 93854 128596 93860 128648
rect 93912 128636 93918 128648
rect 97258 128636 97264 128648
rect 93912 128608 97264 128636
rect 93912 128596 93918 128608
rect 97258 128596 97264 128608
rect 97316 128596 97322 128648
rect 3602 128324 3608 128376
rect 3660 128364 3666 128376
rect 113726 128364 113732 128376
rect 3660 128336 113732 128364
rect 3660 128324 3666 128336
rect 113726 128324 113732 128336
rect 113784 128324 113790 128376
rect 73798 127576 73804 127628
rect 73856 127616 73862 127628
rect 82078 127616 82084 127628
rect 73856 127588 82084 127616
rect 73856 127576 73862 127588
rect 82078 127576 82084 127588
rect 82136 127576 82142 127628
rect 3694 126964 3700 127016
rect 3752 127004 3758 127016
rect 113634 127004 113640 127016
rect 3752 126976 113640 127004
rect 3752 126964 3758 126976
rect 113634 126964 113640 126976
rect 113692 126964 113698 127016
rect 25498 126896 25504 126948
rect 25556 126936 25562 126948
rect 113726 126936 113732 126948
rect 25556 126908 113732 126936
rect 25556 126896 25562 126908
rect 113726 126896 113732 126908
rect 113784 126896 113790 126948
rect 86218 126828 86224 126880
rect 86276 126868 86282 126880
rect 88334 126868 88340 126880
rect 86276 126840 88340 126868
rect 86276 126828 86282 126840
rect 88334 126828 88340 126840
rect 88392 126828 88398 126880
rect 184198 125604 184204 125656
rect 184256 125644 184262 125656
rect 579706 125644 579712 125656
rect 184256 125616 579712 125644
rect 184256 125604 184262 125616
rect 579706 125604 579712 125616
rect 579764 125604 579770 125656
rect 22830 125536 22836 125588
rect 22888 125576 22894 125588
rect 113542 125576 113548 125588
rect 22888 125548 113548 125576
rect 22888 125536 22894 125548
rect 113542 125536 113548 125548
rect 113600 125536 113606 125588
rect 88334 125468 88340 125520
rect 88392 125508 88398 125520
rect 90358 125508 90364 125520
rect 88392 125480 90364 125508
rect 88392 125468 88398 125480
rect 90358 125468 90364 125480
rect 90416 125468 90422 125520
rect 344278 124176 344284 124228
rect 344336 124216 344342 124228
rect 345658 124216 345664 124228
rect 344336 124188 345664 124216
rect 344336 124176 344342 124188
rect 345658 124176 345664 124188
rect 345716 124176 345722 124228
rect 22738 124108 22744 124160
rect 22796 124148 22802 124160
rect 113726 124148 113732 124160
rect 22796 124120 113732 124148
rect 22796 124108 22802 124120
rect 113726 124108 113732 124120
rect 113784 124108 113790 124160
rect 175918 124108 175924 124160
rect 175976 124148 175982 124160
rect 178218 124148 178224 124160
rect 175976 124120 178224 124148
rect 175976 124108 175982 124120
rect 178218 124108 178224 124120
rect 178276 124108 178282 124160
rect 358078 124108 358084 124160
rect 358136 124148 358142 124160
rect 360838 124148 360844 124160
rect 358136 124120 360844 124148
rect 358136 124108 358142 124120
rect 360838 124108 360844 124120
rect 360896 124108 360902 124160
rect 24118 122748 24124 122800
rect 24176 122788 24182 122800
rect 113358 122788 113364 122800
rect 24176 122760 113364 122788
rect 24176 122748 24182 122760
rect 113358 122748 113364 122760
rect 113416 122748 113422 122800
rect 97258 121796 97264 121848
rect 97316 121836 97322 121848
rect 98730 121836 98736 121848
rect 97316 121808 98736 121836
rect 97316 121796 97322 121808
rect 98730 121796 98736 121808
rect 98788 121796 98794 121848
rect 10318 121388 10324 121440
rect 10376 121428 10382 121440
rect 113726 121428 113732 121440
rect 10376 121400 113732 121428
rect 10376 121388 10382 121400
rect 113726 121388 113732 121400
rect 113784 121388 113790 121440
rect 82078 121320 82084 121372
rect 82136 121360 82142 121372
rect 85850 121360 85856 121372
rect 82136 121332 85856 121360
rect 82136 121320 82142 121332
rect 85850 121320 85856 121332
rect 85908 121320 85914 121372
rect 98730 121320 98736 121372
rect 98788 121360 98794 121372
rect 100018 121360 100024 121372
rect 98788 121332 100024 121360
rect 98788 121320 98794 121332
rect 100018 121320 100024 121332
rect 100076 121320 100082 121372
rect 8938 120028 8944 120080
rect 8996 120068 9002 120080
rect 113726 120068 113732 120080
rect 8996 120040 113732 120068
rect 8996 120028 9002 120040
rect 113726 120028 113732 120040
rect 113784 120028 113790 120080
rect 5074 118600 5080 118652
rect 5132 118640 5138 118652
rect 113634 118640 113640 118652
rect 5132 118612 113640 118640
rect 5132 118600 5138 118612
rect 113634 118600 113640 118612
rect 113692 118600 113698 118652
rect 85850 117376 85856 117428
rect 85908 117416 85914 117428
rect 87598 117416 87604 117428
rect 85908 117388 87604 117416
rect 85908 117376 85914 117388
rect 87598 117376 87604 117388
rect 87656 117376 87662 117428
rect 42058 117240 42064 117292
rect 42116 117280 42122 117292
rect 113726 117280 113732 117292
rect 42116 117252 113732 117280
rect 42116 117240 42122 117252
rect 113726 117240 113732 117252
rect 113784 117240 113790 117292
rect 338758 117240 338764 117292
rect 338816 117280 338822 117292
rect 341518 117280 341524 117292
rect 338816 117252 341524 117280
rect 338816 117240 338822 117252
rect 341518 117240 341524 117252
rect 341576 117240 341582 117292
rect 19978 115880 19984 115932
rect 20036 115920 20042 115932
rect 113726 115920 113732 115932
rect 20036 115892 113732 115920
rect 20036 115880 20042 115892
rect 113726 115880 113732 115892
rect 113784 115880 113790 115932
rect 177298 115880 177304 115932
rect 177356 115920 177362 115932
rect 178034 115920 178040 115932
rect 177356 115892 178040 115920
rect 177356 115880 177362 115892
rect 178034 115880 178040 115892
rect 178092 115880 178098 115932
rect 90358 115812 90364 115864
rect 90416 115852 90422 115864
rect 93486 115852 93492 115864
rect 90416 115824 93492 115852
rect 90416 115812 90422 115824
rect 93486 115812 93492 115824
rect 93544 115812 93550 115864
rect 37918 113092 37924 113144
rect 37976 113132 37982 113144
rect 113726 113132 113732 113144
rect 37976 113104 113732 113132
rect 37976 113092 37982 113104
rect 113726 113092 113732 113104
rect 113784 113092 113790 113144
rect 15838 111732 15844 111784
rect 15896 111772 15902 111784
rect 113726 111772 113732 111784
rect 15896 111744 113732 111772
rect 15896 111732 15902 111744
rect 113726 111732 113732 111744
rect 113784 111732 113790 111784
rect 93486 111664 93492 111716
rect 93544 111704 93550 111716
rect 96522 111704 96528 111716
rect 93544 111676 96528 111704
rect 93544 111664 93550 111676
rect 96522 111664 96528 111676
rect 96580 111664 96586 111716
rect 348418 111052 348424 111104
rect 348476 111092 348482 111104
rect 358078 111092 358084 111104
rect 348476 111064 358084 111092
rect 348476 111052 348482 111064
rect 358078 111052 358084 111064
rect 358136 111052 358142 111104
rect 87598 110916 87604 110968
rect 87656 110956 87662 110968
rect 88702 110956 88708 110968
rect 87656 110928 88708 110956
rect 87656 110916 87662 110928
rect 88702 110916 88708 110928
rect 88760 110916 88766 110968
rect 75178 110508 75184 110560
rect 75236 110548 75242 110560
rect 77938 110548 77944 110560
rect 75236 110520 77944 110548
rect 75236 110508 75242 110520
rect 77938 110508 77944 110520
rect 77996 110508 78002 110560
rect 23474 110372 23480 110424
rect 23532 110412 23538 110424
rect 113726 110412 113732 110424
rect 23532 110384 113732 110412
rect 23532 110372 23538 110384
rect 113726 110372 113732 110384
rect 113784 110372 113790 110424
rect 101398 109216 101404 109268
rect 101456 109256 101462 109268
rect 102134 109256 102140 109268
rect 101456 109228 102140 109256
rect 101456 109216 101462 109228
rect 102134 109216 102140 109228
rect 102192 109216 102198 109268
rect 100018 108944 100024 108996
rect 100076 108984 100082 108996
rect 102226 108984 102232 108996
rect 100076 108956 102232 108984
rect 100076 108944 100082 108956
rect 102226 108944 102232 108956
rect 102284 108944 102290 108996
rect 108298 108944 108304 108996
rect 108356 108984 108362 108996
rect 113726 108984 113732 108996
rect 108356 108956 113732 108984
rect 108356 108944 108362 108956
rect 113726 108944 113732 108956
rect 113784 108944 113790 108996
rect 96522 108604 96528 108656
rect 96580 108644 96586 108656
rect 97902 108644 97908 108656
rect 96580 108616 97908 108644
rect 96580 108604 96586 108616
rect 97902 108604 97908 108616
rect 97960 108604 97966 108656
rect 88702 107584 88708 107636
rect 88760 107624 88766 107636
rect 113542 107624 113548 107636
rect 88760 107596 113548 107624
rect 88760 107584 88766 107596
rect 113542 107584 113548 107596
rect 113600 107584 113606 107636
rect 337010 106768 337016 106820
rect 337068 106808 337074 106820
rect 338758 106808 338764 106820
rect 337068 106780 338764 106808
rect 337068 106768 337074 106780
rect 338758 106768 338764 106780
rect 338816 106768 338822 106820
rect 102226 106224 102232 106276
rect 102284 106264 102290 106276
rect 113726 106264 113732 106276
rect 102284 106236 113732 106264
rect 102284 106224 102290 106236
rect 113726 106224 113732 106236
rect 113784 106224 113790 106276
rect 178034 106224 178040 106276
rect 178092 106264 178098 106276
rect 344278 106264 344284 106276
rect 178092 106236 344284 106264
rect 178092 106224 178098 106236
rect 344278 106224 344284 106236
rect 344336 106224 344342 106276
rect 102134 105204 102140 105256
rect 102192 105244 102198 105256
rect 104618 105244 104624 105256
rect 102192 105216 104624 105244
rect 102192 105204 102198 105216
rect 104618 105204 104624 105216
rect 104676 105204 104682 105256
rect 97994 104796 98000 104848
rect 98052 104836 98058 104848
rect 113358 104836 113364 104848
rect 98052 104808 113364 104836
rect 98052 104796 98058 104808
rect 113358 104796 113364 104808
rect 113416 104796 113422 104848
rect 178034 104796 178040 104848
rect 178092 104836 178098 104848
rect 337010 104836 337016 104848
rect 178092 104808 337016 104836
rect 178092 104796 178098 104808
rect 337010 104796 337016 104808
rect 337068 104796 337074 104848
rect 178034 103436 178040 103488
rect 178092 103476 178098 103488
rect 413278 103476 413284 103488
rect 178092 103448 413284 103476
rect 178092 103436 178098 103448
rect 413278 103436 413284 103448
rect 413336 103436 413342 103488
rect 178034 102076 178040 102128
rect 178092 102116 178098 102128
rect 410518 102116 410524 102128
rect 178092 102088 410524 102116
rect 178092 102076 178098 102088
rect 410518 102076 410524 102088
rect 410576 102076 410582 102128
rect 178034 100648 178040 100700
rect 178092 100688 178098 100700
rect 409138 100688 409144 100700
rect 178092 100660 409144 100688
rect 178092 100648 178098 100660
rect 409138 100648 409144 100660
rect 409196 100648 409202 100700
rect 175918 99356 175924 99408
rect 175976 99396 175982 99408
rect 580166 99396 580172 99408
rect 175976 99368 580172 99396
rect 175976 99356 175982 99368
rect 580166 99356 580172 99368
rect 580224 99356 580230 99408
rect 178034 99288 178040 99340
rect 178092 99328 178098 99340
rect 407758 99328 407764 99340
rect 178092 99300 407764 99328
rect 178092 99288 178098 99300
rect 407758 99288 407764 99300
rect 407816 99288 407822 99340
rect 104618 98948 104624 99000
rect 104676 98988 104682 99000
rect 106550 98988 106556 99000
rect 104676 98960 106556 98988
rect 104676 98948 104682 98960
rect 106550 98948 106556 98960
rect 106608 98948 106614 99000
rect 102778 97928 102784 97980
rect 102836 97968 102842 97980
rect 105538 97968 105544 97980
rect 102836 97940 105544 97968
rect 102836 97928 102842 97940
rect 105538 97928 105544 97940
rect 105596 97928 105602 97980
rect 178034 97928 178040 97980
rect 178092 97968 178098 97980
rect 406378 97968 406384 97980
rect 178092 97940 406384 97968
rect 178092 97928 178098 97940
rect 406378 97928 406384 97940
rect 406436 97928 406442 97980
rect 77938 96636 77944 96688
rect 77996 96676 78002 96688
rect 77996 96648 78812 96676
rect 77996 96636 78002 96648
rect 78784 96608 78812 96648
rect 81894 96608 81900 96620
rect 78784 96580 81900 96608
rect 81894 96568 81900 96580
rect 81952 96568 81958 96620
rect 341518 95888 341524 95940
rect 341576 95928 341582 95940
rect 348418 95928 348424 95940
rect 341576 95900 348424 95928
rect 341576 95888 341582 95900
rect 348418 95888 348424 95900
rect 348476 95888 348482 95940
rect 106550 95140 106556 95192
rect 106608 95180 106614 95192
rect 108390 95180 108396 95192
rect 106608 95152 108396 95180
rect 106608 95140 106614 95152
rect 108390 95140 108396 95152
rect 108448 95140 108454 95192
rect 178034 95140 178040 95192
rect 178092 95180 178098 95192
rect 404998 95180 405004 95192
rect 178092 95152 405004 95180
rect 178092 95140 178098 95152
rect 404998 95140 405004 95152
rect 405056 95140 405062 95192
rect 81894 93780 81900 93832
rect 81952 93820 81958 93832
rect 84838 93820 84844 93832
rect 81952 93792 84844 93820
rect 81952 93780 81958 93792
rect 84838 93780 84844 93792
rect 84896 93780 84902 93832
rect 178034 93780 178040 93832
rect 178092 93820 178098 93832
rect 403618 93820 403624 93832
rect 178092 93792 403624 93820
rect 178092 93780 178098 93792
rect 403618 93780 403624 93792
rect 403676 93780 403682 93832
rect 178034 92420 178040 92472
rect 178092 92460 178098 92472
rect 400858 92460 400864 92472
rect 178092 92432 400864 92460
rect 178092 92420 178098 92432
rect 400858 92420 400864 92432
rect 400916 92420 400922 92472
rect 178034 90992 178040 91044
rect 178092 91032 178098 91044
rect 399478 91032 399484 91044
rect 178092 91004 399484 91032
rect 178092 90992 178098 91004
rect 399478 90992 399484 91004
rect 399536 90992 399542 91044
rect 108390 90108 108396 90160
rect 108448 90148 108454 90160
rect 109770 90148 109776 90160
rect 108448 90120 109776 90148
rect 108448 90108 108454 90120
rect 109770 90108 109776 90120
rect 109828 90108 109834 90160
rect 178034 89632 178040 89684
rect 178092 89672 178098 89684
rect 418798 89672 418804 89684
rect 178092 89644 418804 89672
rect 178092 89632 178098 89644
rect 418798 89632 418804 89644
rect 418856 89632 418862 89684
rect 178034 88272 178040 88324
rect 178092 88312 178098 88324
rect 417418 88312 417424 88324
rect 178092 88284 417424 88312
rect 178092 88272 178098 88284
rect 417418 88272 417424 88284
rect 417476 88272 417482 88324
rect 109770 86912 109776 86964
rect 109828 86952 109834 86964
rect 110966 86952 110972 86964
rect 109828 86924 110972 86952
rect 109828 86912 109834 86924
rect 110966 86912 110972 86924
rect 111024 86912 111030 86964
rect 178034 86912 178040 86964
rect 178092 86952 178098 86964
rect 414658 86952 414664 86964
rect 178092 86924 414664 86952
rect 178092 86912 178098 86924
rect 414658 86912 414664 86924
rect 414716 86912 414722 86964
rect 178678 85552 178684 85604
rect 178736 85592 178742 85604
rect 580166 85592 580172 85604
rect 178736 85564 580172 85592
rect 178736 85552 178742 85564
rect 580166 85552 580172 85564
rect 580224 85552 580230 85604
rect 178034 85484 178040 85536
rect 178092 85524 178098 85536
rect 188338 85524 188344 85536
rect 178092 85496 188344 85524
rect 178092 85484 178098 85496
rect 188338 85484 188344 85496
rect 188396 85484 188402 85536
rect 105538 84804 105544 84856
rect 105596 84844 105602 84856
rect 116762 84844 116768 84856
rect 105596 84816 116768 84844
rect 105596 84804 105602 84816
rect 116762 84804 116768 84816
rect 116820 84804 116826 84856
rect 3326 84192 3332 84244
rect 3384 84232 3390 84244
rect 116670 84232 116676 84244
rect 3384 84204 116676 84232
rect 3384 84192 3390 84204
rect 116670 84192 116676 84204
rect 116728 84192 116734 84244
rect 178034 84124 178040 84176
rect 178092 84164 178098 84176
rect 185578 84164 185584 84176
rect 178092 84136 185584 84164
rect 178092 84124 178098 84136
rect 185578 84124 185584 84136
rect 185636 84124 185642 84176
rect 178034 82764 178040 82816
rect 178092 82804 178098 82816
rect 184198 82804 184204 82816
rect 178092 82776 184204 82804
rect 178092 82764 178098 82776
rect 184198 82764 184204 82776
rect 184256 82764 184262 82816
rect 332594 82084 332600 82136
rect 332652 82124 332658 82136
rect 341518 82124 341524 82136
rect 332652 82096 341524 82124
rect 332652 82084 332658 82096
rect 341518 82084 341524 82096
rect 341576 82084 341582 82136
rect 110966 79976 110972 80028
rect 111024 80016 111030 80028
rect 115842 80016 115848 80028
rect 111024 79988 115848 80016
rect 111024 79976 111030 79988
rect 115842 79976 115848 79988
rect 115900 79976 115906 80028
rect 324314 79296 324320 79348
rect 324372 79336 324378 79348
rect 332594 79336 332600 79348
rect 324372 79308 332600 79336
rect 324372 79296 324378 79308
rect 332594 79296 332600 79308
rect 332652 79296 332658 79348
rect 178034 75896 178040 75948
rect 178092 75936 178098 75948
rect 562318 75936 562324 75948
rect 178092 75908 562324 75936
rect 178092 75896 178098 75908
rect 562318 75896 562324 75908
rect 562376 75896 562382 75948
rect 153166 75704 166580 75732
rect 115934 75624 115940 75676
rect 115992 75664 115998 75676
rect 120350 75664 120356 75676
rect 115992 75636 120356 75664
rect 115992 75624 115998 75636
rect 120350 75624 120356 75636
rect 120408 75624 120414 75676
rect 5258 75216 5264 75268
rect 5316 75256 5322 75268
rect 153166 75256 153194 75704
rect 155926 75636 160094 75664
rect 155926 75596 155954 75636
rect 5316 75228 153194 75256
rect 153396 75568 155954 75596
rect 5316 75216 5322 75228
rect 153396 75188 153424 75568
rect 160066 75528 160094 75636
rect 165724 75568 166120 75596
rect 165724 75528 165752 75568
rect 147646 75160 153424 75188
rect 155926 75500 157334 75528
rect 160066 75500 165108 75528
rect 147646 74984 147674 75160
rect 141804 74956 144914 74984
rect 141804 74928 141832 74956
rect 141786 74876 141792 74928
rect 141844 74876 141850 74928
rect 144886 74916 144914 74956
rect 145208 74956 147674 74984
rect 145208 74916 145236 74956
rect 144886 74888 145236 74916
rect 140958 74808 140964 74860
rect 141016 74848 141022 74860
rect 141016 74820 147674 74848
rect 141016 74808 141022 74820
rect 147646 74780 147674 74820
rect 155926 74780 155954 75500
rect 157306 75460 157334 75500
rect 165080 75460 165108 75500
rect 165356 75500 165752 75528
rect 166092 75528 166120 75568
rect 166552 75528 166580 75704
rect 166966 75704 170444 75732
rect 166966 75528 166994 75704
rect 170416 75676 170444 75704
rect 170398 75624 170404 75676
rect 170456 75624 170462 75676
rect 166092 75500 166488 75528
rect 166552 75500 166994 75528
rect 157306 75432 165016 75460
rect 165080 75432 165200 75460
rect 157996 75364 164832 75392
rect 157996 75188 158024 75364
rect 147646 74752 155954 74780
rect 156064 75160 158024 75188
rect 156064 74780 156092 75160
rect 164804 75120 164832 75364
rect 164988 75188 165016 75432
rect 165172 75392 165200 75432
rect 165356 75392 165384 75500
rect 166460 75460 166488 75500
rect 171318 75460 171324 75472
rect 166460 75432 171324 75460
rect 171318 75420 171324 75432
rect 171376 75420 171382 75472
rect 171410 75420 171416 75472
rect 171468 75460 171474 75472
rect 176562 75460 176568 75472
rect 171468 75432 176568 75460
rect 171468 75420 171474 75432
rect 176562 75420 176568 75432
rect 176620 75420 176626 75472
rect 171134 75392 171140 75404
rect 165172 75364 165384 75392
rect 166644 75364 171140 75392
rect 166644 75188 166672 75364
rect 171134 75352 171140 75364
rect 171192 75352 171198 75404
rect 195974 75324 195980 75336
rect 164988 75160 166672 75188
rect 167564 75296 195980 75324
rect 167564 75120 167592 75296
rect 195974 75284 195980 75296
rect 196032 75284 196038 75336
rect 170490 75256 170496 75268
rect 156524 75092 161474 75120
rect 164804 75092 167592 75120
rect 167932 75228 170496 75256
rect 156138 74876 156144 74928
rect 156196 74916 156202 74928
rect 156524 74916 156552 75092
rect 161446 75052 161474 75092
rect 167932 75052 167960 75228
rect 170490 75216 170496 75228
rect 170548 75216 170554 75268
rect 171134 75148 171140 75200
rect 171192 75188 171198 75200
rect 249794 75188 249800 75200
rect 171192 75160 249800 75188
rect 171192 75148 171198 75160
rect 249794 75148 249800 75160
rect 249852 75148 249858 75200
rect 171318 75080 171324 75132
rect 171376 75120 171382 75132
rect 259454 75120 259460 75132
rect 171376 75092 259460 75120
rect 171376 75080 171382 75092
rect 259454 75080 259460 75092
rect 259512 75080 259518 75132
rect 156196 74888 156552 74916
rect 156616 75024 160048 75052
rect 161446 75024 167960 75052
rect 156196 74876 156202 74888
rect 156138 74780 156144 74792
rect 156064 74752 156144 74780
rect 156138 74740 156144 74752
rect 156196 74740 156202 74792
rect 156616 74712 156644 75024
rect 160020 74984 160048 75024
rect 176378 75012 176384 75064
rect 176436 75052 176442 75064
rect 324314 75052 324320 75064
rect 176436 75024 324320 75052
rect 176436 75012 176442 75024
rect 324314 75012 324320 75024
rect 324372 75012 324378 75064
rect 320174 74984 320180 74996
rect 157536 74956 159956 74984
rect 160020 74956 320180 74984
rect 157536 74848 157564 74956
rect 159928 74916 159956 74956
rect 320174 74944 320180 74956
rect 320232 74944 320238 74996
rect 338114 74916 338120 74928
rect 159928 74888 338120 74916
rect 338114 74876 338120 74888
rect 338172 74876 338178 74928
rect 156800 74820 157564 74848
rect 157720 74820 165614 74848
rect 156800 74780 156828 74820
rect 147784 74684 156644 74712
rect 156708 74752 156828 74780
rect 146478 74536 146484 74588
rect 146536 74576 146542 74588
rect 147784 74576 147812 74684
rect 147858 74604 147864 74656
rect 147916 74644 147922 74656
rect 156708 74644 156736 74752
rect 157518 74740 157524 74792
rect 157576 74780 157582 74792
rect 157720 74780 157748 74820
rect 165586 74780 165614 74820
rect 167546 74808 167552 74860
rect 167604 74848 167610 74860
rect 167604 74820 168512 74848
rect 167604 74808 167610 74820
rect 167730 74780 167736 74792
rect 157576 74752 157748 74780
rect 157904 74752 161474 74780
rect 165586 74752 167736 74780
rect 157576 74740 157582 74752
rect 147916 74616 156736 74644
rect 147916 74604 147922 74616
rect 157518 74604 157524 74656
rect 157576 74644 157582 74656
rect 157904 74644 157932 74752
rect 161446 74712 161474 74752
rect 167730 74740 167736 74752
rect 167788 74740 167794 74792
rect 168484 74780 168512 74820
rect 168558 74808 168564 74860
rect 168616 74848 168622 74860
rect 176378 74848 176384 74860
rect 168616 74820 176384 74848
rect 168616 74808 168622 74820
rect 176378 74808 176384 74820
rect 176436 74808 176442 74860
rect 396810 74848 396816 74860
rect 176488 74820 396816 74848
rect 176488 74780 176516 74820
rect 396810 74808 396816 74820
rect 396868 74808 396874 74860
rect 168484 74752 176516 74780
rect 176562 74740 176568 74792
rect 176620 74780 176626 74792
rect 396994 74780 397000 74792
rect 176620 74752 397000 74780
rect 176620 74740 176626 74752
rect 396994 74740 397000 74752
rect 397052 74740 397058 74792
rect 390554 74712 390560 74724
rect 161446 74684 390560 74712
rect 390554 74672 390560 74684
rect 390612 74672 390618 74724
rect 465166 74644 465172 74656
rect 157576 74616 157932 74644
rect 161446 74616 465172 74644
rect 157576 74604 157582 74616
rect 146536 74548 147812 74576
rect 146536 74536 146542 74548
rect 157794 74536 157800 74588
rect 157852 74576 157858 74588
rect 161446 74576 161474 74616
rect 465166 74604 465172 74616
rect 465224 74604 465230 74656
rect 167546 74576 167552 74588
rect 157852 74548 161474 74576
rect 164206 74548 167552 74576
rect 157852 74536 157858 74548
rect 154758 74468 154764 74520
rect 154816 74508 154822 74520
rect 164206 74508 164234 74548
rect 167546 74536 167552 74548
rect 167604 74536 167610 74588
rect 168190 74536 168196 74588
rect 168248 74576 168254 74588
rect 579614 74576 579620 74588
rect 168248 74548 579620 74576
rect 168248 74536 168254 74548
rect 579614 74536 579620 74548
rect 579672 74536 579678 74588
rect 154816 74480 164234 74508
rect 154816 74468 154822 74480
rect 167086 74468 167092 74520
rect 167144 74508 167150 74520
rect 580534 74508 580540 74520
rect 167144 74480 580540 74508
rect 167144 74468 167150 74480
rect 580534 74468 580540 74480
rect 580592 74468 580598 74520
rect 43438 74400 43444 74452
rect 43496 74440 43502 74452
rect 169754 74440 169760 74452
rect 43496 74412 169760 74440
rect 43496 74400 43502 74412
rect 169754 74400 169760 74412
rect 169812 74400 169818 74452
rect 43530 74332 43536 74384
rect 43588 74372 43594 74384
rect 169846 74372 169852 74384
rect 43588 74344 169852 74372
rect 43588 74332 43594 74344
rect 169846 74332 169852 74344
rect 169904 74332 169910 74384
rect 143718 74264 143724 74316
rect 143776 74304 143782 74316
rect 284294 74304 284300 74316
rect 143776 74276 284300 74304
rect 143776 74264 143782 74276
rect 284294 74264 284300 74276
rect 284352 74264 284358 74316
rect 145098 74196 145104 74248
rect 145156 74236 145162 74248
rect 302234 74236 302240 74248
rect 145156 74208 302240 74236
rect 145156 74196 145162 74208
rect 302234 74196 302240 74208
rect 302292 74196 302298 74248
rect 146754 74128 146760 74180
rect 146812 74168 146818 74180
rect 324314 74168 324320 74180
rect 146812 74140 324320 74168
rect 146812 74128 146818 74140
rect 324314 74128 324320 74140
rect 324372 74128 324378 74180
rect 150618 74060 150624 74112
rect 150676 74100 150682 74112
rect 373994 74100 374000 74112
rect 150676 74072 374000 74100
rect 150676 74060 150682 74072
rect 373994 74060 374000 74072
rect 374052 74060 374058 74112
rect 153378 73992 153384 74044
rect 153436 74032 153442 74044
rect 408494 74032 408500 74044
rect 153436 74004 408500 74032
rect 153436 73992 153442 74004
rect 408494 73992 408500 74004
rect 408552 73992 408558 74044
rect 112438 73924 112444 73976
rect 112496 73964 112502 73976
rect 112496 73936 164372 73964
rect 112496 73924 112502 73936
rect 115198 73856 115204 73908
rect 115256 73896 115262 73908
rect 161658 73896 161664 73908
rect 115256 73868 161664 73896
rect 115256 73856 115262 73868
rect 161658 73856 161664 73868
rect 161716 73856 161722 73908
rect 116670 73720 116676 73772
rect 116728 73760 116734 73772
rect 164344 73760 164372 73936
rect 168374 73924 168380 73976
rect 168432 73964 168438 73976
rect 462314 73964 462320 73976
rect 168432 73936 462320 73964
rect 168432 73924 168438 73936
rect 462314 73924 462320 73936
rect 462372 73924 462378 73976
rect 168282 73856 168288 73908
rect 168340 73896 168346 73908
rect 527174 73896 527180 73908
rect 168340 73868 527180 73896
rect 168340 73856 168346 73868
rect 527174 73856 527180 73868
rect 527232 73856 527238 73908
rect 164418 73788 164424 73840
rect 164476 73828 164482 73840
rect 550634 73828 550640 73840
rect 164476 73800 550640 73828
rect 164476 73788 164482 73800
rect 550634 73788 550640 73800
rect 550692 73788 550698 73840
rect 169938 73760 169944 73772
rect 116728 73732 162348 73760
rect 164344 73732 169944 73760
rect 116728 73720 116734 73732
rect 155494 73652 155500 73704
rect 155552 73692 155558 73704
rect 155552 73664 158392 73692
rect 155552 73652 155558 73664
rect 5166 73584 5172 73636
rect 5224 73624 5230 73636
rect 158364 73624 158392 73664
rect 162320 73624 162348 73732
rect 169938 73720 169944 73732
rect 169996 73720 170002 73772
rect 168190 73652 168196 73704
rect 168248 73692 168254 73704
rect 170490 73692 170496 73704
rect 168248 73664 170496 73692
rect 168248 73652 168254 73664
rect 170490 73652 170496 73664
rect 170548 73652 170554 73704
rect 170122 73624 170128 73636
rect 5224 73596 157334 73624
rect 158364 73596 161474 73624
rect 162320 73596 170128 73624
rect 5224 73584 5230 73596
rect 84838 73516 84844 73568
rect 84896 73556 84902 73568
rect 85574 73556 85580 73568
rect 84896 73528 85580 73556
rect 84896 73516 84902 73528
rect 85574 73516 85580 73528
rect 85632 73516 85638 73568
rect 131666 73380 131672 73432
rect 131724 73380 131730 73432
rect 157306 73420 157334 73596
rect 161446 73488 161474 73596
rect 170122 73584 170128 73596
rect 170180 73584 170186 73636
rect 161658 73516 161664 73568
rect 161716 73556 161722 73568
rect 170030 73556 170036 73568
rect 161716 73528 170036 73556
rect 161716 73516 161722 73528
rect 170030 73516 170036 73528
rect 170088 73516 170094 73568
rect 167178 73488 167184 73500
rect 161446 73460 167184 73488
rect 167178 73448 167184 73460
rect 167236 73448 167242 73500
rect 169570 73420 169576 73432
rect 157306 73392 169576 73420
rect 169570 73380 169576 73392
rect 169628 73380 169634 73432
rect 131684 73352 131712 73380
rect 131684 73324 131804 73352
rect 131390 73244 131396 73296
rect 131448 73284 131454 73296
rect 131666 73284 131672 73296
rect 131448 73256 131672 73284
rect 131448 73244 131454 73256
rect 131666 73244 131672 73256
rect 131724 73244 131730 73296
rect 120902 73108 120908 73160
rect 120960 73148 120966 73160
rect 127894 73148 127900 73160
rect 120960 73120 127900 73148
rect 120960 73108 120966 73120
rect 127894 73108 127900 73120
rect 127952 73108 127958 73160
rect 131390 73108 131396 73160
rect 131448 73148 131454 73160
rect 131776 73148 131804 73324
rect 147858 73176 147864 73228
rect 147916 73216 147922 73228
rect 153378 73216 153384 73228
rect 147916 73188 153384 73216
rect 147916 73176 147922 73188
rect 153378 73176 153384 73188
rect 153436 73176 153442 73228
rect 207014 73216 207020 73228
rect 162136 73188 207020 73216
rect 131448 73120 131804 73148
rect 131448 73108 131454 73120
rect 136818 73108 136824 73160
rect 136876 73148 136882 73160
rect 156138 73148 156144 73160
rect 136876 73120 156144 73148
rect 136876 73108 136882 73120
rect 156138 73108 156144 73120
rect 156196 73108 156202 73160
rect 137646 73040 137652 73092
rect 137704 73080 137710 73092
rect 162136 73080 162164 73188
rect 207014 73176 207020 73188
rect 207072 73176 207078 73228
rect 167914 73108 167920 73160
rect 167972 73148 167978 73160
rect 168282 73148 168288 73160
rect 167972 73120 168288 73148
rect 167972 73108 167978 73120
rect 168282 73108 168288 73120
rect 168340 73108 168346 73160
rect 137704 73052 162164 73080
rect 137704 73040 137710 73052
rect 167822 73040 167828 73092
rect 167880 73080 167886 73092
rect 580718 73080 580724 73092
rect 167880 73052 580724 73080
rect 167880 73040 167886 73052
rect 580718 73040 580724 73052
rect 580776 73040 580782 73092
rect 120718 72972 120724 73024
rect 120776 73012 120782 73024
rect 128170 73012 128176 73024
rect 120776 72984 128176 73012
rect 120776 72972 120782 72984
rect 128170 72972 128176 72984
rect 128228 72972 128234 73024
rect 137738 72972 137744 73024
rect 137796 73012 137802 73024
rect 145098 73012 145104 73024
rect 137796 72984 145104 73012
rect 137796 72972 137802 72984
rect 145098 72972 145104 72984
rect 145156 72972 145162 73024
rect 151814 72972 151820 73024
rect 151872 73012 151878 73024
rect 151998 73012 152004 73024
rect 151872 72984 152004 73012
rect 151872 72972 151878 72984
rect 151998 72972 152004 72984
rect 152056 72972 152062 73024
rect 152734 72972 152740 73024
rect 152792 73012 152798 73024
rect 168006 73012 168012 73024
rect 152792 72984 168012 73012
rect 152792 72972 152798 72984
rect 168006 72972 168012 72984
rect 168064 72972 168070 73024
rect 168466 72972 168472 73024
rect 168524 73012 168530 73024
rect 397454 73012 397460 73024
rect 168524 72984 397460 73012
rect 168524 72972 168530 72984
rect 397454 72972 397460 72984
rect 397512 72972 397518 73024
rect 120810 72904 120816 72956
rect 120868 72944 120874 72956
rect 129274 72944 129280 72956
rect 120868 72916 129280 72944
rect 120868 72904 120874 72916
rect 129274 72904 129280 72916
rect 129332 72904 129338 72956
rect 136266 72904 136272 72956
rect 136324 72944 136330 72956
rect 147858 72944 147864 72956
rect 136324 72916 147864 72944
rect 136324 72904 136330 72916
rect 147858 72904 147864 72916
rect 147916 72904 147922 72956
rect 150250 72904 150256 72956
rect 150308 72944 150314 72956
rect 150308 72916 151492 72944
rect 150308 72904 150314 72916
rect 119338 72836 119344 72888
rect 119396 72876 119402 72888
rect 122742 72876 122748 72888
rect 119396 72848 122748 72876
rect 119396 72836 119402 72848
rect 122742 72836 122748 72848
rect 122800 72836 122806 72888
rect 141602 72836 141608 72888
rect 141660 72876 141666 72888
rect 150618 72876 150624 72888
rect 141660 72848 150624 72876
rect 141660 72836 141666 72848
rect 150618 72836 150624 72848
rect 150676 72836 150682 72888
rect 151464 72876 151492 72916
rect 153378 72904 153384 72956
rect 153436 72944 153442 72956
rect 167914 72944 167920 72956
rect 153436 72916 167920 72944
rect 153436 72904 153442 72916
rect 167914 72904 167920 72916
rect 167972 72904 167978 72956
rect 168282 72904 168288 72956
rect 168340 72944 168346 72956
rect 217318 72944 217324 72956
rect 168340 72916 217324 72944
rect 168340 72904 168346 72916
rect 217318 72904 217324 72916
rect 217376 72904 217382 72956
rect 154758 72876 154764 72888
rect 151464 72848 154764 72876
rect 154758 72836 154764 72848
rect 154816 72836 154822 72888
rect 156598 72836 156604 72888
rect 156656 72876 156662 72888
rect 231118 72876 231124 72888
rect 156656 72848 231124 72876
rect 156656 72836 156662 72848
rect 231118 72836 231124 72848
rect 231176 72836 231182 72888
rect 121086 72768 121092 72820
rect 121144 72808 121150 72820
rect 130378 72808 130384 72820
rect 121144 72780 130384 72808
rect 121144 72768 121150 72780
rect 130378 72768 130384 72780
rect 130436 72768 130442 72820
rect 142706 72768 142712 72820
rect 142764 72808 142770 72820
rect 151814 72808 151820 72820
rect 142764 72780 151820 72808
rect 142764 72768 142770 72780
rect 151814 72768 151820 72780
rect 151872 72768 151878 72820
rect 154390 72768 154396 72820
rect 154448 72808 154454 72820
rect 154448 72780 156644 72808
rect 154448 72768 154454 72780
rect 120994 72700 121000 72752
rect 121052 72740 121058 72752
rect 129826 72740 129832 72752
rect 121052 72712 129832 72740
rect 121052 72700 121058 72712
rect 129826 72700 129832 72712
rect 129884 72700 129890 72752
rect 140498 72700 140504 72752
rect 140556 72740 140562 72752
rect 146754 72740 146760 72752
rect 140556 72712 146760 72740
rect 140556 72700 140562 72712
rect 146754 72700 146760 72712
rect 146812 72700 146818 72752
rect 151906 72700 151912 72752
rect 151964 72740 151970 72752
rect 155494 72740 155500 72752
rect 151964 72712 155500 72740
rect 151964 72700 151970 72712
rect 155494 72700 155500 72712
rect 155552 72700 155558 72752
rect 86218 72632 86224 72684
rect 86276 72672 86282 72684
rect 122374 72672 122380 72684
rect 86276 72644 122380 72672
rect 86276 72632 86282 72644
rect 122374 72632 122380 72644
rect 122432 72632 122438 72684
rect 122742 72632 122748 72684
rect 122800 72672 122806 72684
rect 127342 72672 127348 72684
rect 122800 72644 127348 72672
rect 122800 72632 122806 72644
rect 127342 72632 127348 72644
rect 127400 72632 127406 72684
rect 132310 72632 132316 72684
rect 132368 72672 132374 72684
rect 137738 72672 137744 72684
rect 132368 72644 137744 72672
rect 132368 72632 132374 72644
rect 137738 72632 137744 72644
rect 137796 72632 137802 72684
rect 138842 72632 138848 72684
rect 138900 72672 138906 72684
rect 142706 72672 142712 72684
rect 138900 72644 142712 72672
rect 138900 72632 138906 72644
rect 142706 72632 142712 72644
rect 142764 72632 142770 72684
rect 152918 72672 152924 72684
rect 143552 72644 152924 72672
rect 85574 72564 85580 72616
rect 85632 72604 85638 72616
rect 93946 72604 93952 72616
rect 85632 72576 93952 72604
rect 85632 72564 85638 72576
rect 93946 72564 93952 72576
rect 94004 72564 94010 72616
rect 132678 72604 132684 72616
rect 132466 72576 132684 72604
rect 60734 72496 60740 72548
rect 60792 72536 60798 72548
rect 126330 72536 126336 72548
rect 60792 72508 126336 72536
rect 60792 72496 60798 72508
rect 126330 72496 126336 72508
rect 126388 72496 126394 72548
rect 25498 72428 25504 72480
rect 25556 72468 25562 72480
rect 123110 72468 123116 72480
rect 25556 72440 123116 72468
rect 25556 72428 25562 72440
rect 123110 72428 123116 72440
rect 123168 72428 123174 72480
rect 121362 72360 121368 72412
rect 121420 72400 121426 72412
rect 132466 72400 132494 72576
rect 132678 72564 132684 72576
rect 132736 72564 132742 72616
rect 139210 72564 139216 72616
rect 139268 72604 139274 72616
rect 143552 72604 143580 72644
rect 152918 72632 152924 72644
rect 152976 72632 152982 72684
rect 156616 72672 156644 72780
rect 157426 72768 157432 72820
rect 157484 72808 157490 72820
rect 239214 72808 239220 72820
rect 157484 72780 239220 72808
rect 157484 72768 157490 72780
rect 239214 72768 239220 72780
rect 239272 72768 239278 72820
rect 158254 72700 158260 72752
rect 158312 72740 158318 72752
rect 158622 72740 158628 72752
rect 158312 72712 158628 72740
rect 158312 72700 158318 72712
rect 158622 72700 158628 72712
rect 158680 72700 158686 72752
rect 166626 72700 166632 72752
rect 166684 72740 166690 72752
rect 259362 72740 259368 72752
rect 166684 72712 259368 72740
rect 166684 72700 166690 72712
rect 259362 72700 259368 72712
rect 259420 72700 259426 72752
rect 422294 72672 422300 72684
rect 156616 72644 422300 72672
rect 422294 72632 422300 72644
rect 422352 72632 422358 72684
rect 139268 72576 143580 72604
rect 139268 72564 139274 72576
rect 151262 72564 151268 72616
rect 151320 72604 151326 72616
rect 154114 72604 154120 72616
rect 151320 72576 154120 72604
rect 151320 72564 151326 72576
rect 154114 72564 154120 72576
rect 154172 72564 154178 72616
rect 158622 72564 158628 72616
rect 158680 72604 158686 72616
rect 471974 72604 471980 72616
rect 158680 72576 471980 72604
rect 158680 72564 158686 72576
rect 471974 72564 471980 72576
rect 472032 72564 472038 72616
rect 134702 72496 134708 72548
rect 134760 72536 134766 72548
rect 149974 72536 149980 72548
rect 134760 72508 149980 72536
rect 134760 72496 134766 72508
rect 149974 72496 149980 72508
rect 150032 72496 150038 72548
rect 151998 72496 152004 72548
rect 152056 72536 152062 72548
rect 156598 72536 156604 72548
rect 152056 72508 156604 72536
rect 152056 72496 152062 72508
rect 156598 72496 156604 72508
rect 156656 72496 156662 72548
rect 166718 72496 166724 72548
rect 166776 72536 166782 72548
rect 520918 72536 520924 72548
rect 166776 72508 520924 72536
rect 166776 72496 166782 72508
rect 520918 72496 520924 72508
rect 520976 72496 520982 72548
rect 135714 72428 135720 72480
rect 135772 72468 135778 72480
rect 165246 72468 165252 72480
rect 135772 72440 165252 72468
rect 135772 72428 135778 72440
rect 165246 72428 165252 72440
rect 165304 72428 165310 72480
rect 166902 72428 166908 72480
rect 166960 72468 166966 72480
rect 580258 72468 580264 72480
rect 166960 72440 580264 72468
rect 166960 72428 166966 72440
rect 580258 72428 580264 72440
rect 580316 72428 580322 72480
rect 121420 72372 132494 72400
rect 121420 72360 121426 72372
rect 142154 72360 142160 72412
rect 142212 72400 142218 72412
rect 152918 72400 152924 72412
rect 142212 72372 152924 72400
rect 142212 72360 142218 72372
rect 152918 72360 152924 72372
rect 152976 72360 152982 72412
rect 156046 72360 156052 72412
rect 156104 72400 156110 72412
rect 171778 72400 171784 72412
rect 156104 72372 171784 72400
rect 156104 72360 156110 72372
rect 171778 72360 171784 72372
rect 171836 72360 171842 72412
rect 133966 72292 133972 72344
rect 134024 72332 134030 72344
rect 137646 72332 137652 72344
rect 134024 72304 137652 72332
rect 134024 72292 134030 72304
rect 137646 72292 137652 72304
rect 137704 72292 137710 72344
rect 150802 72292 150808 72344
rect 150860 72332 150866 72344
rect 152826 72332 152832 72344
rect 150860 72304 152832 72332
rect 150860 72292 150866 72304
rect 152826 72292 152832 72304
rect 152884 72292 152890 72344
rect 167638 72332 167644 72344
rect 153764 72304 167644 72332
rect 145466 72224 145472 72276
rect 145524 72264 145530 72276
rect 145524 72236 151032 72264
rect 145524 72224 145530 72236
rect 116670 72156 116676 72208
rect 116728 72196 116734 72208
rect 124858 72196 124864 72208
rect 116728 72168 124864 72196
rect 116728 72156 116734 72168
rect 124858 72156 124864 72168
rect 124916 72156 124922 72208
rect 142706 72156 142712 72208
rect 142764 72196 142770 72208
rect 150158 72196 150164 72208
rect 142764 72168 150164 72196
rect 142764 72156 142770 72168
rect 150158 72156 150164 72168
rect 150216 72156 150222 72208
rect 118142 72088 118148 72140
rect 118200 72128 118206 72140
rect 124306 72128 124312 72140
rect 118200 72100 124312 72128
rect 118200 72088 118206 72100
rect 124306 72088 124312 72100
rect 124364 72088 124370 72140
rect 151004 72128 151032 72236
rect 151814 72224 151820 72276
rect 151872 72264 151878 72276
rect 153010 72264 153016 72276
rect 151872 72236 153016 72264
rect 151872 72224 151878 72236
rect 153010 72224 153016 72236
rect 153068 72224 153074 72276
rect 152182 72156 152188 72208
rect 152240 72196 152246 72208
rect 153764 72196 153792 72304
rect 167638 72292 167644 72304
rect 167696 72292 167702 72344
rect 154942 72224 154948 72276
rect 155000 72264 155006 72276
rect 169018 72264 169024 72276
rect 155000 72236 169024 72264
rect 155000 72224 155006 72236
rect 169018 72224 169024 72236
rect 169076 72224 169082 72276
rect 152240 72168 153792 72196
rect 152240 72156 152246 72168
rect 153838 72156 153844 72208
rect 153896 72196 153902 72208
rect 167730 72196 167736 72208
rect 153896 72168 167736 72196
rect 153896 72156 153902 72168
rect 167730 72156 167736 72168
rect 167788 72156 167794 72208
rect 154298 72128 154304 72140
rect 151004 72100 154304 72128
rect 154298 72088 154304 72100
rect 154356 72088 154362 72140
rect 167362 72128 167368 72140
rect 162136 72100 167368 72128
rect 117958 72020 117964 72072
rect 118016 72060 118022 72072
rect 123754 72060 123760 72072
rect 118016 72032 123760 72060
rect 118016 72020 118022 72032
rect 123754 72020 123760 72032
rect 123812 72020 123818 72072
rect 145098 72020 145104 72072
rect 145156 72060 145162 72072
rect 146018 72060 146024 72072
rect 145156 72032 146024 72060
rect 145156 72020 145162 72032
rect 146018 72020 146024 72032
rect 146076 72020 146082 72072
rect 151354 72020 151360 72072
rect 151412 72060 151418 72072
rect 158438 72060 158444 72072
rect 151412 72032 158444 72060
rect 151412 72020 151418 72032
rect 158438 72020 158444 72032
rect 158496 72020 158502 72072
rect 118050 71952 118056 72004
rect 118108 71992 118114 72004
rect 123018 71992 123024 72004
rect 118108 71964 123024 71992
rect 118108 71952 118114 71964
rect 123018 71952 123024 71964
rect 123076 71952 123082 72004
rect 149146 71952 149152 72004
rect 149204 71992 149210 72004
rect 154390 71992 154396 72004
rect 149204 71964 154396 71992
rect 149204 71952 149210 71964
rect 154390 71952 154396 71964
rect 154448 71952 154454 72004
rect 149698 71884 149704 71936
rect 149756 71924 149762 71936
rect 156874 71924 156880 71936
rect 149756 71896 156880 71924
rect 149756 71884 149762 71896
rect 156874 71884 156880 71896
rect 156932 71884 156938 71936
rect 127710 71816 127716 71868
rect 127768 71856 127774 71868
rect 128078 71856 128084 71868
rect 127768 71828 128084 71856
rect 127768 71816 127774 71828
rect 128078 71816 128084 71828
rect 128136 71816 128142 71868
rect 146754 71816 146760 71868
rect 146812 71856 146818 71868
rect 151630 71856 151636 71868
rect 146812 71828 151636 71856
rect 146812 71816 146818 71828
rect 151630 71816 151636 71828
rect 151688 71816 151694 71868
rect 153286 71816 153292 71868
rect 153344 71856 153350 71868
rect 162136 71856 162164 72100
rect 167362 72088 167368 72100
rect 167420 72088 167426 72140
rect 162762 72020 162768 72072
rect 162820 72060 162826 72072
rect 166718 72060 166724 72072
rect 162820 72032 166724 72060
rect 162820 72020 162826 72032
rect 166718 72020 166724 72032
rect 166776 72020 166782 72072
rect 178586 72060 178592 72072
rect 166966 72032 178592 72060
rect 153344 71828 162164 71856
rect 153344 71816 153350 71828
rect 165062 71816 165068 71868
rect 165120 71856 165126 71868
rect 166626 71856 166632 71868
rect 165120 71828 166632 71856
rect 165120 71816 165126 71828
rect 166626 71816 166632 71828
rect 166684 71816 166690 71868
rect 132494 71748 132500 71800
rect 132552 71788 132558 71800
rect 136174 71788 136180 71800
rect 132552 71760 136180 71788
rect 132552 71748 132558 71760
rect 136174 71748 136180 71760
rect 136232 71748 136238 71800
rect 136634 71748 136640 71800
rect 136692 71788 136698 71800
rect 143258 71788 143264 71800
rect 136692 71760 143264 71788
rect 136692 71748 136698 71760
rect 143258 71748 143264 71760
rect 143316 71748 143322 71800
rect 145834 71748 145840 71800
rect 145892 71788 145898 71800
rect 147306 71788 147312 71800
rect 145892 71760 147312 71788
rect 145892 71748 145898 71760
rect 147306 71748 147312 71760
rect 147364 71748 147370 71800
rect 3510 71680 3516 71732
rect 3568 71720 3574 71732
rect 166966 71720 166994 72032
rect 178586 72020 178592 72032
rect 178644 72020 178650 72072
rect 167270 71952 167276 72004
rect 167328 71992 167334 72004
rect 580166 71992 580172 72004
rect 167328 71964 580172 71992
rect 167328 71952 167334 71964
rect 580166 71952 580172 71964
rect 580224 71952 580230 72004
rect 3568 71692 166994 71720
rect 3568 71680 3574 71692
rect 93946 71612 93952 71664
rect 94004 71652 94010 71664
rect 168650 71652 168656 71664
rect 94004 71624 168656 71652
rect 94004 71612 94010 71624
rect 168650 71612 168656 71624
rect 168708 71612 168714 71664
rect 127618 71544 127624 71596
rect 127676 71584 127682 71596
rect 168742 71584 168748 71596
rect 127676 71556 168748 71584
rect 127676 71544 127682 71556
rect 168742 71544 168748 71556
rect 168800 71544 168806 71596
rect 168926 71516 168932 71528
rect 122806 71488 168932 71516
rect 116762 71068 116768 71120
rect 116820 71108 116826 71120
rect 122806 71108 122834 71488
rect 168926 71476 168932 71488
rect 168984 71476 168990 71528
rect 168834 71448 168840 71460
rect 116820 71080 122834 71108
rect 132466 71420 168840 71448
rect 116820 71068 116826 71080
rect 116578 70932 116584 70984
rect 116636 70972 116642 70984
rect 127618 70972 127624 70984
rect 116636 70944 127624 70972
rect 116636 70932 116642 70944
rect 127618 70932 127624 70944
rect 127676 70932 127682 70984
rect 120350 70864 120356 70916
rect 120408 70904 120414 70916
rect 132466 70904 132494 71420
rect 168834 71408 168840 71420
rect 168892 71408 168898 71460
rect 259362 71000 259368 71052
rect 259420 71040 259426 71052
rect 581086 71040 581092 71052
rect 259420 71012 581092 71040
rect 259420 71000 259426 71012
rect 581086 71000 581092 71012
rect 581144 71000 581150 71052
rect 120408 70876 132494 70904
rect 120408 70864 120414 70876
rect 123018 69912 123024 69964
rect 123076 69952 123082 69964
rect 123570 69952 123576 69964
rect 123076 69924 123576 69952
rect 123076 69912 123082 69924
rect 123570 69912 123576 69924
rect 123628 69912 123634 69964
rect 129090 69912 129096 69964
rect 129148 69952 129154 69964
rect 129642 69952 129648 69964
rect 129148 69924 129648 69952
rect 129148 69912 129154 69924
rect 129642 69912 129648 69924
rect 129700 69912 129706 69964
rect 138750 69912 138756 69964
rect 138808 69912 138814 69964
rect 121914 69844 121920 69896
rect 121972 69884 121978 69896
rect 122558 69884 122564 69896
rect 121972 69856 122564 69884
rect 121972 69844 121978 69856
rect 122558 69844 122564 69856
rect 122616 69844 122622 69896
rect 125778 69844 125784 69896
rect 125836 69884 125842 69896
rect 126606 69884 126612 69896
rect 125836 69856 126612 69884
rect 125836 69844 125842 69856
rect 126606 69844 126612 69856
rect 126664 69844 126670 69896
rect 130470 69884 130476 69896
rect 130028 69856 130476 69884
rect 122374 69776 122380 69828
rect 122432 69816 122438 69828
rect 122650 69816 122656 69828
rect 122432 69788 122656 69816
rect 122432 69776 122438 69788
rect 122650 69776 122656 69788
rect 122708 69776 122714 69828
rect 122926 69776 122932 69828
rect 122984 69816 122990 69828
rect 124122 69816 124128 69828
rect 122984 69788 124128 69816
rect 122984 69776 122990 69788
rect 124122 69776 124128 69788
rect 124180 69776 124186 69828
rect 124950 69816 124956 69828
rect 124600 69788 124956 69816
rect 123110 69708 123116 69760
rect 123168 69748 123174 69760
rect 123846 69748 123852 69760
rect 123168 69720 123852 69748
rect 123168 69708 123174 69720
rect 123846 69708 123852 69720
rect 123904 69708 123910 69760
rect 121730 69640 121736 69692
rect 121788 69680 121794 69692
rect 122190 69680 122196 69692
rect 121788 69652 122196 69680
rect 121788 69640 121794 69652
rect 122190 69640 122196 69652
rect 122248 69640 122254 69692
rect 123202 69640 123208 69692
rect 123260 69680 123266 69692
rect 123754 69680 123760 69692
rect 123260 69652 123760 69680
rect 123260 69640 123266 69652
rect 123754 69640 123760 69652
rect 123812 69640 123818 69692
rect 124600 69624 124628 69788
rect 124950 69776 124956 69788
rect 125008 69776 125014 69828
rect 126054 69708 126060 69760
rect 126112 69748 126118 69760
rect 126606 69748 126612 69760
rect 126112 69720 126612 69748
rect 126112 69708 126118 69720
rect 126606 69708 126612 69720
rect 126664 69708 126670 69760
rect 126330 69640 126336 69692
rect 126388 69680 126394 69692
rect 126790 69680 126796 69692
rect 126388 69652 126796 69680
rect 126388 69640 126394 69652
rect 126790 69640 126796 69652
rect 126848 69640 126854 69692
rect 127710 69640 127716 69692
rect 127768 69680 127774 69692
rect 128170 69680 128176 69692
rect 127768 69652 128176 69680
rect 127768 69640 127774 69652
rect 128170 69640 128176 69652
rect 128228 69640 128234 69692
rect 128538 69640 128544 69692
rect 128596 69680 128602 69692
rect 128814 69680 128820 69692
rect 128596 69652 128820 69680
rect 128596 69640 128602 69652
rect 128814 69640 128820 69652
rect 128872 69640 128878 69692
rect 128998 69640 129004 69692
rect 129056 69680 129062 69692
rect 129182 69680 129188 69692
rect 129056 69652 129188 69680
rect 129056 69640 129062 69652
rect 129182 69640 129188 69652
rect 129240 69640 129246 69692
rect 130028 69624 130056 69856
rect 130470 69844 130476 69856
rect 130528 69844 130534 69896
rect 130102 69776 130108 69828
rect 130160 69776 130166 69828
rect 130562 69776 130568 69828
rect 130620 69776 130626 69828
rect 138106 69776 138112 69828
rect 138164 69816 138170 69828
rect 138164 69788 138704 69816
rect 138164 69776 138170 69788
rect 122098 69572 122104 69624
rect 122156 69612 122162 69624
rect 122558 69612 122564 69624
rect 122156 69584 122564 69612
rect 122156 69572 122162 69584
rect 122558 69572 122564 69584
rect 122616 69572 122622 69624
rect 123386 69572 123392 69624
rect 123444 69612 123450 69624
rect 123938 69612 123944 69624
rect 123444 69584 123944 69612
rect 123444 69572 123450 69584
rect 123938 69572 123944 69584
rect 123996 69572 124002 69624
rect 124582 69572 124588 69624
rect 124640 69572 124646 69624
rect 125686 69572 125692 69624
rect 125744 69612 125750 69624
rect 126882 69612 126888 69624
rect 125744 69584 126888 69612
rect 125744 69572 125750 69584
rect 126882 69572 126888 69584
rect 126940 69572 126946 69624
rect 128630 69572 128636 69624
rect 128688 69612 128694 69624
rect 129734 69612 129740 69624
rect 128688 69584 129740 69612
rect 128688 69572 128694 69584
rect 129734 69572 129740 69584
rect 129792 69572 129798 69624
rect 130010 69572 130016 69624
rect 130068 69572 130074 69624
rect 124490 69504 124496 69556
rect 124548 69544 124554 69556
rect 125318 69544 125324 69556
rect 124548 69516 125324 69544
rect 124548 69504 124554 69516
rect 125318 69504 125324 69516
rect 125376 69504 125382 69556
rect 130120 69544 130148 69776
rect 130580 69680 130608 69776
rect 130212 69652 130608 69680
rect 130212 69624 130240 69652
rect 138676 69624 138704 69788
rect 138768 69692 138796 69912
rect 138750 69640 138756 69692
rect 138808 69640 138814 69692
rect 156598 69640 156604 69692
rect 156656 69680 156662 69692
rect 156966 69680 156972 69692
rect 156656 69652 156972 69680
rect 156656 69640 156662 69652
rect 156966 69640 156972 69652
rect 157024 69640 157030 69692
rect 167546 69680 167552 69692
rect 167288 69652 167552 69680
rect 167288 69624 167316 69652
rect 167546 69640 167552 69652
rect 167604 69640 167610 69692
rect 130194 69572 130200 69624
rect 130252 69572 130258 69624
rect 130562 69572 130568 69624
rect 130620 69612 130626 69624
rect 130930 69612 130936 69624
rect 130620 69584 130936 69612
rect 130620 69572 130626 69584
rect 130930 69572 130936 69584
rect 130988 69572 130994 69624
rect 138658 69572 138664 69624
rect 138716 69572 138722 69624
rect 167270 69572 167276 69624
rect 167328 69572 167334 69624
rect 130470 69544 130476 69556
rect 130120 69516 130476 69544
rect 130470 69504 130476 69516
rect 130528 69504 130534 69556
rect 124858 69436 124864 69488
rect 124916 69476 124922 69488
rect 125410 69476 125416 69488
rect 124916 69448 125416 69476
rect 124916 69436 124922 69448
rect 125410 69436 125416 69448
rect 125468 69436 125474 69488
rect 130102 69436 130108 69488
rect 130160 69476 130166 69488
rect 130838 69476 130844 69488
rect 130160 69448 130844 69476
rect 130160 69436 130166 69448
rect 130838 69436 130844 69448
rect 130896 69436 130902 69488
rect 167546 69436 167552 69488
rect 167604 69476 167610 69488
rect 167914 69476 167920 69488
rect 167604 69448 167920 69476
rect 167604 69436 167610 69448
rect 167914 69436 167920 69448
rect 167972 69436 167978 69488
rect 154758 68824 154764 68876
rect 154816 68864 154822 68876
rect 158346 68864 158352 68876
rect 154816 68836 158352 68864
rect 154816 68824 154822 68836
rect 158346 68824 158352 68836
rect 158404 68824 158410 68876
rect 131390 68280 131396 68332
rect 131448 68280 131454 68332
rect 239214 68280 239220 68332
rect 239272 68320 239278 68332
rect 460934 68320 460940 68332
rect 239272 68292 460940 68320
rect 239272 68280 239278 68292
rect 460934 68280 460940 68292
rect 460992 68280 460998 68332
rect 127434 68184 127440 68196
rect 127360 68156 127440 68184
rect 127360 67924 127388 68156
rect 127434 68144 127440 68156
rect 127492 68144 127498 68196
rect 131298 67940 131304 67992
rect 131356 67980 131362 67992
rect 131408 67980 131436 68280
rect 131356 67952 131436 67980
rect 131356 67940 131362 67952
rect 127342 67872 127348 67924
rect 127400 67872 127406 67924
rect 123294 67804 123300 67856
rect 123352 67844 123358 67856
rect 123662 67844 123668 67856
rect 123352 67816 123668 67844
rect 123352 67804 123358 67816
rect 123662 67804 123668 67816
rect 123720 67804 123726 67856
rect 125962 67804 125968 67856
rect 126020 67844 126026 67856
rect 126238 67844 126244 67856
rect 126020 67816 126244 67844
rect 126020 67804 126026 67816
rect 126238 67804 126244 67816
rect 126296 67804 126302 67856
rect 127434 67804 127440 67856
rect 127492 67844 127498 67856
rect 127894 67844 127900 67856
rect 127492 67816 127900 67844
rect 127492 67804 127498 67816
rect 127894 67804 127900 67816
rect 127952 67804 127958 67856
rect 128722 67804 128728 67856
rect 128780 67844 128786 67856
rect 129090 67844 129096 67856
rect 128780 67816 129096 67844
rect 128780 67804 128786 67816
rect 129090 67804 129096 67816
rect 129148 67804 129154 67856
rect 127250 67736 127256 67788
rect 127308 67776 127314 67788
rect 128262 67776 128268 67788
rect 127308 67748 128268 67776
rect 127308 67736 127314 67748
rect 128262 67736 128268 67748
rect 128320 67736 128326 67788
rect 128998 67736 129004 67788
rect 129056 67776 129062 67788
rect 129550 67776 129556 67788
rect 129056 67748 129556 67776
rect 129056 67736 129062 67748
rect 129550 67736 129556 67748
rect 129608 67736 129614 67788
rect 123662 67668 123668 67720
rect 123720 67708 123726 67720
rect 124030 67708 124036 67720
rect 123720 67680 124036 67708
rect 123720 67668 123726 67680
rect 124030 67668 124036 67680
rect 124088 67668 124094 67720
rect 128722 67668 128728 67720
rect 128780 67708 128786 67720
rect 129458 67708 129464 67720
rect 128780 67680 129464 67708
rect 128780 67668 128786 67680
rect 129458 67668 129464 67680
rect 129516 67668 129522 67720
rect 126054 67532 126060 67584
rect 126112 67572 126118 67584
rect 126422 67572 126428 67584
rect 126112 67544 126428 67572
rect 126112 67532 126118 67544
rect 126422 67532 126428 67544
rect 126480 67532 126486 67584
rect 125962 67464 125968 67516
rect 126020 67504 126026 67516
rect 126698 67504 126704 67516
rect 126020 67476 126704 67504
rect 126020 67464 126026 67476
rect 126698 67464 126704 67476
rect 126756 67464 126762 67516
rect 122006 67232 122012 67244
rect 103486 67204 122012 67232
rect 5534 66852 5540 66904
rect 5592 66892 5598 66904
rect 103486 66892 103514 67204
rect 122006 67192 122012 67204
rect 122064 67192 122070 67244
rect 5592 66864 103514 66892
rect 5592 66852 5598 66864
rect 121638 66852 121644 66904
rect 121696 66892 121702 66904
rect 122282 66892 122288 66904
rect 121696 66864 122288 66892
rect 121696 66852 121702 66864
rect 122282 66852 122288 66864
rect 122340 66852 122346 66904
rect 122190 66784 122196 66836
rect 122248 66824 122254 66836
rect 122742 66824 122748 66836
rect 122248 66796 122748 66824
rect 122248 66784 122254 66796
rect 122742 66784 122748 66796
rect 122800 66784 122806 66836
rect 124766 66172 124772 66224
rect 124824 66212 124830 66224
rect 125042 66212 125048 66224
rect 124824 66184 125048 66212
rect 124824 66172 124830 66184
rect 125042 66172 125048 66184
rect 125100 66172 125106 66224
rect 114370 60664 114376 60716
rect 114428 60704 114434 60716
rect 580166 60704 580172 60716
rect 114428 60676 580172 60704
rect 114428 60664 114434 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 163498 58624 163504 58676
rect 163556 58664 163562 58676
rect 326338 58664 326344 58676
rect 163556 58636 326344 58664
rect 163556 58624 163562 58636
rect 326338 58624 326344 58636
rect 326396 58624 326402 58676
rect 15194 54476 15200 54528
rect 15252 54516 15258 54528
rect 119338 54516 119344 54528
rect 15252 54488 119344 54516
rect 15252 54476 15258 54488
rect 119338 54476 119344 54488
rect 119396 54476 119402 54528
rect 113174 51076 113180 51128
rect 113232 51116 113238 51128
rect 121086 51116 121092 51128
rect 113232 51088 121092 51116
rect 113232 51076 113238 51088
rect 121086 51076 121092 51088
rect 121144 51076 121150 51128
rect 178678 46860 178684 46912
rect 178736 46900 178742 46912
rect 580166 46900 580172 46912
rect 178736 46872 580172 46900
rect 178736 46860 178742 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 3510 45500 3516 45552
rect 3568 45540 3574 45552
rect 170214 45540 170220 45552
rect 3568 45512 170220 45540
rect 3568 45500 3574 45512
rect 170214 45500 170220 45512
rect 170272 45500 170278 45552
rect 106274 43392 106280 43444
rect 106332 43432 106338 43444
rect 120994 43432 121000 43444
rect 106332 43404 121000 43432
rect 106332 43392 106338 43404
rect 120994 43392 121000 43404
rect 121052 43392 121058 43444
rect 153102 40672 153108 40724
rect 153160 40712 153166 40724
rect 226334 40712 226340 40724
rect 153160 40684 226340 40712
rect 153160 40672 153166 40684
rect 226334 40672 226340 40684
rect 226392 40672 226398 40724
rect 155494 36660 155500 36712
rect 155552 36700 155558 36712
rect 390646 36700 390652 36712
rect 155552 36672 390652 36700
rect 155552 36660 155558 36672
rect 390646 36660 390652 36672
rect 390704 36660 390710 36712
rect 152458 36592 152464 36644
rect 152516 36632 152522 36644
rect 397454 36632 397460 36644
rect 152516 36604 397460 36632
rect 152516 36592 152522 36604
rect 397454 36592 397460 36604
rect 397512 36592 397518 36644
rect 157794 36524 157800 36576
rect 157852 36564 157858 36576
rect 456794 36564 456800 36576
rect 157852 36536 456800 36564
rect 157852 36524 157858 36536
rect 456794 36524 456800 36536
rect 456852 36524 456858 36576
rect 145558 35844 145564 35896
rect 145616 35884 145622 35896
rect 307754 35884 307760 35896
rect 145616 35856 307760 35884
rect 145616 35844 145622 35856
rect 307754 35844 307760 35856
rect 307812 35844 307818 35896
rect 147306 35776 147312 35828
rect 147364 35816 147370 35828
rect 311894 35816 311900 35828
rect 147364 35788 311900 35816
rect 147364 35776 147370 35788
rect 311894 35776 311900 35788
rect 311952 35776 311958 35828
rect 146386 35708 146392 35760
rect 146444 35748 146450 35760
rect 318794 35748 318800 35760
rect 146444 35720 318800 35748
rect 146444 35708 146450 35720
rect 318794 35708 318800 35720
rect 318852 35708 318858 35760
rect 146662 35640 146668 35692
rect 146720 35680 146726 35692
rect 322934 35680 322940 35692
rect 146720 35652 322940 35680
rect 146720 35640 146726 35652
rect 322934 35640 322940 35652
rect 322992 35640 322998 35692
rect 146938 35572 146944 35624
rect 146996 35612 147002 35624
rect 325694 35612 325700 35624
rect 146996 35584 325700 35612
rect 146996 35572 147002 35584
rect 325694 35572 325700 35584
rect 325752 35572 325758 35624
rect 147766 35504 147772 35556
rect 147824 35544 147830 35556
rect 336734 35544 336740 35556
rect 147824 35516 336740 35544
rect 147824 35504 147830 35516
rect 336734 35504 336740 35516
rect 336792 35504 336798 35556
rect 148594 35436 148600 35488
rect 148652 35476 148658 35488
rect 347774 35476 347780 35488
rect 148652 35448 347780 35476
rect 148652 35436 148658 35448
rect 347774 35436 347780 35448
rect 347832 35436 347838 35488
rect 154482 35368 154488 35420
rect 154540 35408 154546 35420
rect 354674 35408 354680 35420
rect 154540 35380 354680 35408
rect 154540 35368 154546 35380
rect 354674 35368 354680 35380
rect 354732 35368 354738 35420
rect 149422 35300 149428 35352
rect 149480 35340 149486 35352
rect 357434 35340 357440 35352
rect 149480 35312 357440 35340
rect 149480 35300 149486 35312
rect 357434 35300 357440 35312
rect 357492 35300 357498 35352
rect 158346 35232 158352 35284
rect 158404 35272 158410 35284
rect 368474 35272 368480 35284
rect 158404 35244 368480 35272
rect 158404 35232 158410 35244
rect 368474 35232 368480 35244
rect 368532 35232 368538 35284
rect 158438 35164 158444 35216
rect 158496 35204 158502 35216
rect 382274 35204 382280 35216
rect 158496 35176 382280 35204
rect 158496 35164 158502 35176
rect 382274 35164 382280 35176
rect 382332 35164 382338 35216
rect 145282 35096 145288 35148
rect 145340 35136 145346 35148
rect 304994 35136 305000 35148
rect 145340 35108 305000 35136
rect 145340 35096 145346 35108
rect 304994 35096 305000 35108
rect 305052 35096 305058 35148
rect 138658 34416 138664 34468
rect 138716 34456 138722 34468
rect 212534 34456 212540 34468
rect 138716 34428 212540 34456
rect 138716 34416 138722 34428
rect 212534 34416 212540 34428
rect 212592 34416 212598 34468
rect 138382 34348 138388 34400
rect 138440 34388 138446 34400
rect 216674 34388 216680 34400
rect 138440 34360 216680 34388
rect 138440 34348 138446 34360
rect 216674 34348 216680 34360
rect 216732 34348 216738 34400
rect 138842 34280 138848 34332
rect 138900 34320 138906 34332
rect 219434 34320 219440 34332
rect 138900 34292 219440 34320
rect 138900 34280 138906 34292
rect 219434 34280 219440 34292
rect 219492 34280 219498 34332
rect 139762 34212 139768 34264
rect 139820 34252 139826 34264
rect 234614 34252 234620 34264
rect 139820 34224 234620 34252
rect 139820 34212 139826 34224
rect 234614 34212 234620 34224
rect 234672 34212 234678 34264
rect 140866 34144 140872 34196
rect 140924 34184 140930 34196
rect 248414 34184 248420 34196
rect 140924 34156 248420 34184
rect 140924 34144 140930 34156
rect 248414 34144 248420 34156
rect 248472 34144 248478 34196
rect 141418 34076 141424 34128
rect 141476 34116 141482 34128
rect 255314 34116 255320 34128
rect 141476 34088 255320 34116
rect 141476 34076 141482 34088
rect 255314 34076 255320 34088
rect 255372 34076 255378 34128
rect 142522 34008 142528 34060
rect 142580 34048 142586 34060
rect 269114 34048 269120 34060
rect 142580 34020 269120 34048
rect 142580 34008 142586 34020
rect 269114 34008 269120 34020
rect 269172 34008 269178 34060
rect 143074 33940 143080 33992
rect 143132 33980 143138 33992
rect 276014 33980 276020 33992
rect 143132 33952 276020 33980
rect 143132 33940 143138 33952
rect 276014 33940 276020 33952
rect 276072 33940 276078 33992
rect 143626 33872 143632 33924
rect 143684 33912 143690 33924
rect 284386 33912 284392 33924
rect 143684 33884 284392 33912
rect 143684 33872 143690 33884
rect 284386 33872 284392 33884
rect 284444 33872 284450 33924
rect 144178 33804 144184 33856
rect 144236 33844 144242 33856
rect 291194 33844 291200 33856
rect 144236 33816 291200 33844
rect 144236 33804 144242 33816
rect 291194 33804 291200 33816
rect 291252 33804 291258 33856
rect 145006 33736 145012 33788
rect 145064 33776 145070 33788
rect 300854 33776 300860 33788
rect 145064 33748 300860 33776
rect 145064 33736 145070 33748
rect 300854 33736 300860 33748
rect 300912 33736 300918 33788
rect 2866 33056 2872 33108
rect 2924 33096 2930 33108
rect 175550 33096 175556 33108
rect 2924 33068 175556 33096
rect 2924 33056 2930 33068
rect 175550 33056 175556 33068
rect 175608 33056 175614 33108
rect 135346 32920 135352 32972
rect 135404 32960 135410 32972
rect 176654 32960 176660 32972
rect 135404 32932 176660 32960
rect 135404 32920 135410 32932
rect 176654 32920 176660 32932
rect 176712 32920 176718 32972
rect 135622 32852 135628 32904
rect 135680 32892 135686 32904
rect 180794 32892 180800 32904
rect 135680 32864 180800 32892
rect 135680 32852 135686 32864
rect 180794 32852 180800 32864
rect 180852 32852 180858 32904
rect 135898 32784 135904 32836
rect 135956 32824 135962 32836
rect 184934 32824 184940 32836
rect 135956 32796 184940 32824
rect 135956 32784 135962 32796
rect 184934 32784 184940 32796
rect 184992 32784 184998 32836
rect 136726 32716 136732 32768
rect 136784 32756 136790 32768
rect 194594 32756 194600 32768
rect 136784 32728 194600 32756
rect 136784 32716 136790 32728
rect 194594 32716 194600 32728
rect 194652 32716 194658 32768
rect 137002 32648 137008 32700
rect 137060 32688 137066 32700
rect 198734 32688 198740 32700
rect 137060 32660 198740 32688
rect 137060 32648 137066 32660
rect 198734 32648 198740 32660
rect 198792 32648 198798 32700
rect 137554 32580 137560 32632
rect 137612 32620 137618 32632
rect 205634 32620 205640 32632
rect 137612 32592 205640 32620
rect 137612 32580 137618 32592
rect 205634 32580 205640 32592
rect 205692 32580 205698 32632
rect 142246 32512 142252 32564
rect 142304 32552 142310 32564
rect 266354 32552 266360 32564
rect 142304 32524 266360 32552
rect 142304 32512 142310 32524
rect 266354 32512 266360 32524
rect 266412 32512 266418 32564
rect 164326 32444 164332 32496
rect 164384 32484 164390 32496
rect 549254 32484 549260 32496
rect 164384 32456 549260 32484
rect 164384 32444 164390 32456
rect 549254 32444 549260 32456
rect 549312 32444 549318 32496
rect 166258 32376 166264 32428
rect 166316 32416 166322 32428
rect 574094 32416 574100 32428
rect 166316 32388 574100 32416
rect 166316 32376 166322 32388
rect 574094 32376 574100 32388
rect 574152 32376 574158 32428
rect 157610 31696 157616 31748
rect 157668 31736 157674 31748
rect 463694 31736 463700 31748
rect 157668 31708 463700 31736
rect 157668 31696 157674 31708
rect 463694 31696 463700 31708
rect 463752 31696 463758 31748
rect 158162 31628 158168 31680
rect 158220 31668 158226 31680
rect 470594 31668 470600 31680
rect 158220 31640 470600 31668
rect 158220 31628 158226 31640
rect 470594 31628 470600 31640
rect 470652 31628 470658 31680
rect 158714 31560 158720 31612
rect 158772 31600 158778 31612
rect 477494 31600 477500 31612
rect 158772 31572 477500 31600
rect 158772 31560 158778 31572
rect 477494 31560 477500 31572
rect 477552 31560 477558 31612
rect 159082 31492 159088 31544
rect 159140 31532 159146 31544
rect 481634 31532 481640 31544
rect 159140 31504 481640 31532
rect 159140 31492 159146 31504
rect 481634 31492 481640 31504
rect 481692 31492 481698 31544
rect 161014 31424 161020 31476
rect 161072 31464 161078 31476
rect 490006 31464 490012 31476
rect 161072 31436 490012 31464
rect 161072 31424 161078 31436
rect 490006 31424 490012 31436
rect 490064 31424 490070 31476
rect 160186 31356 160192 31408
rect 160244 31396 160250 31408
rect 496814 31396 496820 31408
rect 160244 31368 496820 31396
rect 160244 31356 160250 31368
rect 496814 31356 496820 31368
rect 496872 31356 496878 31408
rect 160738 31288 160744 31340
rect 160796 31328 160802 31340
rect 503714 31328 503720 31340
rect 160796 31300 503720 31328
rect 160796 31288 160802 31300
rect 503714 31288 503720 31300
rect 503772 31288 503778 31340
rect 162578 31220 162584 31272
rect 162636 31260 162642 31272
rect 510614 31260 510620 31272
rect 162636 31232 510620 31260
rect 162636 31220 162642 31232
rect 510614 31220 510620 31232
rect 510672 31220 510678 31272
rect 161842 31152 161848 31204
rect 161900 31192 161906 31204
rect 517514 31192 517520 31204
rect 161900 31164 517520 31192
rect 161900 31152 161906 31164
rect 517514 31152 517520 31164
rect 517572 31152 517578 31204
rect 166718 31084 166724 31136
rect 166776 31124 166782 31136
rect 524414 31124 524420 31136
rect 166776 31096 524420 31124
rect 166776 31084 166782 31096
rect 524414 31084 524420 31096
rect 524472 31084 524478 31136
rect 162118 31016 162124 31068
rect 162176 31056 162182 31068
rect 521654 31056 521660 31068
rect 162176 31028 521660 31056
rect 162176 31016 162182 31028
rect 521654 31016 521660 31028
rect 521712 31016 521718 31068
rect 154298 30268 154304 30320
rect 154356 30308 154362 30320
rect 307846 30308 307852 30320
rect 154356 30280 307852 30308
rect 154356 30268 154362 30280
rect 307846 30268 307852 30280
rect 307904 30268 307910 30320
rect 144914 30200 144920 30252
rect 144972 30240 144978 30252
rect 299474 30240 299480 30252
rect 144972 30212 299480 30240
rect 144972 30200 144978 30212
rect 299474 30200 299480 30212
rect 299532 30200 299538 30252
rect 145190 30132 145196 30184
rect 145248 30172 145254 30184
rect 303614 30172 303620 30184
rect 145248 30144 303620 30172
rect 145248 30132 145254 30144
rect 303614 30132 303620 30144
rect 303672 30132 303678 30184
rect 150710 30064 150716 30116
rect 150768 30104 150774 30116
rect 374086 30104 374092 30116
rect 150768 30076 374092 30104
rect 150768 30064 150774 30076
rect 374086 30064 374092 30076
rect 374144 30064 374150 30116
rect 154206 29996 154212 30048
rect 154264 30036 154270 30048
rect 382366 30036 382372 30048
rect 154264 30008 382372 30036
rect 154264 29996 154270 30008
rect 382366 29996 382372 30008
rect 382424 29996 382430 30048
rect 156966 29928 156972 29980
rect 157024 29968 157030 29980
rect 389174 29968 389180 29980
rect 157024 29940 389180 29968
rect 157024 29928 157030 29940
rect 389174 29928 389180 29940
rect 389232 29928 389238 29980
rect 155126 29860 155132 29912
rect 155184 29900 155190 29912
rect 431954 29900 431960 29912
rect 155184 29872 431960 29900
rect 155184 29860 155190 29872
rect 431954 29860 431960 29872
rect 432012 29860 432018 29912
rect 157058 29792 157064 29844
rect 157116 29832 157122 29844
rect 438854 29832 438860 29844
rect 157116 29804 438860 29832
rect 157116 29792 157122 29804
rect 438854 29792 438860 29804
rect 438912 29792 438918 29844
rect 155954 29724 155960 29776
rect 156012 29764 156018 29776
rect 441614 29764 441620 29776
rect 156012 29736 441620 29764
rect 156012 29724 156018 29736
rect 441614 29724 441620 29736
rect 441672 29724 441678 29776
rect 156230 29656 156236 29708
rect 156288 29696 156294 29708
rect 445754 29696 445760 29708
rect 156288 29668 445760 29696
rect 156288 29656 156294 29668
rect 445754 29656 445760 29668
rect 445812 29656 445818 29708
rect 156782 29588 156788 29640
rect 156840 29628 156846 29640
rect 452654 29628 452660 29640
rect 156840 29600 452660 29628
rect 156840 29588 156846 29600
rect 452654 29588 452660 29600
rect 452712 29588 452718 29640
rect 139394 28908 139400 28960
rect 139452 28948 139458 28960
rect 229094 28948 229100 28960
rect 139452 28920 229100 28948
rect 139452 28908 139458 28920
rect 229094 28908 229100 28920
rect 229152 28908 229158 28960
rect 151538 28840 151544 28892
rect 151596 28880 151602 28892
rect 242894 28880 242900 28892
rect 151596 28852 242900 28880
rect 151596 28840 151602 28852
rect 242894 28840 242900 28852
rect 242952 28840 242958 28892
rect 140222 28772 140228 28824
rect 140280 28812 140286 28824
rect 240134 28812 240140 28824
rect 140280 28784 240140 28812
rect 140280 28772 140286 28784
rect 240134 28772 240140 28784
rect 240192 28772 240198 28824
rect 140774 28704 140780 28756
rect 140832 28744 140838 28756
rect 247034 28744 247040 28756
rect 140832 28716 247040 28744
rect 140832 28704 140838 28716
rect 247034 28704 247040 28716
rect 247092 28704 247098 28756
rect 150618 28636 150624 28688
rect 150676 28676 150682 28688
rect 258074 28676 258080 28688
rect 150676 28648 258080 28676
rect 150676 28636 150682 28648
rect 258074 28636 258080 28648
rect 258132 28636 258138 28688
rect 141050 28568 141056 28620
rect 141108 28608 141114 28620
rect 251174 28608 251180 28620
rect 141108 28580 251180 28608
rect 141108 28568 141114 28580
rect 251174 28568 251180 28580
rect 251232 28568 251238 28620
rect 152918 28500 152924 28552
rect 152976 28540 152982 28552
rect 264974 28540 264980 28552
rect 152976 28512 264980 28540
rect 152976 28500 152982 28512
rect 264974 28500 264980 28512
rect 265032 28500 265038 28552
rect 153010 28432 153016 28484
rect 153068 28472 153074 28484
rect 271874 28472 271880 28484
rect 153068 28444 271880 28472
rect 153068 28432 153074 28444
rect 271874 28432 271880 28444
rect 271932 28432 271938 28484
rect 150434 28364 150440 28416
rect 150492 28404 150498 28416
rect 371234 28404 371240 28416
rect 150492 28376 371240 28404
rect 150492 28364 150498 28376
rect 371234 28364 371240 28376
rect 371292 28364 371298 28416
rect 152826 28296 152832 28348
rect 152884 28336 152890 28348
rect 375374 28336 375380 28348
rect 152884 28308 375380 28336
rect 152884 28296 152890 28308
rect 375374 28296 375380 28308
rect 375432 28296 375438 28348
rect 165982 28228 165988 28280
rect 166040 28268 166046 28280
rect 571334 28268 571340 28280
rect 166040 28240 571340 28268
rect 166040 28228 166046 28240
rect 571334 28228 571340 28240
rect 571392 28228 571398 28280
rect 138290 28160 138296 28212
rect 138348 28200 138354 28212
rect 215294 28200 215300 28212
rect 138348 28172 215300 28200
rect 138348 28160 138354 28172
rect 215294 28160 215300 28172
rect 215352 28160 215358 28212
rect 138106 28092 138112 28144
rect 138164 28132 138170 28144
rect 211154 28132 211160 28144
rect 138164 28104 211160 28132
rect 138164 28092 138170 28104
rect 211154 28092 211160 28104
rect 211212 28092 211218 28144
rect 150158 28024 150164 28076
rect 150216 28064 150222 28076
rect 222194 28064 222200 28076
rect 150216 28036 222200 28064
rect 150216 28024 150222 28036
rect 222194 28024 222200 28036
rect 222252 28024 222258 28076
rect 143258 27548 143264 27600
rect 143316 27588 143322 27600
rect 193214 27588 193220 27600
rect 143316 27560 193220 27588
rect 143316 27548 143322 27560
rect 193214 27548 193220 27560
rect 193272 27548 193278 27600
rect 136082 27480 136088 27532
rect 136140 27520 136146 27532
rect 186314 27520 186320 27532
rect 136140 27492 186320 27520
rect 136140 27480 136146 27492
rect 186314 27480 186320 27492
rect 186372 27480 186378 27532
rect 136910 27412 136916 27464
rect 136968 27452 136974 27464
rect 197354 27452 197360 27464
rect 136968 27424 197360 27452
rect 136968 27412 136974 27424
rect 197354 27412 197360 27424
rect 197412 27412 197418 27464
rect 146018 27344 146024 27396
rect 146076 27384 146082 27396
rect 208394 27384 208400 27396
rect 146076 27356 208400 27384
rect 146076 27344 146082 27356
rect 208394 27344 208400 27356
rect 208452 27344 208458 27396
rect 137186 27276 137192 27328
rect 137244 27316 137250 27328
rect 201494 27316 201500 27328
rect 137244 27288 201500 27316
rect 137244 27276 137250 27288
rect 201494 27276 201500 27288
rect 201552 27276 201558 27328
rect 137462 27208 137468 27260
rect 137520 27248 137526 27260
rect 204254 27248 204260 27260
rect 137520 27220 204260 27248
rect 137520 27208 137526 27220
rect 204254 27208 204260 27220
rect 204312 27208 204318 27260
rect 138566 27140 138572 27192
rect 138624 27180 138630 27192
rect 218054 27180 218060 27192
rect 138624 27152 218060 27180
rect 138624 27140 138630 27152
rect 218054 27140 218060 27152
rect 218112 27140 218118 27192
rect 139670 27072 139676 27124
rect 139728 27112 139734 27124
rect 233234 27112 233240 27124
rect 139728 27084 233240 27112
rect 139728 27072 139734 27084
rect 233234 27072 233240 27084
rect 233292 27072 233298 27124
rect 148318 27004 148324 27056
rect 148376 27044 148382 27056
rect 343634 27044 343640 27056
rect 148376 27016 343640 27044
rect 148376 27004 148382 27016
rect 343634 27004 343640 27016
rect 343692 27004 343698 27056
rect 154574 26936 154580 26988
rect 154632 26976 154638 26988
rect 423674 26976 423680 26988
rect 154632 26948 423680 26976
rect 154632 26936 154638 26948
rect 423674 26936 423680 26948
rect 423732 26936 423738 26988
rect 157978 26868 157984 26920
rect 158036 26908 158042 26920
rect 467834 26908 467840 26920
rect 158036 26880 467840 26908
rect 158036 26868 158042 26880
rect 467834 26868 467840 26880
rect 467892 26868 467898 26920
rect 135806 26188 135812 26240
rect 135864 26228 135870 26240
rect 183554 26228 183560 26240
rect 135864 26200 183560 26228
rect 135864 26188 135870 26200
rect 183554 26188 183560 26200
rect 183612 26188 183618 26240
rect 139946 26120 139952 26172
rect 140004 26160 140010 26172
rect 235994 26160 236000 26172
rect 140004 26132 236000 26160
rect 140004 26120 140010 26132
rect 235994 26120 236000 26132
rect 236052 26120 236058 26172
rect 141878 26052 141884 26104
rect 141936 26092 141942 26104
rect 260834 26092 260840 26104
rect 141936 26064 260840 26092
rect 141936 26052 141942 26064
rect 260834 26052 260840 26064
rect 260892 26052 260898 26104
rect 144362 25984 144368 26036
rect 144420 26024 144426 26036
rect 292574 26024 292580 26036
rect 144420 25996 292580 26024
rect 144420 25984 144426 25996
rect 292574 25984 292580 25996
rect 292632 25984 292638 26036
rect 149330 25916 149336 25968
rect 149388 25956 149394 25968
rect 357526 25956 357532 25968
rect 149388 25928 357532 25956
rect 149388 25916 149394 25928
rect 357526 25916 357532 25928
rect 357584 25916 357590 25968
rect 150526 25848 150532 25900
rect 150584 25888 150590 25900
rect 372614 25888 372620 25900
rect 150584 25860 372620 25888
rect 150584 25848 150590 25860
rect 372614 25848 372620 25860
rect 372672 25848 372678 25900
rect 153746 25780 153752 25832
rect 153804 25820 153810 25832
rect 414014 25820 414020 25832
rect 153804 25792 414020 25820
rect 153804 25780 153810 25792
rect 414014 25780 414020 25792
rect 414072 25780 414078 25832
rect 164786 25712 164792 25764
rect 164844 25752 164850 25764
rect 556154 25752 556160 25764
rect 164844 25724 556160 25752
rect 164844 25712 164850 25724
rect 556154 25712 556160 25724
rect 556212 25712 556218 25764
rect 166626 25644 166632 25696
rect 166684 25684 166690 25696
rect 558914 25684 558920 25696
rect 166684 25656 558920 25684
rect 166684 25644 166690 25656
rect 558914 25644 558920 25656
rect 558972 25644 558978 25696
rect 165614 25576 165620 25628
rect 165672 25616 165678 25628
rect 565814 25616 565820 25628
rect 165672 25588 565820 25616
rect 165672 25576 165678 25588
rect 565814 25576 565820 25588
rect 565872 25576 565878 25628
rect 81434 25508 81440 25560
rect 81492 25548 81498 25560
rect 120902 25548 120908 25560
rect 81492 25520 120908 25548
rect 81492 25508 81498 25520
rect 120902 25508 120908 25520
rect 120960 25508 120966 25560
rect 166166 25508 166172 25560
rect 166224 25548 166230 25560
rect 572714 25548 572720 25560
rect 166224 25520 572720 25548
rect 166224 25508 166230 25520
rect 572714 25508 572720 25520
rect 572772 25508 572778 25560
rect 135530 25440 135536 25492
rect 135588 25480 135594 25492
rect 179414 25480 179420 25492
rect 135588 25452 179420 25480
rect 135588 25440 135594 25452
rect 179414 25440 179420 25452
rect 179472 25440 179478 25492
rect 135254 25372 135260 25424
rect 135312 25412 135318 25424
rect 176746 25412 176752 25424
rect 135312 25384 176752 25412
rect 135312 25372 135318 25384
rect 176746 25372 176752 25384
rect 176804 25372 176810 25424
rect 141326 24760 141332 24812
rect 141384 24800 141390 24812
rect 253934 24800 253940 24812
rect 141384 24772 253940 24800
rect 141384 24760 141390 24772
rect 253934 24760 253940 24772
rect 253992 24760 253998 24812
rect 143534 24692 143540 24744
rect 143592 24732 143598 24744
rect 282914 24732 282920 24744
rect 143592 24704 282920 24732
rect 143592 24692 143598 24704
rect 282914 24692 282920 24704
rect 282972 24692 282978 24744
rect 153194 24624 153200 24676
rect 153252 24664 153258 24676
rect 407206 24664 407212 24676
rect 153252 24636 407212 24664
rect 153252 24624 153258 24636
rect 407206 24624 407212 24636
rect 407264 24624 407270 24676
rect 162854 24556 162860 24608
rect 162912 24596 162918 24608
rect 531314 24596 531320 24608
rect 162912 24568 531320 24596
rect 162912 24556 162918 24568
rect 531314 24556 531320 24568
rect 531372 24556 531378 24608
rect 163130 24488 163136 24540
rect 163188 24528 163194 24540
rect 534074 24528 534080 24540
rect 163188 24500 534080 24528
rect 163188 24488 163194 24500
rect 534074 24488 534080 24500
rect 534132 24488 534138 24540
rect 163406 24420 163412 24472
rect 163464 24460 163470 24472
rect 538214 24460 538220 24472
rect 163464 24432 538220 24460
rect 163464 24420 163470 24432
rect 538214 24420 538220 24432
rect 538272 24420 538278 24472
rect 163682 24352 163688 24404
rect 163740 24392 163746 24404
rect 540974 24392 540980 24404
rect 163740 24364 540980 24392
rect 163740 24352 163746 24364
rect 540974 24352 540980 24364
rect 541032 24352 541038 24404
rect 164234 24284 164240 24336
rect 164292 24324 164298 24336
rect 547874 24324 547880 24336
rect 164292 24296 547880 24324
rect 164292 24284 164298 24296
rect 547874 24284 547880 24296
rect 547932 24284 547938 24336
rect 164510 24216 164516 24268
rect 164568 24256 164574 24268
rect 552014 24256 552020 24268
rect 164568 24228 552020 24256
rect 164568 24216 164574 24228
rect 552014 24216 552020 24228
rect 552072 24216 552078 24268
rect 165706 24148 165712 24200
rect 165764 24188 165770 24200
rect 567194 24188 567200 24200
rect 165764 24160 567200 24188
rect 165764 24148 165770 24160
rect 567194 24148 567200 24160
rect 567252 24148 567258 24200
rect 165890 24080 165896 24132
rect 165948 24120 165954 24132
rect 569954 24120 569960 24132
rect 165948 24092 569960 24120
rect 165948 24080 165954 24092
rect 569954 24080 569960 24092
rect 570012 24080 570018 24132
rect 157334 23400 157340 23452
rect 157392 23440 157398 23452
rect 459554 23440 459560 23452
rect 157392 23412 459560 23440
rect 157392 23400 157398 23412
rect 459554 23400 459560 23412
rect 459612 23400 459618 23452
rect 160094 23332 160100 23384
rect 160152 23372 160158 23384
rect 495434 23372 495440 23384
rect 160152 23344 495440 23372
rect 160152 23332 160158 23344
rect 495434 23332 495440 23344
rect 495492 23332 495498 23384
rect 160370 23264 160376 23316
rect 160428 23304 160434 23316
rect 498286 23304 498292 23316
rect 160428 23276 498292 23304
rect 160428 23264 160434 23276
rect 498286 23264 498292 23276
rect 498344 23264 498350 23316
rect 160646 23196 160652 23248
rect 160704 23236 160710 23248
rect 502334 23236 502340 23248
rect 160704 23208 502340 23236
rect 160704 23196 160710 23208
rect 502334 23196 502340 23208
rect 502392 23196 502398 23248
rect 160922 23128 160928 23180
rect 160980 23168 160986 23180
rect 506474 23168 506480 23180
rect 160980 23140 506480 23168
rect 160980 23128 160986 23140
rect 506474 23128 506480 23140
rect 506532 23128 506538 23180
rect 161474 23060 161480 23112
rect 161532 23100 161538 23112
rect 513374 23100 513380 23112
rect 161532 23072 513380 23100
rect 161532 23060 161538 23072
rect 513374 23060 513380 23072
rect 513432 23060 513438 23112
rect 161750 22992 161756 23044
rect 161808 23032 161814 23044
rect 516134 23032 516140 23044
rect 161808 23004 516140 23032
rect 161808 22992 161814 23004
rect 516134 22992 516140 23004
rect 516192 22992 516198 23044
rect 162026 22924 162032 22976
rect 162084 22964 162090 22976
rect 520274 22964 520280 22976
rect 162084 22936 520280 22964
rect 162084 22924 162090 22936
rect 520274 22924 520280 22936
rect 520332 22924 520338 22976
rect 162302 22856 162308 22908
rect 162360 22896 162366 22908
rect 523034 22896 523040 22908
rect 162360 22868 523040 22896
rect 162360 22856 162366 22868
rect 523034 22856 523040 22868
rect 523092 22856 523098 22908
rect 165154 22788 165160 22840
rect 165212 22828 165218 22840
rect 560294 22828 560300 22840
rect 165212 22800 560300 22828
rect 165212 22788 165218 22800
rect 560294 22788 560300 22800
rect 560352 22788 560358 22840
rect 114462 22720 114468 22772
rect 114520 22760 114526 22772
rect 580166 22760 580172 22772
rect 114520 22732 580172 22760
rect 114520 22720 114526 22732
rect 580166 22720 580172 22732
rect 580224 22720 580230 22772
rect 3510 22652 3516 22704
rect 3568 22692 3574 22704
rect 170306 22692 170312 22704
rect 3568 22664 170312 22692
rect 3568 22652 3574 22664
rect 170306 22652 170312 22664
rect 170364 22652 170370 22704
rect 148042 21972 148048 22024
rect 148100 22012 148106 22024
rect 340874 22012 340880 22024
rect 148100 21984 340880 22012
rect 148100 21972 148106 21984
rect 340874 21972 340880 21984
rect 340932 21972 340938 22024
rect 156874 21904 156880 21956
rect 156932 21944 156938 21956
rect 361574 21944 361580 21956
rect 156932 21916 361580 21944
rect 156932 21904 156938 21916
rect 361574 21904 361580 21916
rect 361632 21904 361638 21956
rect 155034 21836 155040 21888
rect 155092 21876 155098 21888
rect 430574 21876 430580 21888
rect 155092 21848 430580 21876
rect 155092 21836 155098 21848
rect 430574 21836 430580 21848
rect 430632 21836 430638 21888
rect 155218 21768 155224 21820
rect 155276 21808 155282 21820
rect 432046 21808 432052 21820
rect 155276 21780 432052 21808
rect 155276 21768 155282 21780
rect 432046 21768 432052 21780
rect 432104 21768 432110 21820
rect 156322 21700 156328 21752
rect 156380 21740 156386 21752
rect 447134 21740 447140 21752
rect 156380 21712 447140 21740
rect 156380 21700 156386 21712
rect 447134 21700 447140 21712
rect 447192 21700 447198 21752
rect 156414 21632 156420 21684
rect 156472 21672 156478 21684
rect 448514 21672 448520 21684
rect 156472 21644 448520 21672
rect 156472 21632 156478 21644
rect 448514 21632 448520 21644
rect 448572 21632 448578 21684
rect 158990 21564 158996 21616
rect 159048 21604 159054 21616
rect 481726 21604 481732 21616
rect 159048 21576 481732 21604
rect 159048 21564 159054 21576
rect 481726 21564 481732 21576
rect 481784 21564 481790 21616
rect 159266 21496 159272 21548
rect 159324 21536 159330 21548
rect 484394 21536 484400 21548
rect 159324 21508 484400 21536
rect 159324 21496 159330 21508
rect 484394 21496 484400 21508
rect 484452 21496 484458 21548
rect 159542 21428 159548 21480
rect 159600 21468 159606 21480
rect 488534 21468 488540 21480
rect 159600 21440 488540 21468
rect 159600 21428 159606 21440
rect 488534 21428 488540 21440
rect 488592 21428 488598 21480
rect 159818 21360 159824 21412
rect 159876 21400 159882 21412
rect 491294 21400 491300 21412
rect 159876 21372 491300 21400
rect 159876 21360 159882 21372
rect 491294 21360 491300 21372
rect 491352 21360 491358 21412
rect 140038 20408 140044 20460
rect 140096 20448 140102 20460
rect 237374 20448 237380 20460
rect 140096 20420 237380 20448
rect 140096 20408 140102 20420
rect 237374 20408 237380 20420
rect 237432 20408 237438 20460
rect 141694 20340 141700 20392
rect 141752 20380 141758 20392
rect 259546 20380 259552 20392
rect 141752 20352 259552 20380
rect 141752 20340 141758 20352
rect 259546 20340 259552 20352
rect 259604 20340 259610 20392
rect 147214 20272 147220 20324
rect 147272 20312 147278 20324
rect 329834 20312 329840 20324
rect 147272 20284 329840 20312
rect 147272 20272 147278 20284
rect 329834 20272 329840 20284
rect 329892 20272 329898 20324
rect 139486 20204 139492 20256
rect 139544 20244 139550 20256
rect 230474 20244 230480 20256
rect 139544 20216 230480 20244
rect 139544 20204 139550 20216
rect 230474 20204 230480 20216
rect 230532 20204 230538 20256
rect 231118 20204 231124 20256
rect 231176 20244 231182 20256
rect 449894 20244 449900 20256
rect 231176 20216 449900 20244
rect 231176 20204 231182 20216
rect 449894 20204 449900 20216
rect 449952 20204 449958 20256
rect 152274 20136 152280 20188
rect 152332 20176 152338 20188
rect 394694 20176 394700 20188
rect 152332 20148 394700 20176
rect 152332 20136 152338 20148
rect 394694 20136 394700 20148
rect 394752 20136 394758 20188
rect 152550 20068 152556 20120
rect 152608 20108 152614 20120
rect 398834 20108 398840 20120
rect 152608 20080 398840 20108
rect 152608 20068 152614 20080
rect 398834 20068 398840 20080
rect 398892 20068 398898 20120
rect 153654 20000 153660 20052
rect 153712 20040 153718 20052
rect 412634 20040 412640 20052
rect 153712 20012 412640 20040
rect 153712 20000 153718 20012
rect 412634 20000 412640 20012
rect 412692 20000 412698 20052
rect 158070 19932 158076 19984
rect 158128 19972 158134 19984
rect 469214 19972 469220 19984
rect 158128 19944 469220 19972
rect 158128 19932 158134 19944
rect 469214 19932 469220 19944
rect 469272 19932 469278 19984
rect 141142 19048 141148 19100
rect 141200 19088 141206 19100
rect 251266 19088 251272 19100
rect 141200 19060 251272 19088
rect 141200 19048 141206 19060
rect 251266 19048 251272 19060
rect 251324 19048 251330 19100
rect 163774 18980 163780 19032
rect 163832 19020 163838 19032
rect 312538 19020 312544 19032
rect 163832 18992 312544 19020
rect 163832 18980 163838 18992
rect 312538 18980 312544 18992
rect 312596 18980 312602 19032
rect 149514 18912 149520 18964
rect 149572 18952 149578 18964
rect 358814 18952 358820 18964
rect 149572 18924 358820 18952
rect 149572 18912 149578 18924
rect 358814 18912 358820 18924
rect 358872 18912 358878 18964
rect 150894 18844 150900 18896
rect 150952 18884 150958 18896
rect 376754 18884 376760 18896
rect 150952 18856 376760 18884
rect 150952 18844 150958 18856
rect 376754 18844 376760 18856
rect 376812 18844 376818 18896
rect 151170 18776 151176 18828
rect 151228 18816 151234 18828
rect 380894 18816 380900 18828
rect 151228 18788 380900 18816
rect 151228 18776 151234 18788
rect 380894 18776 380900 18788
rect 380952 18776 380958 18828
rect 156690 18708 156696 18760
rect 156748 18748 156754 18760
rect 451274 18748 451280 18760
rect 156748 18720 451280 18748
rect 156748 18708 156754 18720
rect 451274 18708 451280 18720
rect 451332 18708 451338 18760
rect 163222 18640 163228 18692
rect 163280 18680 163286 18692
rect 535454 18680 535460 18692
rect 163280 18652 535460 18680
rect 163280 18640 163286 18652
rect 535454 18640 535460 18652
rect 535512 18640 535518 18692
rect 35894 18572 35900 18624
rect 35952 18612 35958 18624
rect 118142 18612 118148 18624
rect 35952 18584 118148 18612
rect 35952 18572 35958 18584
rect 118142 18572 118148 18584
rect 118200 18572 118206 18624
rect 164602 18572 164608 18624
rect 164660 18612 164666 18624
rect 553394 18612 553400 18624
rect 164660 18584 553400 18612
rect 164660 18572 164666 18584
rect 553394 18572 553400 18584
rect 553452 18572 553458 18624
rect 142798 17620 142804 17672
rect 142856 17660 142862 17672
rect 273254 17660 273260 17672
rect 142856 17632 273260 17660
rect 142856 17620 142862 17632
rect 273254 17620 273260 17632
rect 273312 17620 273318 17672
rect 147030 17552 147036 17604
rect 147088 17592 147094 17604
rect 327074 17592 327080 17604
rect 147088 17564 327080 17592
rect 147088 17552 147094 17564
rect 327074 17552 327080 17564
rect 327132 17552 327138 17604
rect 154850 17484 154856 17536
rect 154908 17524 154914 17536
rect 427814 17524 427820 17536
rect 154908 17496 427820 17524
rect 154908 17484 154914 17496
rect 427814 17484 427820 17496
rect 427872 17484 427878 17536
rect 155310 17416 155316 17468
rect 155368 17456 155374 17468
rect 433334 17456 433340 17468
rect 155368 17428 433340 17456
rect 155368 17416 155374 17428
rect 433334 17416 433340 17428
rect 433392 17416 433398 17468
rect 155402 17348 155408 17400
rect 155460 17388 155466 17400
rect 434714 17388 434720 17400
rect 155460 17360 434720 17388
rect 155460 17348 155466 17360
rect 434714 17348 434720 17360
rect 434772 17348 434778 17400
rect 155586 17280 155592 17332
rect 155644 17320 155650 17332
rect 437474 17320 437480 17332
rect 155644 17292 437480 17320
rect 155644 17280 155650 17292
rect 437474 17280 437480 17292
rect 437532 17280 437538 17332
rect 164878 17212 164884 17264
rect 164936 17252 164942 17264
rect 556246 17252 556252 17264
rect 164936 17224 556252 17252
rect 164936 17212 164942 17224
rect 556246 17212 556252 17224
rect 556304 17212 556310 17264
rect 142890 16396 142896 16448
rect 142948 16436 142954 16448
rect 274818 16436 274824 16448
rect 142948 16408 274824 16436
rect 142948 16396 142954 16408
rect 274818 16396 274824 16408
rect 274876 16396 274882 16448
rect 143902 16328 143908 16380
rect 143960 16368 143966 16380
rect 287330 16368 287336 16380
rect 143960 16340 287336 16368
rect 143960 16328 143966 16340
rect 287330 16328 287336 16340
rect 287388 16328 287394 16380
rect 143994 16260 144000 16312
rect 144052 16300 144058 16312
rect 288986 16300 288992 16312
rect 144052 16272 288992 16300
rect 144052 16260 144058 16272
rect 288986 16260 288992 16272
rect 289044 16260 289050 16312
rect 144270 16192 144276 16244
rect 144328 16232 144334 16244
rect 292666 16232 292672 16244
rect 144328 16204 292672 16232
rect 144328 16192 144334 16204
rect 292666 16192 292672 16204
rect 292724 16192 292730 16244
rect 148502 16124 148508 16176
rect 148560 16164 148566 16176
rect 346946 16164 346952 16176
rect 148560 16136 346952 16164
rect 148560 16124 148566 16136
rect 346946 16124 346952 16136
rect 347004 16124 347010 16176
rect 149054 16056 149060 16108
rect 149112 16096 149118 16108
rect 353570 16096 353576 16108
rect 149112 16068 353576 16096
rect 149112 16056 149118 16068
rect 353570 16056 353576 16068
rect 353628 16056 353634 16108
rect 153930 15988 153936 16040
rect 153988 16028 153994 16040
rect 415486 16028 415492 16040
rect 153988 16000 415492 16028
rect 153988 15988 153994 16000
rect 415486 15988 415492 16000
rect 415544 15988 415550 16040
rect 171778 15920 171784 15972
rect 171836 15960 171842 15972
rect 443362 15960 443368 15972
rect 171836 15932 443368 15960
rect 171836 15920 171842 15932
rect 443362 15920 443368 15932
rect 443420 15920 443426 15972
rect 162946 15852 162952 15904
rect 163004 15892 163010 15904
rect 532050 15892 532056 15904
rect 163004 15864 532056 15892
rect 163004 15852 163010 15864
rect 532050 15852 532056 15864
rect 532108 15852 532114 15904
rect 141234 14900 141240 14952
rect 141292 14940 141298 14952
rect 253474 14940 253480 14952
rect 141292 14912 253480 14940
rect 141292 14900 141298 14912
rect 253474 14900 253480 14912
rect 253532 14900 253538 14952
rect 141510 14832 141516 14884
rect 141568 14872 141574 14884
rect 256694 14872 256700 14884
rect 141568 14844 256700 14872
rect 141568 14832 141574 14844
rect 256694 14832 256700 14844
rect 256752 14832 256758 14884
rect 142338 14764 142344 14816
rect 142396 14804 142402 14816
rect 267734 14804 267740 14816
rect 142396 14776 267740 14804
rect 142396 14764 142402 14776
rect 267734 14764 267740 14776
rect 267792 14764 267798 14816
rect 142614 14696 142620 14748
rect 142672 14736 142678 14748
rect 270770 14736 270776 14748
rect 142672 14708 270776 14736
rect 142672 14696 142678 14708
rect 270770 14696 270776 14708
rect 270828 14696 270834 14748
rect 149606 14628 149612 14680
rect 149664 14668 149670 14680
rect 361114 14668 361120 14680
rect 149664 14640 361120 14668
rect 149664 14628 149670 14640
rect 361114 14628 361120 14640
rect 361172 14628 361178 14680
rect 151446 14560 151452 14612
rect 151504 14600 151510 14612
rect 384298 14600 384304 14612
rect 151504 14572 384304 14600
rect 151504 14560 151510 14572
rect 384298 14560 384304 14572
rect 384356 14560 384362 14612
rect 154666 14492 154672 14544
rect 154724 14532 154730 14544
rect 425698 14532 425704 14544
rect 154724 14504 425704 14532
rect 154724 14492 154730 14504
rect 425698 14492 425704 14504
rect 425756 14492 425762 14544
rect 157886 14424 157892 14476
rect 157944 14464 157950 14476
rect 467466 14464 467472 14476
rect 157944 14436 467472 14464
rect 157944 14424 157950 14436
rect 467466 14424 467472 14436
rect 467524 14424 467530 14476
rect 139578 13404 139584 13456
rect 139636 13444 139642 13456
rect 231854 13444 231860 13456
rect 139636 13416 231860 13444
rect 139636 13404 139642 13416
rect 231854 13404 231860 13416
rect 231912 13404 231918 13456
rect 140130 13336 140136 13388
rect 140188 13376 140194 13388
rect 239306 13376 239312 13388
rect 140188 13348 239312 13376
rect 140188 13336 140194 13348
rect 239306 13336 239312 13348
rect 239364 13336 239370 13388
rect 146846 13268 146852 13320
rect 146904 13308 146910 13320
rect 324406 13308 324412 13320
rect 146904 13280 324412 13308
rect 146904 13268 146910 13280
rect 324406 13268 324412 13280
rect 324464 13268 324470 13320
rect 147122 13200 147128 13252
rect 147180 13240 147186 13252
rect 328730 13240 328736 13252
rect 147180 13212 328736 13240
rect 147180 13200 147186 13212
rect 328730 13200 328736 13212
rect 328788 13200 328794 13252
rect 149790 13132 149796 13184
rect 149848 13172 149854 13184
rect 363506 13172 363512 13184
rect 149848 13144 363512 13172
rect 149848 13132 149854 13144
rect 363506 13132 363512 13144
rect 363564 13132 363570 13184
rect 14274 13064 14280 13116
rect 14332 13104 14338 13116
rect 122098 13104 122104 13116
rect 14332 13076 122104 13104
rect 14332 13064 14338 13076
rect 122098 13064 122104 13076
rect 122156 13064 122162 13116
rect 150986 13064 150992 13116
rect 151044 13104 151050 13116
rect 378410 13104 378416 13116
rect 151044 13076 378416 13104
rect 151044 13064 151050 13076
rect 378410 13064 378416 13076
rect 378468 13064 378474 13116
rect 157702 12248 157708 12300
rect 157760 12288 157766 12300
rect 169110 12288 169116 12300
rect 157760 12260 169116 12288
rect 157760 12248 157766 12260
rect 169110 12248 169116 12260
rect 169168 12248 169174 12300
rect 138198 12180 138204 12232
rect 138256 12220 138262 12232
rect 214466 12220 214472 12232
rect 138256 12192 214472 12220
rect 138256 12180 138262 12192
rect 214466 12180 214472 12192
rect 214524 12180 214530 12232
rect 138474 12112 138480 12164
rect 138532 12152 138538 12164
rect 218146 12152 218152 12164
rect 138532 12124 218152 12152
rect 138532 12112 138538 12124
rect 218146 12112 218152 12124
rect 218204 12112 218210 12164
rect 138750 12044 138756 12096
rect 138808 12084 138814 12096
rect 221090 12084 221096 12096
rect 138808 12056 221096 12084
rect 138808 12044 138814 12056
rect 221090 12044 221096 12056
rect 221148 12044 221154 12096
rect 146570 11976 146576 12028
rect 146628 12016 146634 12028
rect 322106 12016 322112 12028
rect 146628 11988 322112 12016
rect 146628 11976 146634 11988
rect 322106 11976 322112 11988
rect 322164 11976 322170 12028
rect 148226 11908 148232 11960
rect 148284 11948 148290 11960
rect 342898 11948 342904 11960
rect 148284 11920 342904 11948
rect 148284 11908 148290 11920
rect 342898 11908 342904 11920
rect 342956 11908 342962 11960
rect 148410 11840 148416 11892
rect 148468 11880 148474 11892
rect 345290 11880 345296 11892
rect 148468 11852 345296 11880
rect 148468 11840 148474 11852
rect 345290 11840 345296 11852
rect 345348 11840 345354 11892
rect 149238 11772 149244 11824
rect 149296 11812 149302 11824
rect 356330 11812 356336 11824
rect 149296 11784 356336 11812
rect 149296 11772 149302 11784
rect 356330 11772 356336 11784
rect 356388 11772 356394 11824
rect 159358 11704 159364 11756
rect 159416 11744 159422 11756
rect 486418 11744 486424 11756
rect 159416 11716 486424 11744
rect 159416 11704 159422 11716
rect 486418 11704 486424 11716
rect 486476 11704 486482 11756
rect 176654 11636 176660 11688
rect 176712 11676 176718 11688
rect 177850 11676 177856 11688
rect 176712 11648 177856 11676
rect 176712 11636 176718 11648
rect 177850 11636 177856 11648
rect 177908 11636 177914 11688
rect 218054 11636 218060 11688
rect 218112 11676 218118 11688
rect 219250 11676 219256 11688
rect 218112 11648 219256 11676
rect 218112 11636 218118 11648
rect 219250 11636 219256 11648
rect 219308 11636 219314 11688
rect 242894 11636 242900 11688
rect 242952 11676 242958 11688
rect 244090 11676 244096 11688
rect 242952 11648 244096 11676
rect 242952 11636 242958 11648
rect 244090 11636 244096 11648
rect 244148 11636 244154 11688
rect 259454 11636 259460 11688
rect 259512 11676 259518 11688
rect 260650 11676 260656 11688
rect 259512 11648 260656 11676
rect 259512 11636 259518 11648
rect 260650 11636 260656 11648
rect 260708 11636 260714 11688
rect 110506 10956 110512 11008
rect 110564 10996 110570 11008
rect 130470 10996 130476 11008
rect 110564 10968 130476 10996
rect 110564 10956 110570 10968
rect 130470 10956 130476 10968
rect 130528 10956 130534 11008
rect 102134 10888 102140 10940
rect 102192 10928 102198 10940
rect 128998 10928 129004 10940
rect 102192 10900 129004 10928
rect 102192 10888 102198 10900
rect 128998 10888 129004 10900
rect 129056 10888 129062 10940
rect 95786 10820 95792 10872
rect 95844 10860 95850 10872
rect 129182 10860 129188 10872
rect 95844 10832 129188 10860
rect 95844 10820 95850 10832
rect 129182 10820 129188 10832
rect 129240 10820 129246 10872
rect 134794 10820 134800 10872
rect 134852 10860 134858 10872
rect 170306 10860 170312 10872
rect 134852 10832 170312 10860
rect 134852 10820 134858 10832
rect 170306 10820 170312 10832
rect 170364 10820 170370 10872
rect 92474 10752 92480 10804
rect 92532 10792 92538 10804
rect 129090 10792 129096 10804
rect 92532 10764 129096 10792
rect 92532 10752 92538 10764
rect 129090 10752 129096 10764
rect 129148 10752 129154 10804
rect 137094 10752 137100 10804
rect 137152 10792 137158 10804
rect 200298 10792 200304 10804
rect 137152 10764 200304 10792
rect 137152 10752 137158 10764
rect 200298 10752 200304 10764
rect 200356 10752 200362 10804
rect 74994 10684 75000 10736
rect 75052 10724 75058 10736
rect 122190 10724 122196 10736
rect 75052 10696 122196 10724
rect 75052 10684 75058 10696
rect 122190 10684 122196 10696
rect 122248 10684 122254 10736
rect 137370 10684 137376 10736
rect 137428 10724 137434 10736
rect 203426 10724 203432 10736
rect 137428 10696 203432 10724
rect 137428 10684 137434 10696
rect 203426 10684 203432 10696
rect 203484 10684 203490 10736
rect 78122 10616 78128 10668
rect 78180 10656 78186 10668
rect 127802 10656 127808 10668
rect 78180 10628 127808 10656
rect 78180 10616 78186 10628
rect 127802 10616 127808 10628
rect 127860 10616 127866 10668
rect 142982 10616 142988 10668
rect 143040 10656 143046 10668
rect 276106 10656 276112 10668
rect 143040 10628 276112 10656
rect 143040 10616 143046 10628
rect 276106 10616 276112 10628
rect 276164 10616 276170 10668
rect 67634 10548 67640 10600
rect 67692 10588 67698 10600
rect 126330 10588 126336 10600
rect 67692 10560 126336 10588
rect 67692 10548 67698 10560
rect 126330 10548 126336 10560
rect 126388 10548 126394 10600
rect 144454 10548 144460 10600
rect 144512 10588 144518 10600
rect 294874 10588 294880 10600
rect 144512 10560 294880 10588
rect 144512 10548 144518 10560
rect 294874 10548 294880 10560
rect 294932 10548 294938 10600
rect 64322 10480 64328 10532
rect 64380 10520 64386 10532
rect 126422 10520 126428 10532
rect 64380 10492 126428 10520
rect 64380 10480 64386 10492
rect 126422 10480 126428 10492
rect 126480 10480 126486 10532
rect 145926 10480 145932 10532
rect 145984 10520 145990 10532
rect 313826 10520 313832 10532
rect 145984 10492 313832 10520
rect 145984 10480 145990 10492
rect 313826 10480 313832 10492
rect 313884 10480 313890 10532
rect 46658 10412 46664 10464
rect 46716 10452 46722 10464
rect 125042 10452 125048 10464
rect 46716 10424 125048 10452
rect 46716 10412 46722 10424
rect 125042 10412 125048 10424
rect 125100 10412 125106 10464
rect 146294 10412 146300 10464
rect 146352 10452 146358 10464
rect 318058 10452 318064 10464
rect 146352 10424 318064 10452
rect 146352 10412 146358 10424
rect 318058 10412 318064 10424
rect 318116 10412 318122 10464
rect 31938 10344 31944 10396
rect 31996 10384 32002 10396
rect 123662 10384 123668 10396
rect 31996 10356 123668 10384
rect 31996 10344 32002 10356
rect 123662 10344 123668 10356
rect 123720 10344 123726 10396
rect 152642 10344 152648 10396
rect 152700 10384 152706 10396
rect 398926 10384 398932 10396
rect 152700 10356 398932 10384
rect 152700 10344 152706 10356
rect 398926 10344 398932 10356
rect 398984 10344 398990 10396
rect 25314 10276 25320 10328
rect 25372 10316 25378 10328
rect 123570 10316 123576 10328
rect 25372 10288 123576 10316
rect 25372 10276 25378 10288
rect 123570 10276 123576 10288
rect 123628 10276 123634 10328
rect 156506 10276 156512 10328
rect 156564 10316 156570 10328
rect 448606 10316 448612 10328
rect 156564 10288 448612 10316
rect 156564 10276 156570 10288
rect 448606 10276 448612 10288
rect 448664 10276 448670 10328
rect 117314 10208 117320 10260
rect 117372 10248 117378 10260
rect 130378 10248 130384 10260
rect 117372 10220 130384 10248
rect 117372 10208 117378 10220
rect 130378 10208 130384 10220
rect 130436 10208 130442 10260
rect 120626 10140 120632 10192
rect 120684 10180 120690 10192
rect 130562 10180 130568 10192
rect 120684 10152 130568 10180
rect 120684 10140 120690 10152
rect 130562 10140 130568 10152
rect 130620 10140 130626 10192
rect 116394 9596 116400 9648
rect 116452 9636 116458 9648
rect 130194 9636 130200 9648
rect 116452 9608 130200 9636
rect 116452 9596 116458 9608
rect 130194 9596 130200 9608
rect 130252 9596 130258 9648
rect 135438 9596 135444 9648
rect 135496 9636 135502 9648
rect 179046 9636 179052 9648
rect 135496 9608 179052 9636
rect 135496 9596 135502 9608
rect 179046 9596 179052 9608
rect 179104 9596 179110 9648
rect 112806 9528 112812 9580
rect 112864 9568 112870 9580
rect 130286 9568 130292 9580
rect 112864 9540 130292 9568
rect 112864 9528 112870 9540
rect 130286 9528 130292 9540
rect 130344 9528 130350 9580
rect 135990 9528 135996 9580
rect 136048 9568 136054 9580
rect 186130 9568 186136 9580
rect 136048 9540 186136 9568
rect 136048 9528 136054 9540
rect 186130 9528 186136 9540
rect 186188 9528 186194 9580
rect 60826 9460 60832 9512
rect 60884 9500 60890 9512
rect 126146 9500 126152 9512
rect 60884 9472 126152 9500
rect 60884 9460 60890 9472
rect 126146 9460 126152 9472
rect 126204 9460 126210 9512
rect 145374 9460 145380 9512
rect 145432 9500 145438 9512
rect 306742 9500 306748 9512
rect 145432 9472 306748 9500
rect 145432 9460 145438 9472
rect 306742 9460 306748 9472
rect 306800 9460 306806 9512
rect 57238 9392 57244 9444
rect 57296 9432 57302 9444
rect 126238 9432 126244 9444
rect 57296 9404 126244 9432
rect 57296 9392 57302 9404
rect 126238 9392 126244 9404
rect 126296 9392 126302 9444
rect 145650 9392 145656 9444
rect 145708 9432 145714 9444
rect 310238 9432 310244 9444
rect 145708 9404 310244 9432
rect 145708 9392 145714 9404
rect 310238 9392 310244 9404
rect 310296 9392 310302 9444
rect 43070 9324 43076 9376
rect 43128 9364 43134 9376
rect 116670 9364 116676 9376
rect 43128 9336 116676 9364
rect 43128 9324 43134 9336
rect 116670 9324 116676 9336
rect 116728 9324 116734 9376
rect 145742 9324 145748 9376
rect 145800 9364 145806 9376
rect 311434 9364 311440 9376
rect 145800 9336 311440 9364
rect 145800 9324 145806 9336
rect 311434 9324 311440 9336
rect 311492 9324 311498 9376
rect 50154 9256 50160 9308
rect 50212 9296 50218 9308
rect 124858 9296 124864 9308
rect 50212 9268 124864 9296
rect 50212 9256 50218 9268
rect 124858 9256 124864 9268
rect 124916 9256 124922 9308
rect 147950 9256 147956 9308
rect 148008 9296 148014 9308
rect 339862 9296 339868 9308
rect 148008 9268 339868 9296
rect 148008 9256 148014 9268
rect 339862 9256 339868 9268
rect 339920 9256 339926 9308
rect 45462 9188 45468 9240
rect 45520 9228 45526 9240
rect 124766 9228 124772 9240
rect 45520 9200 124772 9228
rect 45520 9188 45526 9200
rect 124766 9188 124772 9200
rect 124824 9188 124830 9240
rect 148134 9188 148140 9240
rect 148192 9228 148198 9240
rect 342162 9228 342168 9240
rect 148192 9200 342168 9228
rect 148192 9188 148198 9200
rect 342162 9188 342168 9200
rect 342220 9188 342226 9240
rect 41874 9120 41880 9172
rect 41932 9160 41938 9172
rect 124950 9160 124956 9172
rect 41932 9132 124956 9160
rect 41932 9120 41938 9132
rect 124950 9120 124956 9132
rect 125008 9120 125014 9172
rect 152090 9120 152096 9172
rect 152148 9160 152154 9172
rect 393038 9160 393044 9172
rect 152148 9132 393044 9160
rect 152148 9120 152154 9132
rect 393038 9120 393044 9132
rect 393096 9120 393102 9172
rect 31294 9052 31300 9104
rect 31352 9092 31358 9104
rect 123386 9092 123392 9104
rect 31352 9064 123392 9092
rect 31352 9052 31358 9064
rect 123386 9052 123392 9064
rect 123444 9052 123450 9104
rect 153470 9052 153476 9104
rect 153528 9092 153534 9104
rect 410794 9092 410800 9104
rect 153528 9064 410800 9092
rect 153528 9052 153534 9064
rect 410794 9052 410800 9064
rect 410852 9052 410858 9104
rect 24210 8984 24216 9036
rect 24268 9024 24274 9036
rect 123478 9024 123484 9036
rect 24268 8996 123484 9024
rect 24268 8984 24274 8996
rect 123478 8984 123484 8996
rect 123536 8984 123542 9036
rect 153562 8984 153568 9036
rect 153620 9024 153626 9036
rect 411898 9024 411904 9036
rect 153620 8996 411904 9024
rect 153620 8984 153626 8996
rect 411898 8984 411904 8996
rect 411956 8984 411962 9036
rect 9950 8916 9956 8968
rect 10008 8956 10014 8968
rect 122006 8956 122012 8968
rect 10008 8928 122012 8956
rect 10008 8916 10014 8928
rect 122006 8916 122012 8928
rect 122064 8916 122070 8968
rect 166074 8916 166080 8968
rect 166132 8956 166138 8968
rect 572714 8956 572720 8968
rect 166132 8928 572720 8956
rect 166132 8916 166138 8928
rect 572714 8916 572720 8928
rect 572772 8916 572778 8968
rect 134886 8848 134892 8900
rect 134944 8888 134950 8900
rect 171962 8888 171968 8900
rect 134944 8860 171968 8888
rect 134944 8848 134950 8860
rect 171962 8848 171968 8860
rect 172020 8848 172026 8900
rect 98638 8236 98644 8288
rect 98696 8276 98702 8288
rect 128906 8276 128912 8288
rect 98696 8248 128912 8276
rect 98696 8236 98702 8248
rect 128906 8236 128912 8248
rect 128964 8236 128970 8288
rect 95142 8168 95148 8220
rect 95200 8208 95206 8220
rect 128814 8208 128820 8220
rect 95200 8180 128820 8208
rect 95200 8168 95206 8180
rect 128814 8168 128820 8180
rect 128872 8168 128878 8220
rect 84470 8100 84476 8152
rect 84528 8140 84534 8152
rect 127710 8140 127716 8152
rect 84528 8112 127716 8140
rect 84528 8100 84534 8112
rect 127710 8100 127716 8112
rect 127768 8100 127774 8152
rect 80882 8032 80888 8084
rect 80940 8072 80946 8084
rect 127434 8072 127440 8084
rect 80940 8044 127440 8072
rect 80940 8032 80946 8044
rect 127434 8032 127440 8044
rect 127492 8032 127498 8084
rect 77386 7964 77392 8016
rect 77444 8004 77450 8016
rect 127618 8004 127624 8016
rect 77444 7976 127624 8004
rect 77444 7964 77450 7976
rect 127618 7964 127624 7976
rect 127676 7964 127682 8016
rect 142430 7964 142436 8016
rect 142488 8004 142494 8016
rect 268838 8004 268844 8016
rect 142488 7976 268844 8004
rect 142488 7964 142494 7976
rect 268838 7964 268844 7976
rect 268896 7964 268902 8016
rect 73798 7896 73804 7948
rect 73856 7936 73862 7948
rect 127526 7936 127532 7948
rect 73856 7908 127532 7936
rect 73856 7896 73862 7908
rect 127526 7896 127532 7908
rect 127584 7896 127590 7948
rect 144086 7896 144092 7948
rect 144144 7936 144150 7948
rect 290182 7936 290188 7948
rect 144144 7908 290188 7936
rect 144144 7896 144150 7908
rect 290182 7896 290188 7908
rect 290240 7896 290246 7948
rect 66714 7828 66720 7880
rect 66772 7868 66778 7880
rect 125962 7868 125968 7880
rect 66772 7840 125968 7868
rect 66772 7828 66778 7840
rect 125962 7828 125968 7840
rect 126020 7828 126026 7880
rect 147674 7828 147680 7880
rect 147732 7868 147738 7880
rect 336274 7868 336280 7880
rect 147732 7840 336280 7868
rect 147732 7828 147738 7840
rect 336274 7828 336280 7840
rect 336332 7828 336338 7880
rect 63218 7760 63224 7812
rect 63276 7800 63282 7812
rect 126054 7800 126060 7812
rect 63276 7772 126060 7800
rect 63276 7760 63282 7772
rect 126054 7760 126060 7772
rect 126112 7760 126118 7812
rect 154022 7760 154028 7812
rect 154080 7800 154086 7812
rect 417878 7800 417884 7812
rect 154080 7772 417884 7800
rect 154080 7760 154086 7772
rect 417878 7760 417884 7772
rect 417936 7760 417942 7812
rect 27706 7692 27712 7744
rect 27764 7732 27770 7744
rect 123294 7732 123300 7744
rect 27764 7704 123300 7732
rect 27764 7692 27770 7704
rect 123294 7692 123300 7704
rect 123352 7692 123358 7744
rect 164694 7692 164700 7744
rect 164752 7732 164758 7744
rect 554958 7732 554964 7744
rect 164752 7704 554964 7732
rect 164752 7692 164758 7704
rect 554958 7692 554964 7704
rect 555016 7692 555022 7744
rect 19426 7624 19432 7676
rect 19484 7664 19490 7676
rect 118050 7664 118056 7676
rect 19484 7636 118056 7664
rect 19484 7624 19490 7636
rect 118050 7624 118056 7636
rect 118108 7624 118114 7676
rect 119890 7624 119896 7676
rect 119948 7664 119954 7676
rect 130102 7664 130108 7676
rect 119948 7636 130108 7664
rect 119948 7624 119954 7636
rect 130102 7624 130108 7636
rect 130160 7624 130166 7676
rect 164970 7624 164976 7676
rect 165028 7664 165034 7676
rect 558546 7664 558552 7676
rect 165028 7636 558552 7664
rect 165028 7624 165034 7636
rect 558546 7624 558552 7636
rect 558604 7624 558610 7676
rect 23014 7556 23020 7608
rect 23072 7596 23078 7608
rect 123202 7596 123208 7608
rect 23072 7568 123208 7596
rect 23072 7556 23078 7568
rect 123202 7556 123208 7568
rect 123260 7556 123266 7608
rect 165798 7556 165804 7608
rect 165856 7596 165862 7608
rect 569126 7596 569132 7608
rect 165856 7568 569132 7596
rect 165856 7556 165862 7568
rect 569126 7556 569132 7568
rect 569184 7556 569190 7608
rect 102226 7488 102232 7540
rect 102284 7528 102290 7540
rect 128722 7528 128728 7540
rect 102284 7500 128728 7528
rect 102284 7488 102290 7500
rect 128722 7488 128728 7500
rect 128780 7488 128786 7540
rect 481634 7488 481640 7540
rect 481692 7528 481698 7540
rect 482462 7528 482468 7540
rect 481692 7500 482468 7528
rect 481692 7488 481698 7500
rect 482462 7488 482468 7500
rect 482520 7488 482526 7540
rect 115198 6808 115204 6860
rect 115256 6848 115262 6860
rect 130010 6848 130016 6860
rect 115256 6820 130016 6848
rect 115256 6808 115262 6820
rect 130010 6808 130016 6820
rect 130068 6808 130074 6860
rect 562318 6808 562324 6860
rect 562376 6848 562382 6860
rect 580166 6848 580172 6860
rect 562376 6820 580172 6848
rect 562376 6808 562382 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 99834 6740 99840 6792
rect 99892 6780 99898 6792
rect 120810 6780 120816 6792
rect 99892 6752 120816 6780
rect 99892 6740 99898 6752
rect 120810 6740 120816 6752
rect 120868 6740 120874 6792
rect 59630 6672 59636 6724
rect 59688 6712 59694 6724
rect 125870 6712 125876 6724
rect 59688 6684 125876 6712
rect 59688 6672 59694 6684
rect 125870 6672 125876 6684
rect 125928 6672 125934 6724
rect 139854 6672 139860 6724
rect 139912 6712 139918 6724
rect 235810 6712 235816 6724
rect 139912 6684 235816 6712
rect 139912 6672 139918 6684
rect 235810 6672 235816 6684
rect 235868 6672 235874 6724
rect 11146 6604 11152 6656
rect 11204 6644 11210 6656
rect 86218 6644 86224 6656
rect 11204 6616 86224 6644
rect 11204 6604 11210 6616
rect 86218 6604 86224 6616
rect 86276 6604 86282 6656
rect 104526 6604 104532 6656
rect 104584 6644 104590 6656
rect 128630 6644 128636 6656
rect 104584 6616 128636 6644
rect 104584 6604 104590 6616
rect 128630 6604 128636 6616
rect 128688 6604 128694 6656
rect 143810 6604 143816 6656
rect 143868 6644 143874 6656
rect 286594 6644 286600 6656
rect 143868 6616 286600 6644
rect 143868 6604 143874 6616
rect 286594 6604 286600 6616
rect 286652 6604 286658 6656
rect 48958 6536 48964 6588
rect 49016 6576 49022 6588
rect 124490 6576 124496 6588
rect 49016 6548 124496 6576
rect 49016 6536 49022 6548
rect 124490 6536 124496 6548
rect 124548 6536 124554 6588
rect 151078 6536 151084 6588
rect 151136 6576 151142 6588
rect 379974 6576 379980 6588
rect 151136 6548 379980 6576
rect 151136 6536 151142 6548
rect 379974 6536 379980 6548
rect 380032 6536 380038 6588
rect 44266 6468 44272 6520
rect 44324 6508 44330 6520
rect 124582 6508 124588 6520
rect 44324 6480 124588 6508
rect 44324 6468 44330 6480
rect 124582 6468 124588 6480
rect 124640 6468 124646 6520
rect 152366 6468 152372 6520
rect 152424 6508 152430 6520
rect 396534 6508 396540 6520
rect 152424 6480 396540 6508
rect 152424 6468 152430 6480
rect 396534 6468 396540 6480
rect 396592 6468 396598 6520
rect 40678 6400 40684 6452
rect 40736 6440 40742 6452
rect 124674 6440 124680 6452
rect 40736 6412 124680 6440
rect 40736 6400 40742 6412
rect 124674 6400 124680 6412
rect 124732 6400 124738 6452
rect 169018 6400 169024 6452
rect 169076 6440 169082 6452
rect 429654 6440 429660 6452
rect 169076 6412 429660 6440
rect 169076 6400 169082 6412
rect 429654 6400 429660 6412
rect 429712 6400 429718 6452
rect 30098 6332 30104 6384
rect 30156 6372 30162 6384
rect 123110 6372 123116 6384
rect 30156 6344 123116 6372
rect 30156 6332 30162 6344
rect 123110 6332 123116 6344
rect 123168 6332 123174 6384
rect 167178 6332 167184 6384
rect 167236 6372 167242 6384
rect 436738 6372 436744 6384
rect 167236 6344 436744 6372
rect 167236 6332 167242 6344
rect 436738 6332 436744 6344
rect 436796 6332 436802 6384
rect 13538 6264 13544 6316
rect 13596 6304 13602 6316
rect 121914 6304 121920 6316
rect 13596 6276 121920 6304
rect 13596 6264 13602 6276
rect 121914 6264 121920 6276
rect 121972 6264 121978 6316
rect 161566 6264 161572 6316
rect 161624 6304 161630 6316
rect 514754 6304 514760 6316
rect 161624 6276 514760 6304
rect 161624 6264 161630 6276
rect 514754 6264 514760 6276
rect 514812 6264 514818 6316
rect 8754 6196 8760 6248
rect 8812 6236 8818 6248
rect 121730 6236 121736 6248
rect 8812 6208 121736 6236
rect 8812 6196 8818 6208
rect 121730 6196 121736 6208
rect 121788 6196 121794 6248
rect 163590 6196 163596 6248
rect 163648 6236 163654 6248
rect 540790 6236 540796 6248
rect 163648 6208 540796 6236
rect 163648 6196 163654 6208
rect 540790 6196 540796 6208
rect 540848 6196 540854 6248
rect 4062 6128 4068 6180
rect 4120 6168 4126 6180
rect 121822 6168 121828 6180
rect 4120 6140 121828 6168
rect 4120 6128 4126 6140
rect 121822 6128 121828 6140
rect 121880 6128 121886 6180
rect 163866 6128 163872 6180
rect 163924 6168 163930 6180
rect 544378 6168 544384 6180
rect 163924 6140 544384 6168
rect 163924 6128 163930 6140
rect 544378 6128 544384 6140
rect 544436 6128 544442 6180
rect 97442 5448 97448 5500
rect 97500 5488 97506 5500
rect 129642 5488 129648 5500
rect 97500 5460 129648 5488
rect 97500 5448 97506 5460
rect 129642 5448 129648 5460
rect 129700 5448 129706 5500
rect 93946 5380 93952 5432
rect 94004 5420 94010 5432
rect 128538 5420 128544 5432
rect 94004 5392 128544 5420
rect 94004 5380 94010 5392
rect 128538 5380 128544 5392
rect 128596 5380 128602 5432
rect 132586 5380 132592 5432
rect 132644 5420 132650 5432
rect 142430 5420 142436 5432
rect 132644 5392 142436 5420
rect 132644 5380 132650 5392
rect 142430 5380 142436 5392
rect 142488 5380 142494 5432
rect 85666 5312 85672 5364
rect 85724 5352 85730 5364
rect 120718 5352 120724 5364
rect 85724 5324 120724 5352
rect 85724 5312 85730 5324
rect 120718 5312 120724 5324
rect 120776 5312 120782 5364
rect 132770 5312 132776 5364
rect 132828 5352 132834 5364
rect 144730 5352 144736 5364
rect 132828 5324 144736 5352
rect 132828 5312 132834 5324
rect 144730 5312 144736 5324
rect 144788 5312 144794 5364
rect 86862 5244 86868 5296
rect 86920 5284 86926 5296
rect 127250 5284 127256 5296
rect 86920 5256 127256 5284
rect 86920 5244 86926 5256
rect 127250 5244 127256 5256
rect 127308 5244 127314 5296
rect 134518 5244 134524 5296
rect 134576 5284 134582 5296
rect 167178 5284 167184 5296
rect 134576 5256 167184 5284
rect 134576 5244 134582 5256
rect 167178 5244 167184 5256
rect 167236 5244 167242 5296
rect 76190 5176 76196 5228
rect 76248 5216 76254 5228
rect 127342 5216 127348 5228
rect 76248 5188 127348 5216
rect 76248 5176 76254 5188
rect 127342 5176 127348 5188
rect 127400 5176 127406 5228
rect 137278 5176 137284 5228
rect 137336 5216 137342 5228
rect 202690 5216 202696 5228
rect 137336 5188 202696 5216
rect 137336 5176 137342 5188
rect 202690 5176 202696 5188
rect 202748 5176 202754 5228
rect 72602 5108 72608 5160
rect 72660 5148 72666 5160
rect 127158 5148 127164 5160
rect 72660 5120 127164 5148
rect 72660 5108 72666 5120
rect 127158 5108 127164 5120
rect 127216 5108 127222 5160
rect 133046 5108 133052 5160
rect 133104 5148 133110 5160
rect 148318 5148 148324 5160
rect 133104 5120 148324 5148
rect 133104 5108 133110 5120
rect 148318 5108 148324 5120
rect 148376 5108 148382 5160
rect 149882 5108 149888 5160
rect 149940 5148 149946 5160
rect 364610 5148 364616 5160
rect 149940 5120 364616 5148
rect 149940 5108 149946 5120
rect 364610 5108 364616 5120
rect 364668 5108 364674 5160
rect 404998 5108 405004 5160
rect 405056 5148 405062 5160
rect 479334 5148 479340 5160
rect 405056 5120 479340 5148
rect 405056 5108 405062 5120
rect 479334 5108 479340 5120
rect 479392 5108 479398 5160
rect 65518 5040 65524 5092
rect 65576 5080 65582 5092
rect 125778 5080 125784 5092
rect 65576 5052 125784 5080
rect 65576 5040 65582 5052
rect 125778 5040 125784 5052
rect 125836 5040 125842 5092
rect 133138 5040 133144 5092
rect 133196 5080 133202 5092
rect 149514 5080 149520 5092
rect 133196 5052 149520 5080
rect 133196 5040 133202 5052
rect 149514 5040 149520 5052
rect 149572 5040 149578 5092
rect 160462 5040 160468 5092
rect 160520 5080 160526 5092
rect 500586 5080 500592 5092
rect 160520 5052 500592 5080
rect 160520 5040 160526 5052
rect 500586 5040 500592 5052
rect 500644 5040 500650 5092
rect 33594 4972 33600 5024
rect 33652 5012 33658 5024
rect 122926 5012 122932 5024
rect 33652 4984 122932 5012
rect 33652 4972 33658 4984
rect 122926 4972 122932 4984
rect 122984 4972 122990 5024
rect 133414 4972 133420 5024
rect 133472 5012 133478 5024
rect 153010 5012 153016 5024
rect 133472 4984 153016 5012
rect 133472 4972 133478 4984
rect 153010 4972 153016 4984
rect 153068 4972 153074 5024
rect 160554 4972 160560 5024
rect 160612 5012 160618 5024
rect 501782 5012 501788 5024
rect 160612 4984 501788 5012
rect 160612 4972 160618 4984
rect 501782 4972 501788 4984
rect 501840 4972 501846 5024
rect 28902 4904 28908 4956
rect 28960 4944 28966 4956
rect 117958 4944 117964 4956
rect 28960 4916 117964 4944
rect 28960 4904 28966 4916
rect 117958 4904 117964 4916
rect 118016 4904 118022 4956
rect 118786 4904 118792 4956
rect 118844 4944 118850 4956
rect 130838 4944 130844 4956
rect 118844 4916 130844 4944
rect 118844 4904 118850 4916
rect 130838 4904 130844 4916
rect 130896 4904 130902 4956
rect 133322 4904 133328 4956
rect 133380 4944 133386 4956
rect 151814 4944 151820 4956
rect 133380 4916 151820 4944
rect 133380 4904 133386 4916
rect 151814 4904 151820 4916
rect 151872 4904 151878 4956
rect 161934 4904 161940 4956
rect 161992 4944 161998 4956
rect 519538 4944 519544 4956
rect 161992 4916 519544 4944
rect 161992 4904 161998 4916
rect 519538 4904 519544 4916
rect 519596 4904 519602 4956
rect 5258 4836 5264 4888
rect 5316 4876 5322 4888
rect 22738 4876 22744 4888
rect 5316 4848 22744 4876
rect 5316 4836 5322 4848
rect 22738 4836 22744 4848
rect 22796 4836 22802 4888
rect 26510 4836 26516 4888
rect 26568 4876 26574 4888
rect 123018 4876 123024 4888
rect 26568 4848 123024 4876
rect 26568 4836 26574 4848
rect 123018 4836 123024 4848
rect 123076 4836 123082 4888
rect 133874 4836 133880 4888
rect 133932 4876 133938 4888
rect 158898 4876 158904 4888
rect 133932 4848 158904 4876
rect 133932 4836 133938 4848
rect 158898 4836 158904 4848
rect 158956 4836 158962 4888
rect 162210 4836 162216 4888
rect 162268 4876 162274 4888
rect 523034 4876 523040 4888
rect 162268 4848 523040 4876
rect 162268 4836 162274 4848
rect 523034 4836 523040 4848
rect 523092 4836 523098 4888
rect 21818 4768 21824 4820
rect 21876 4808 21882 4820
rect 123754 4808 123760 4820
rect 21876 4780 123760 4808
rect 21876 4768 21882 4780
rect 123754 4768 123760 4780
rect 123812 4768 123818 4820
rect 134242 4768 134248 4820
rect 134300 4808 134306 4820
rect 163682 4808 163688 4820
rect 134300 4780 163688 4808
rect 134300 4768 134306 4780
rect 163682 4768 163688 4780
rect 163740 4768 163746 4820
rect 166902 4768 166908 4820
rect 166960 4808 166966 4820
rect 577406 4808 577412 4820
rect 166960 4780 577412 4808
rect 166960 4768 166966 4780
rect 577406 4768 577412 4780
rect 577464 4768 577470 4820
rect 111610 4700 111616 4752
rect 111668 4740 111674 4752
rect 129918 4740 129924 4752
rect 111668 4712 129924 4740
rect 111668 4700 111674 4712
rect 129918 4700 129924 4712
rect 129976 4700 129982 4752
rect 117222 4632 117228 4684
rect 117280 4672 117286 4684
rect 129366 4672 129372 4684
rect 117280 4644 129372 4672
rect 117280 4632 117286 4644
rect 129366 4632 129372 4644
rect 129424 4632 129430 4684
rect 101030 4088 101036 4140
rect 101088 4128 101094 4140
rect 117222 4128 117228 4140
rect 101088 4100 117228 4128
rect 101088 4088 101094 4100
rect 117222 4088 117228 4100
rect 117280 4088 117286 4140
rect 121362 4088 121368 4140
rect 121420 4128 121426 4140
rect 143534 4128 143540 4140
rect 121420 4100 143540 4128
rect 121420 4088 121426 4100
rect 143534 4088 143540 4100
rect 143592 4088 143598 4140
rect 167546 4088 167552 4140
rect 167604 4128 167610 4140
rect 189718 4128 189724 4140
rect 167604 4100 189724 4128
rect 167604 4088 167610 4100
rect 189718 4088 189724 4100
rect 189776 4088 189782 4140
rect 276014 4088 276020 4140
rect 276072 4128 276078 4140
rect 276750 4128 276756 4140
rect 276072 4100 276756 4128
rect 276072 4088 276078 4100
rect 276750 4088 276756 4100
rect 276808 4088 276814 4140
rect 284294 4088 284300 4140
rect 284352 4128 284358 4140
rect 285030 4128 285036 4140
rect 284352 4100 285036 4128
rect 284352 4088 284358 4100
rect 285030 4088 285036 4100
rect 285088 4088 285094 4140
rect 292574 4088 292580 4140
rect 292632 4128 292638 4140
rect 293310 4128 293316 4140
rect 292632 4100 293316 4128
rect 292632 4088 292638 4100
rect 293310 4088 293316 4100
rect 293368 4088 293374 4140
rect 312538 4088 312544 4140
rect 312596 4128 312602 4140
rect 543182 4128 543188 4140
rect 312596 4100 543188 4128
rect 312596 4088 312602 4100
rect 543182 4088 543188 4100
rect 543240 4088 543246 4140
rect 83274 4020 83280 4072
rect 83332 4060 83338 4072
rect 127986 4060 127992 4072
rect 83332 4032 127992 4060
rect 83332 4020 83338 4032
rect 127986 4020 127992 4032
rect 128044 4020 128050 4072
rect 131850 4020 131856 4072
rect 131908 4060 131914 4072
rect 132954 4060 132960 4072
rect 131908 4032 132960 4060
rect 131908 4020 131914 4032
rect 132954 4020 132960 4032
rect 133012 4020 133018 4072
rect 133064 4032 135576 4060
rect 79686 3952 79692 4004
rect 79744 3992 79750 4004
rect 128078 3992 128084 4004
rect 79744 3964 128084 3992
rect 79744 3952 79750 3964
rect 128078 3952 128084 3964
rect 128136 3952 128142 4004
rect 132862 3952 132868 4004
rect 132920 3992 132926 4004
rect 133064 3992 133092 4032
rect 132920 3964 133092 3992
rect 132920 3952 132926 3964
rect 134058 3952 134064 4004
rect 134116 3992 134122 4004
rect 135548 3992 135576 4032
rect 146938 4020 146944 4072
rect 146996 4060 147002 4072
rect 160094 4060 160100 4072
rect 146996 4032 160100 4060
rect 146996 4020 147002 4032
rect 160094 4020 160100 4032
rect 160152 4020 160158 4072
rect 168098 4020 168104 4072
rect 168156 4060 168162 4072
rect 401318 4060 401324 4072
rect 168156 4032 401324 4060
rect 168156 4020 168162 4032
rect 401318 4020 401324 4032
rect 401376 4020 401382 4072
rect 145926 3992 145932 4004
rect 134116 3964 135484 3992
rect 135548 3964 145932 3992
rect 134116 3952 134122 3964
rect 69106 3884 69112 3936
rect 69164 3924 69170 3936
rect 125686 3924 125692 3936
rect 69164 3896 125692 3924
rect 69164 3884 69170 3896
rect 125686 3884 125692 3896
rect 125744 3884 125750 3936
rect 132034 3884 132040 3936
rect 132092 3924 132098 3936
rect 135254 3924 135260 3936
rect 132092 3896 135260 3924
rect 132092 3884 132098 3896
rect 135254 3884 135260 3896
rect 135312 3884 135318 3936
rect 135456 3924 135484 3964
rect 145926 3952 145932 3964
rect 145984 3952 145990 4004
rect 167362 3952 167368 4004
rect 167420 3992 167426 4004
rect 408402 3992 408408 4004
rect 167420 3964 408408 3992
rect 167420 3952 167426 3964
rect 408402 3952 408408 3964
rect 408460 3952 408466 4004
rect 161290 3924 161296 3936
rect 135456 3896 161296 3924
rect 161290 3884 161296 3896
rect 161348 3884 161354 3936
rect 167638 3884 167644 3936
rect 167696 3924 167702 3936
rect 415394 3924 415400 3936
rect 167696 3896 415400 3924
rect 167696 3884 167702 3896
rect 415394 3884 415400 3896
rect 415452 3884 415458 3936
rect 58434 3816 58440 3868
rect 58492 3856 58498 3868
rect 126606 3856 126612 3868
rect 58492 3828 126612 3856
rect 58492 3816 58498 3828
rect 126606 3816 126612 3828
rect 126664 3816 126670 3868
rect 134150 3816 134156 3868
rect 134208 3856 134214 3868
rect 162486 3856 162492 3868
rect 134208 3828 162492 3856
rect 134208 3816 134214 3828
rect 162486 3816 162492 3828
rect 162544 3816 162550 3868
rect 167270 3816 167276 3868
rect 167328 3856 167334 3868
rect 427262 3856 427268 3868
rect 167328 3828 427268 3856
rect 167328 3816 167334 3828
rect 427262 3816 427268 3828
rect 427320 3816 427326 3868
rect 51350 3748 51356 3800
rect 51408 3788 51414 3800
rect 125502 3788 125508 3800
rect 51408 3760 125508 3788
rect 51408 3748 51414 3760
rect 125502 3748 125508 3760
rect 125560 3748 125566 3800
rect 134334 3748 134340 3800
rect 134392 3788 134398 3800
rect 164878 3788 164884 3800
rect 134392 3760 164884 3788
rect 134392 3748 134398 3760
rect 164878 3748 164884 3760
rect 164936 3748 164942 3800
rect 168190 3748 168196 3800
rect 168248 3788 168254 3800
rect 445018 3788 445024 3800
rect 168248 3760 445024 3788
rect 168248 3748 168254 3760
rect 445018 3748 445024 3760
rect 445076 3748 445082 3800
rect 445110 3748 445116 3800
rect 445168 3788 445174 3800
rect 546678 3788 546684 3800
rect 445168 3760 546684 3788
rect 445168 3748 445174 3760
rect 546678 3748 546684 3760
rect 546736 3748 546742 3800
rect 47854 3680 47860 3732
rect 47912 3720 47918 3732
rect 125318 3720 125324 3732
rect 47912 3692 125324 3720
rect 47912 3680 47918 3692
rect 125318 3680 125324 3692
rect 125376 3680 125382 3732
rect 134426 3680 134432 3732
rect 134484 3720 134490 3732
rect 166074 3720 166080 3732
rect 134484 3692 166080 3720
rect 134484 3680 134490 3692
rect 166074 3680 166080 3692
rect 166132 3680 166138 3732
rect 167730 3680 167736 3732
rect 167788 3720 167794 3732
rect 462774 3720 462780 3732
rect 167788 3692 462780 3720
rect 167788 3680 167794 3692
rect 462774 3680 462780 3692
rect 462832 3680 462838 3732
rect 39574 3612 39580 3664
rect 39632 3652 39638 3664
rect 124306 3652 124312 3664
rect 39632 3624 124312 3652
rect 39632 3612 39638 3624
rect 124306 3612 124312 3624
rect 124364 3612 124370 3664
rect 134610 3612 134616 3664
rect 134668 3652 134674 3664
rect 168374 3652 168380 3664
rect 134668 3624 168380 3652
rect 134668 3612 134674 3624
rect 168374 3612 168380 3624
rect 168432 3612 168438 3664
rect 169110 3612 169116 3664
rect 169168 3652 169174 3664
rect 465166 3652 465172 3664
rect 169168 3624 465172 3652
rect 169168 3612 169174 3624
rect 465166 3612 465172 3624
rect 465224 3612 465230 3664
rect 12342 3544 12348 3596
rect 12400 3584 12406 3596
rect 122650 3584 122656 3596
rect 12400 3556 122656 3584
rect 12400 3544 12406 3556
rect 122650 3544 122656 3556
rect 122708 3544 122714 3596
rect 133046 3544 133052 3596
rect 133104 3584 133110 3596
rect 147122 3584 147128 3596
rect 133104 3556 147128 3584
rect 133104 3544 133110 3556
rect 147122 3544 147128 3556
rect 147180 3544 147186 3596
rect 159174 3544 159180 3596
rect 159232 3584 159238 3596
rect 484026 3584 484032 3596
rect 159232 3556 484032 3584
rect 159232 3544 159238 3556
rect 484026 3544 484032 3556
rect 484084 3544 484090 3596
rect 7650 3476 7656 3528
rect 7708 3516 7714 3528
rect 122558 3516 122564 3528
rect 7708 3488 122564 3516
rect 7708 3476 7714 3488
rect 122558 3476 122564 3488
rect 122616 3476 122622 3528
rect 125870 3476 125876 3528
rect 125928 3516 125934 3528
rect 131206 3516 131212 3528
rect 125928 3488 131212 3516
rect 125928 3476 125934 3488
rect 131206 3476 131212 3488
rect 131264 3476 131270 3528
rect 133230 3476 133236 3528
rect 133288 3516 133294 3528
rect 150618 3516 150624 3528
rect 133288 3488 150624 3516
rect 133288 3476 133294 3488
rect 150618 3476 150624 3488
rect 150676 3476 150682 3528
rect 159450 3476 159456 3528
rect 159508 3516 159514 3528
rect 478046 3516 478052 3528
rect 159508 3488 478052 3516
rect 159508 3476 159514 3488
rect 478046 3476 478052 3488
rect 478104 3476 478110 3528
rect 478156 3488 483014 3516
rect 2866 3408 2872 3460
rect 2924 3448 2930 3460
rect 122190 3448 122196 3460
rect 2924 3420 122196 3448
rect 2924 3408 2930 3420
rect 122190 3408 122196 3420
rect 122248 3408 122254 3460
rect 126974 3408 126980 3460
rect 127032 3448 127038 3460
rect 131574 3448 131580 3460
rect 127032 3420 131580 3448
rect 127032 3408 127038 3420
rect 131574 3408 131580 3420
rect 131632 3408 131638 3460
rect 133506 3408 133512 3460
rect 133564 3448 133570 3460
rect 154206 3448 154212 3460
rect 133564 3420 154212 3448
rect 133564 3408 133570 3420
rect 154206 3408 154212 3420
rect 154264 3408 154270 3460
rect 159726 3408 159732 3460
rect 159784 3448 159790 3460
rect 478156 3448 478184 3488
rect 159784 3420 478184 3448
rect 482986 3448 483014 3488
rect 491110 3448 491116 3460
rect 482986 3420 491116 3448
rect 159784 3408 159790 3420
rect 491110 3408 491116 3420
rect 491168 3408 491174 3460
rect 520918 3408 520924 3460
rect 520976 3448 520982 3460
rect 582190 3448 582196 3460
rect 520976 3420 582196 3448
rect 520976 3408 520982 3420
rect 582190 3408 582196 3420
rect 582248 3408 582254 3460
rect 102134 3340 102140 3392
rect 102192 3380 102198 3392
rect 103330 3380 103336 3392
rect 102192 3352 103336 3380
rect 102192 3340 102198 3352
rect 103330 3340 103336 3352
rect 103388 3340 103394 3392
rect 122282 3340 122288 3392
rect 122340 3380 122346 3392
rect 131022 3380 131028 3392
rect 122340 3352 131028 3380
rect 122340 3340 122346 3352
rect 131022 3340 131028 3352
rect 131080 3340 131086 3392
rect 131942 3340 131948 3392
rect 132000 3380 132006 3392
rect 134150 3380 134156 3392
rect 132000 3352 134156 3380
rect 132000 3340 132006 3352
rect 134150 3340 134156 3352
rect 134208 3340 134214 3392
rect 137738 3340 137744 3392
rect 137796 3380 137802 3392
rect 146938 3380 146944 3392
rect 137796 3352 146944 3380
rect 137796 3340 137802 3352
rect 146938 3340 146944 3352
rect 146996 3340 147002 3392
rect 167454 3340 167460 3392
rect 167512 3380 167518 3392
rect 394234 3380 394240 3392
rect 167512 3352 394240 3380
rect 167512 3340 167518 3352
rect 394234 3340 394240 3352
rect 394292 3340 394298 3392
rect 398926 3340 398932 3392
rect 398984 3380 398990 3392
rect 400122 3380 400128 3392
rect 398984 3352 400128 3380
rect 398984 3340 398990 3352
rect 400122 3340 400128 3352
rect 400180 3340 400186 3392
rect 415486 3340 415492 3392
rect 415544 3380 415550 3392
rect 416682 3380 416688 3392
rect 415544 3352 416688 3380
rect 415544 3340 415550 3352
rect 416682 3340 416688 3352
rect 416740 3340 416746 3392
rect 423674 3340 423680 3392
rect 423732 3380 423738 3392
rect 424962 3380 424968 3392
rect 423732 3352 424968 3380
rect 423732 3340 423738 3352
rect 424962 3340 424968 3352
rect 425020 3340 425026 3392
rect 440326 3340 440332 3392
rect 440384 3380 440390 3392
rect 441522 3380 441528 3392
rect 440384 3352 441528 3380
rect 440384 3340 440390 3352
rect 441522 3340 441528 3352
rect 441580 3340 441586 3392
rect 448606 3340 448612 3392
rect 448664 3380 448670 3392
rect 449802 3380 449808 3392
rect 448664 3352 449808 3380
rect 448664 3340 448670 3352
rect 449802 3340 449808 3352
rect 449860 3340 449866 3392
rect 456794 3340 456800 3392
rect 456852 3380 456858 3392
rect 458082 3380 458088 3392
rect 456852 3352 458088 3380
rect 456852 3340 456858 3352
rect 458082 3340 458088 3352
rect 458140 3340 458146 3392
rect 473354 3340 473360 3392
rect 473412 3380 473418 3392
rect 474182 3380 474188 3392
rect 473412 3352 474188 3380
rect 473412 3340 473418 3352
rect 474182 3340 474188 3352
rect 474240 3340 474246 3392
rect 478046 3340 478052 3392
rect 478104 3380 478110 3392
rect 487614 3380 487620 3392
rect 478104 3352 487620 3380
rect 478104 3340 478110 3352
rect 487614 3340 487620 3352
rect 487672 3340 487678 3392
rect 132126 3272 132132 3324
rect 132184 3312 132190 3324
rect 136450 3312 136456 3324
rect 132184 3284 136456 3312
rect 132184 3272 132190 3284
rect 136450 3272 136456 3284
rect 136508 3272 136514 3324
rect 150066 3272 150072 3324
rect 150124 3312 150130 3324
rect 169570 3312 169576 3324
rect 150124 3284 169576 3312
rect 150124 3272 150130 3284
rect 169570 3272 169576 3284
rect 169628 3272 169634 3324
rect 169662 3272 169668 3324
rect 169720 3312 169726 3324
rect 175458 3312 175464 3324
rect 169720 3284 175464 3312
rect 169720 3272 169726 3284
rect 175458 3272 175464 3284
rect 175516 3272 175522 3324
rect 193214 3272 193220 3324
rect 193272 3312 193278 3324
rect 194410 3312 194416 3324
rect 193272 3284 194416 3312
rect 193272 3272 193278 3284
rect 194410 3272 194416 3284
rect 194468 3272 194474 3324
rect 226334 3272 226340 3324
rect 226392 3312 226398 3324
rect 227530 3312 227536 3324
rect 226392 3284 227536 3312
rect 226392 3272 226398 3284
rect 227530 3272 227536 3284
rect 227588 3272 227594 3324
rect 299474 3272 299480 3324
rect 299532 3312 299538 3324
rect 300762 3312 300768 3324
rect 299532 3284 300768 3312
rect 299532 3272 299538 3284
rect 300762 3272 300768 3284
rect 300820 3272 300826 3324
rect 307754 3272 307760 3324
rect 307812 3312 307818 3324
rect 309042 3312 309048 3324
rect 307812 3284 309048 3312
rect 307812 3272 307818 3284
rect 309042 3272 309048 3284
rect 309100 3272 309106 3324
rect 316034 3272 316040 3324
rect 316092 3312 316098 3324
rect 317322 3312 317328 3324
rect 316092 3284 317328 3312
rect 316092 3272 316098 3284
rect 317322 3272 317328 3284
rect 317380 3272 317386 3324
rect 324406 3272 324412 3324
rect 324464 3312 324470 3324
rect 325602 3312 325608 3324
rect 324464 3284 325608 3312
rect 324464 3272 324470 3284
rect 325602 3272 325608 3284
rect 325660 3272 325666 3324
rect 332594 3272 332600 3324
rect 332652 3312 332658 3324
rect 333882 3312 333888 3324
rect 332652 3284 333888 3312
rect 332652 3272 332658 3284
rect 333882 3272 333888 3284
rect 333940 3272 333946 3324
rect 539594 3312 539600 3324
rect 335326 3284 539600 3312
rect 20622 3204 20628 3256
rect 20680 3244 20686 3256
rect 25498 3244 25504 3256
rect 20680 3216 25504 3244
rect 20680 3204 20686 3216
rect 25498 3204 25504 3216
rect 25556 3204 25562 3256
rect 165246 3204 165252 3256
rect 165304 3244 165310 3256
rect 182542 3244 182548 3256
rect 165304 3216 182548 3244
rect 165304 3204 165310 3216
rect 182542 3204 182548 3216
rect 182600 3204 182606 3256
rect 326430 3204 326436 3256
rect 326488 3244 326494 3256
rect 335326 3244 335354 3284
rect 539594 3272 539600 3284
rect 539652 3272 539658 3324
rect 326488 3216 335354 3244
rect 326488 3204 326494 3216
rect 349154 3204 349160 3256
rect 349212 3244 349218 3256
rect 350442 3244 350448 3256
rect 349212 3216 350448 3244
rect 349212 3204 349218 3216
rect 350442 3204 350448 3216
rect 350500 3204 350506 3256
rect 357434 3204 357440 3256
rect 357492 3244 357498 3256
rect 358722 3244 358728 3256
rect 357492 3216 358728 3244
rect 357492 3204 357498 3216
rect 358722 3204 358728 3216
rect 358780 3204 358786 3256
rect 365714 3204 365720 3256
rect 365772 3244 365778 3256
rect 367002 3244 367008 3256
rect 365772 3216 367008 3244
rect 365772 3204 365778 3216
rect 367002 3204 367008 3216
rect 367060 3204 367066 3256
rect 374086 3204 374092 3256
rect 374144 3244 374150 3256
rect 375282 3244 375288 3256
rect 374144 3216 375288 3244
rect 374144 3204 374150 3216
rect 375282 3204 375288 3216
rect 375340 3204 375346 3256
rect 382274 3204 382280 3256
rect 382332 3244 382338 3256
rect 383562 3244 383568 3256
rect 382332 3216 383568 3244
rect 382332 3204 382338 3216
rect 383562 3204 383568 3216
rect 383620 3204 383626 3256
rect 390554 3204 390560 3256
rect 390612 3244 390618 3256
rect 391842 3244 391848 3256
rect 390612 3216 391848 3244
rect 390612 3204 390618 3216
rect 391842 3204 391848 3216
rect 391900 3204 391906 3256
rect 128170 3068 128176 3120
rect 128228 3108 128234 3120
rect 131390 3108 131396 3120
rect 128228 3080 131396 3108
rect 128228 3068 128234 3080
rect 131390 3068 131396 3080
rect 131448 3068 131454 3120
rect 129366 3000 129372 3052
rect 129424 3040 129430 3052
rect 131482 3040 131488 3052
rect 129424 3012 131488 3040
rect 129424 3000 129430 3012
rect 131482 3000 131488 3012
rect 131540 3000 131546 3052
rect 136174 2932 136180 2984
rect 136232 2972 136238 2984
rect 141234 2972 141240 2984
rect 136232 2944 141240 2972
rect 136232 2932 136238 2944
rect 141234 2932 141240 2944
rect 141292 2932 141298 2984
rect 432046 1776 432052 1828
rect 432104 1816 432110 1828
rect 433242 1816 433248 1828
rect 432104 1788 433248 1816
rect 432104 1776 432110 1788
rect 433242 1776 433248 1788
rect 433300 1776 433306 1828
<< via1 >>
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 201500 702992 201552 703044
rect 202788 702992 202840 703044
rect 413284 700408 413336 700460
rect 429844 700408 429896 700460
rect 410524 700340 410576 700392
rect 494796 700340 494848 700392
rect 409144 700272 409196 700324
rect 559656 700272 559708 700324
rect 348792 699796 348844 699848
rect 351184 699796 351236 699848
rect 153016 699660 153068 699712
rect 154120 699660 154172 699712
rect 215208 699592 215260 699644
rect 218980 699660 219032 699712
rect 262864 699592 262916 699644
rect 267648 699660 267700 699712
rect 282184 699660 282236 699712
rect 283840 699660 283892 699712
rect 332508 699660 332560 699712
rect 336004 699660 336056 699712
rect 364984 698096 365036 698148
rect 369124 698096 369176 698148
rect 146944 696872 146996 696924
rect 153016 696940 153068 696992
rect 211804 693608 211856 693660
rect 215208 693608 215260 693660
rect 226984 693404 227036 693456
rect 234620 693404 234672 693456
rect 351184 690616 351236 690668
rect 359464 690616 359516 690668
rect 369124 690344 369176 690396
rect 371240 690344 371292 690396
rect 145656 688644 145708 688696
rect 146944 688644 146996 688696
rect 191104 687896 191156 687948
rect 201500 687896 201552 687948
rect 371240 687896 371292 687948
rect 377404 687896 377456 687948
rect 336004 684428 336056 684480
rect 341248 684428 341300 684480
rect 144184 683952 144236 684004
rect 145656 683952 145708 684004
rect 299480 681164 299532 681216
rect 305000 681164 305052 681216
rect 187976 680552 188028 680604
rect 191104 680552 191156 680604
rect 359464 679260 359516 679312
rect 362224 679260 362276 679312
rect 341248 679124 341300 679176
rect 344284 679124 344336 679176
rect 280896 678988 280948 679040
rect 282184 678988 282236 679040
rect 377404 678920 377456 678972
rect 385684 678920 385736 678972
rect 185584 677560 185636 677612
rect 187976 677560 188028 677612
rect 279424 677016 279476 677068
rect 280896 677016 280948 677068
rect 221464 676744 221516 676796
rect 226984 676744 227036 676796
rect 305000 675588 305052 675640
rect 307760 675588 307812 675640
rect 259460 674976 259512 675028
rect 262864 674976 262916 675028
rect 307760 672732 307812 672784
rect 319904 672732 319956 672784
rect 215300 672052 215352 672104
rect 221464 672052 221516 672104
rect 255688 671984 255740 672036
rect 259460 672052 259512 672104
rect 3516 670692 3568 670744
rect 15844 670692 15896 670744
rect 140320 670624 140372 670676
rect 144184 670692 144236 670744
rect 407764 670692 407816 670744
rect 580172 670692 580224 670744
rect 362224 669944 362276 669996
rect 383936 669944 383988 669996
rect 253204 669332 253256 669384
rect 255688 669332 255740 669384
rect 344284 669264 344336 669316
rect 346676 669264 346728 669316
rect 138664 667904 138716 667956
rect 140320 667904 140372 667956
rect 204904 667156 204956 667208
rect 215300 667156 215352 667208
rect 383936 665796 383988 665848
rect 395344 665796 395396 665848
rect 210424 665116 210476 665168
rect 211804 665116 211856 665168
rect 319904 665116 319956 665168
rect 324964 665116 325016 665168
rect 385684 665116 385736 665168
rect 389824 665116 389876 665168
rect 197268 664436 197320 664488
rect 204904 664436 204956 664488
rect 346676 664436 346728 664488
rect 364984 664436 365036 664488
rect 277492 662396 277544 662448
rect 279424 662396 279476 662448
rect 191104 661036 191156 661088
rect 197268 661036 197320 661088
rect 276664 660560 276716 660612
rect 277492 660560 277544 660612
rect 389824 656820 389876 656872
rect 392584 656820 392636 656872
rect 136732 651380 136784 651432
rect 138664 651380 138716 651432
rect 178040 650632 178092 650684
rect 191104 650632 191156 650684
rect 170404 647844 170456 647896
rect 178040 647844 178092 647896
rect 133696 646824 133748 646876
rect 136732 646824 136784 646876
rect 392584 646144 392636 646196
rect 395528 646144 395580 646196
rect 131764 644444 131816 644496
rect 133696 644444 133748 644496
rect 181444 640296 181496 640348
rect 185584 640296 185636 640348
rect 272524 640228 272576 640280
rect 276664 640296 276716 640348
rect 207664 636216 207716 636268
rect 210424 636216 210476 636268
rect 324964 635468 325016 635520
rect 329196 635468 329248 635520
rect 155224 632680 155276 632732
rect 170404 632680 170456 632732
rect 128360 632068 128412 632120
rect 131764 632068 131816 632120
rect 127624 629688 127676 629740
rect 128360 629688 128412 629740
rect 329196 629212 329248 629264
rect 331864 629212 331916 629264
rect 364984 626492 365036 626544
rect 369124 626492 369176 626544
rect 204904 625200 204956 625252
rect 207664 625200 207716 625252
rect 124220 623704 124272 623756
rect 127624 623772 127676 623824
rect 175924 622684 175976 622736
rect 181444 622684 181496 622736
rect 123484 620984 123536 621036
rect 124220 620984 124272 621036
rect 3516 618264 3568 618316
rect 37924 618264 37976 618316
rect 406384 616836 406436 616888
rect 579988 616836 580040 616888
rect 169024 616088 169076 616140
rect 175924 616088 175976 616140
rect 270500 614116 270552 614168
rect 272524 614116 272576 614168
rect 331864 611260 331916 611312
rect 337384 611260 337436 611312
rect 203524 609220 203576 609272
rect 204904 609220 204956 609272
rect 263600 609220 263652 609272
rect 270500 609220 270552 609272
rect 262864 606568 262916 606620
rect 263600 606568 263652 606620
rect 251916 601672 251968 601724
rect 253204 601672 253256 601724
rect 120724 600244 120776 600296
rect 123484 600312 123536 600364
rect 261484 598612 261536 598664
rect 262864 598612 262916 598664
rect 250444 596912 250496 596964
rect 251916 596912 251968 596964
rect 337384 592220 337436 592272
rect 339500 592220 339552 592272
rect 112444 591268 112496 591320
rect 120724 591268 120776 591320
rect 339500 590588 339552 590640
rect 343640 590588 343692 590640
rect 343640 587596 343692 587648
rect 347044 587596 347096 587648
rect 246304 586440 246356 586492
rect 250444 586508 250496 586560
rect 369124 582224 369176 582276
rect 373264 582224 373316 582276
rect 144184 571956 144236 572008
rect 155224 571956 155276 572008
rect 3332 565836 3384 565888
rect 19984 565836 20036 565888
rect 111064 565836 111116 565888
rect 112444 565836 112496 565888
rect 243544 564408 243596 564460
rect 246304 564408 246356 564460
rect 140780 563048 140832 563100
rect 144184 563048 144236 563100
rect 260104 563048 260156 563100
rect 261484 563048 261536 563100
rect 405004 563048 405056 563100
rect 580172 563048 580224 563100
rect 373264 562980 373316 563032
rect 376668 562980 376720 563032
rect 347044 562300 347096 562352
rect 349804 562300 349856 562352
rect 127624 560940 127676 560992
rect 140780 560940 140832 560992
rect 376668 559512 376720 559564
rect 383660 559512 383712 559564
rect 202144 558832 202196 558884
rect 203524 558832 203576 558884
rect 383660 556724 383712 556776
rect 389824 556724 389876 556776
rect 349804 555432 349856 555484
rect 368388 555432 368440 555484
rect 117228 554004 117280 554056
rect 127624 554004 127676 554056
rect 2780 553800 2832 553852
rect 4804 553800 4856 553852
rect 109684 551284 109736 551336
rect 111064 551284 111116 551336
rect 104992 549856 105044 549908
rect 117228 549856 117280 549908
rect 368388 549856 368440 549908
rect 382924 549856 382976 549908
rect 94504 542988 94556 543040
rect 104992 542988 105044 543040
rect 389824 537956 389876 538008
rect 395160 537956 395212 538008
rect 83464 537548 83516 537600
rect 94504 537548 94556 537600
rect 62672 537480 62724 537532
rect 169760 537480 169812 537532
rect 395160 534080 395212 534132
rect 397552 534080 397604 534132
rect 61384 532992 61436 533044
rect 62672 532992 62724 533044
rect 257068 528572 257120 528624
rect 260104 528572 260156 528624
rect 382924 528028 382976 528080
rect 386328 528028 386380 528080
rect 386328 522928 386380 522980
rect 391204 522928 391256 522980
rect 255964 522112 256016 522164
rect 257068 522112 257120 522164
rect 239404 520208 239456 520260
rect 243544 520276 243596 520328
rect 105544 516060 105596 516112
rect 109684 516128 109736 516180
rect 3332 514768 3384 514820
rect 42064 514768 42116 514820
rect 80060 512932 80112 512984
rect 83464 512932 83516 512984
rect 253204 511912 253256 511964
rect 255964 511912 256016 511964
rect 403624 510620 403676 510672
rect 579804 510620 579856 510672
rect 69480 509872 69532 509924
rect 80060 509872 80112 509924
rect 117964 508512 118016 508564
rect 136640 508512 136692 508564
rect 61476 504364 61528 504416
rect 69480 504364 69532 504416
rect 200764 502936 200816 502988
rect 202144 502936 202196 502988
rect 2780 501032 2832 501084
rect 4896 501032 4948 501084
rect 158720 498788 158772 498840
rect 169024 498788 169076 498840
rect 391204 498380 391256 498432
rect 393964 498380 394016 498432
rect 250444 493960 250496 494012
rect 253204 494028 253256 494080
rect 150440 490560 150492 490612
rect 158720 490560 158772 490612
rect 116584 487160 116636 487212
rect 117964 487160 118016 487212
rect 146024 487160 146076 487212
rect 150440 487160 150492 487212
rect 237380 486480 237432 486532
rect 239404 486480 239456 486532
rect 142804 484304 142856 484356
rect 146024 484304 146076 484356
rect 236644 482536 236696 482588
rect 237380 482536 237432 482588
rect 135168 479476 135220 479528
rect 142804 479476 142856 479528
rect 249432 478864 249484 478916
rect 250444 478864 250496 478916
rect 129740 476280 129792 476332
rect 135168 476280 135220 476332
rect 393964 475396 394016 475448
rect 395436 475396 395488 475448
rect 58624 474648 58676 474700
rect 61476 474648 61528 474700
rect 247684 474376 247736 474428
rect 249432 474376 249484 474428
rect 115204 472948 115256 473000
rect 116584 472948 116636 473000
rect 199384 471996 199436 472048
rect 200764 471996 200816 472048
rect 120724 471248 120776 471300
rect 129740 471248 129792 471300
rect 198004 469208 198056 469260
rect 199384 469208 199436 469260
rect 55864 466420 55916 466472
rect 58624 466420 58676 466472
rect 2780 462544 2832 462596
rect 5080 462544 5132 462596
rect 193864 456696 193916 456748
rect 198004 456764 198056 456816
rect 400864 456764 400916 456816
rect 579988 456764 580040 456816
rect 46204 451868 46256 451920
rect 55864 451868 55916 451920
rect 117964 449896 118016 449948
rect 120724 449896 120776 449948
rect 2780 448808 2832 448860
rect 4988 448808 5040 448860
rect 399576 444388 399628 444440
rect 580080 444388 580132 444440
rect 45100 428272 45152 428324
rect 46204 428272 46256 428324
rect 111064 427048 111116 427100
rect 117964 427048 118016 427100
rect 192484 425688 192536 425740
rect 193864 425688 193916 425740
rect 244924 419432 244976 419484
rect 247684 419500 247736 419552
rect 398104 418140 398156 418192
rect 580080 418140 580132 418192
rect 102784 412632 102836 412684
rect 105544 412632 105596 412684
rect 3332 409912 3384 409964
rect 8944 409912 8996 409964
rect 399484 404336 399536 404388
rect 580080 404336 580132 404388
rect 243544 404268 243596 404320
rect 244924 404268 244976 404320
rect 2780 397468 2832 397520
rect 5172 397468 5224 397520
rect 235264 394612 235316 394664
rect 236644 394612 236696 394664
rect 101404 391960 101456 392012
rect 102784 391960 102836 392012
rect 189724 391960 189776 392012
rect 192484 391960 192536 392012
rect 108304 390532 108356 390584
rect 111064 390532 111116 390584
rect 396724 378156 396776 378208
rect 580080 378156 580132 378208
rect 58624 376592 58676 376644
rect 61384 376592 61436 376644
rect 239404 371220 239456 371272
rect 243544 371220 243596 371272
rect 188436 369860 188488 369912
rect 189724 369860 189776 369912
rect 98644 368432 98696 368484
rect 101404 368500 101456 368552
rect 186964 365508 187016 365560
rect 188436 365508 188488 365560
rect 396908 364352 396960 364404
rect 579804 364352 579856 364404
rect 232504 360204 232556 360256
rect 235264 360204 235316 360256
rect 3332 357416 3384 357468
rect 10324 357416 10376 357468
rect 69664 356668 69716 356720
rect 115204 356668 115256 356720
rect 99012 353948 99064 354000
rect 108304 353948 108356 354000
rect 185584 353268 185636 353320
rect 186964 353268 187016 353320
rect 235264 352044 235316 352096
rect 239404 352044 239456 352096
rect 418804 351908 418856 351960
rect 580080 351908 580132 351960
rect 94504 348848 94556 348900
rect 99012 348848 99064 348900
rect 229744 348780 229796 348832
rect 232504 348780 232556 348832
rect 56876 346332 56928 346384
rect 58624 346332 58676 346384
rect 2780 345176 2832 345228
rect 5264 345176 5316 345228
rect 233976 342252 234028 342304
rect 235264 342252 235316 342304
rect 232504 340008 232556 340060
rect 233976 340008 234028 340060
rect 68284 339668 68336 339720
rect 69664 339668 69716 339720
rect 97264 338784 97316 338836
rect 98644 338784 98696 338836
rect 55864 338240 55916 338292
rect 56876 338240 56928 338292
rect 87604 336744 87656 336796
rect 94504 336744 94556 336796
rect 225328 335248 225380 335300
rect 229744 335316 229796 335368
rect 231216 333956 231268 334008
rect 232504 333956 232556 334008
rect 95884 329060 95936 329112
rect 97264 329060 97316 329112
rect 224224 328992 224276 329044
rect 225328 328992 225380 329044
rect 229836 326272 229888 326324
rect 231216 326272 231268 326324
rect 396816 324300 396868 324352
rect 580080 324300 580132 324352
rect 81716 323552 81768 323604
rect 87604 323552 87656 323604
rect 227720 323552 227772 323604
rect 229836 323552 229888 323604
rect 53104 323348 53156 323400
rect 55864 323348 55916 323400
rect 221464 322940 221516 322992
rect 224224 322940 224276 322992
rect 94780 321716 94832 321768
rect 95884 321716 95936 321768
rect 182456 320764 182508 320816
rect 185584 320764 185636 320816
rect 91100 319744 91152 319796
rect 94780 319744 94832 319796
rect 85580 318724 85632 318776
rect 88340 318724 88392 318776
rect 180800 318656 180852 318708
rect 182456 318656 182508 318708
rect 223120 318248 223172 318300
rect 227720 318248 227772 318300
rect 88340 317364 88392 317416
rect 91100 317432 91152 317484
rect 79232 316752 79284 316804
rect 81716 316752 81768 316804
rect 62764 313896 62816 313948
rect 104900 313896 104952 313948
rect 178684 313624 178736 313676
rect 180800 313624 180852 313676
rect 79324 313352 79376 313404
rect 85580 313352 85632 313404
rect 220084 313284 220136 313336
rect 221464 313284 221516 313336
rect 220176 311856 220228 311908
rect 223120 311856 223172 311908
rect 397092 311856 397144 311908
rect 580080 311856 580132 311908
rect 69664 311108 69716 311160
rect 79232 311108 79284 311160
rect 85396 309408 85448 309460
rect 88248 309408 88300 309460
rect 81348 307776 81400 307828
rect 85396 307776 85448 307828
rect 3240 304988 3292 305040
rect 24124 304988 24176 305040
rect 51724 304988 51776 305040
rect 53104 304988 53156 305040
rect 67180 303628 67232 303680
rect 69664 303628 69716 303680
rect 57244 301452 57296 301504
rect 79324 301452 79376 301504
rect 61384 301044 61436 301096
rect 62764 301044 62816 301096
rect 79324 300296 79376 300348
rect 81348 300296 81400 300348
rect 66904 300160 66956 300212
rect 68284 300160 68336 300212
rect 51816 300092 51868 300144
rect 67180 300092 67232 300144
rect 417424 298120 417476 298172
rect 580080 298120 580132 298172
rect 3240 292544 3292 292596
rect 43444 292544 43496 292596
rect 76564 292544 76616 292596
rect 79324 292544 79376 292596
rect 218060 292544 218112 292596
rect 220176 292544 220228 292596
rect 215944 289824 215996 289876
rect 218060 289824 218112 289876
rect 55864 288328 55916 288380
rect 57244 288328 57296 288380
rect 49608 287580 49660 287632
rect 51816 287580 51868 287632
rect 46204 284316 46256 284368
rect 49608 284316 49660 284368
rect 72056 281936 72108 281988
rect 76564 281936 76616 281988
rect 60004 280780 60056 280832
rect 61384 280780 61436 280832
rect 213920 279964 213972 280016
rect 215944 279964 215996 280016
rect 69480 279692 69532 279744
rect 72056 279692 72108 279744
rect 175924 276020 175976 276072
rect 178684 276020 178736 276072
rect 218060 276020 218112 276072
rect 220084 276020 220136 276072
rect 204168 275272 204220 275324
rect 213920 275272 213972 275324
rect 45008 274728 45060 274780
rect 46204 274728 46256 274780
rect 57980 274660 58032 274712
rect 60004 274660 60056 274712
rect 54484 272892 54536 272944
rect 55864 272892 55916 272944
rect 202144 271872 202196 271924
rect 204168 271872 204220 271924
rect 397000 271872 397052 271924
rect 579804 271872 579856 271924
rect 65524 270444 65576 270496
rect 69480 270512 69532 270564
rect 213368 270444 213420 270496
rect 217968 270512 218020 270564
rect 52368 269084 52420 269136
rect 57888 269084 57940 269136
rect 63500 266500 63552 266552
rect 66904 266500 66956 266552
rect 51080 266364 51132 266416
rect 54484 266364 54536 266416
rect 197728 266296 197780 266348
rect 202144 266364 202196 266416
rect 208400 264188 208452 264240
rect 213368 264188 213420 264240
rect 50344 262828 50396 262880
rect 63500 262828 63552 262880
rect 195244 261808 195296 261860
rect 197728 261808 197780 261860
rect 189080 261468 189132 261520
rect 208308 261468 208360 261520
rect 50896 261196 50948 261248
rect 52368 261196 52420 261248
rect 174268 260788 174320 260840
rect 175924 260788 175976 260840
rect 47584 260448 47636 260500
rect 51080 260448 51132 260500
rect 60648 259360 60700 259412
rect 65524 259428 65576 259480
rect 185584 259360 185636 259412
rect 189080 259428 189132 259480
rect 49240 258952 49292 259004
rect 50896 258952 50948 259004
rect 397184 258068 397236 258120
rect 579988 258068 580040 258120
rect 47492 256708 47544 256760
rect 49240 256708 49292 256760
rect 193864 256708 193916 256760
rect 195244 256708 195296 256760
rect 3148 253920 3200 253972
rect 22744 253920 22796 253972
rect 45836 253920 45888 253972
rect 47492 253920 47544 253972
rect 48688 252560 48740 252612
rect 50344 252560 50396 252612
rect 173164 252492 173216 252544
rect 174268 252492 174320 252544
rect 57980 251880 58032 251932
rect 60648 251880 60700 251932
rect 47676 251812 47728 251864
rect 71780 251812 71832 251864
rect 46940 249432 46992 249484
rect 48688 249432 48740 249484
rect 52460 249024 52512 249076
rect 57980 249024 58032 249076
rect 49700 247052 49752 247104
rect 51724 247052 51776 247104
rect 166264 246984 166316 247036
rect 173164 247052 173216 247104
rect 182916 246984 182968 247036
rect 185584 247052 185636 247104
rect 414664 244264 414716 244316
rect 579988 244264 580040 244316
rect 44824 243856 44876 243908
rect 46848 243856 46900 243908
rect 45744 243516 45796 243568
rect 49700 243516 49752 243568
rect 47124 241680 47176 241732
rect 52368 241680 52420 241732
rect 45652 241408 45704 241460
rect 47676 241408 47728 241460
rect 45560 241340 45612 241392
rect 47584 241340 47636 241392
rect 45376 240864 45428 240916
rect 166264 240864 166316 240916
rect 45284 240796 45336 240848
rect 182916 240796 182968 240848
rect 44916 240728 44968 240780
rect 193864 240728 193916 240780
rect 3056 240116 3108 240168
rect 43536 240116 43588 240168
rect 47124 240116 47176 240168
rect 45468 240048 45520 240100
rect 395436 240048 395488 240100
rect 396540 240048 396592 240100
rect 396540 238824 396592 238876
rect 45192 238756 45244 238808
rect 45836 238756 45888 238808
rect 396540 238688 396592 238740
rect 44824 233180 44876 233232
rect 45836 233180 45888 233232
rect 45192 232908 45244 232960
rect 45468 232364 45520 232416
rect 86316 232364 86368 232416
rect 45376 232296 45428 232348
rect 46848 232296 46900 232348
rect 46940 232296 46992 232348
rect 45284 232228 45336 232280
rect 46204 232228 46256 232280
rect 45744 232160 45796 232212
rect 53196 232160 53248 232212
rect 394700 232092 394752 232144
rect 396540 232092 396592 232144
rect 44916 231140 44968 231192
rect 52368 231140 52420 231192
rect 86316 231140 86368 231192
rect 153200 231140 153252 231192
rect 4068 231072 4120 231124
rect 177856 231072 177908 231124
rect 46204 230392 46256 230444
rect 48964 230392 49016 230444
rect 387800 230392 387852 230444
rect 394700 230460 394752 230512
rect 45836 230324 45888 230376
rect 47584 230324 47636 230376
rect 46940 230256 46992 230308
rect 52460 230256 52512 230308
rect 166264 229712 166316 229764
rect 176660 229712 176712 229764
rect 391940 229100 391992 229152
rect 394608 229100 394660 229152
rect 157984 228420 158036 228472
rect 266544 228420 266596 228472
rect 297364 228420 297416 228472
rect 327080 228420 327132 228472
rect 117228 228352 117280 228404
rect 138664 228352 138716 228404
rect 153200 228352 153252 228404
rect 165068 228352 165120 228404
rect 236644 228352 236696 228404
rect 386512 228352 386564 228404
rect 46940 228284 46992 228336
rect 52552 228284 52604 228336
rect 52368 228080 52420 228132
rect 53840 228080 53892 228132
rect 53196 227536 53248 227588
rect 57244 227536 57296 227588
rect 165068 227196 165120 227248
rect 170404 227196 170456 227248
rect 52552 226992 52604 227044
rect 59268 226992 59320 227044
rect 53840 226312 53892 226364
rect 56968 226244 57020 226296
rect 387800 224884 387852 224936
rect 391848 224952 391900 225004
rect 384948 223660 385000 223712
rect 387708 223660 387760 223712
rect 59268 223592 59320 223644
rect 52460 223524 52512 223576
rect 55772 223524 55824 223576
rect 66996 223524 67048 223576
rect 387064 223524 387116 223576
rect 390376 223524 390428 223576
rect 56968 222844 57020 222896
rect 58624 222844 58676 222896
rect 45008 220804 45060 220856
rect 47676 220804 47728 220856
rect 48964 220804 49016 220856
rect 53932 220736 53984 220788
rect 55772 220736 55824 220788
rect 62764 220736 62816 220788
rect 66996 220736 67048 220788
rect 69664 220736 69716 220788
rect 385040 220464 385092 220516
rect 387708 220464 387760 220516
rect 381360 219444 381412 219496
rect 384948 219444 385000 219496
rect 384304 218084 384356 218136
rect 387064 218084 387116 218136
rect 115848 218016 115900 218068
rect 579804 218016 579856 218068
rect 47584 217404 47636 217456
rect 53840 217404 53892 217456
rect 58624 216656 58676 216708
rect 65524 216588 65576 216640
rect 53932 215908 53984 215960
rect 63408 215908 63460 215960
rect 53840 215296 53892 215348
rect 56692 215228 56744 215280
rect 3148 213936 3200 213988
rect 175372 213936 175424 213988
rect 380900 213868 380952 213920
rect 385040 213936 385092 213988
rect 378784 213596 378836 213648
rect 381360 213596 381412 213648
rect 57244 213188 57296 213240
rect 71044 213188 71096 213240
rect 378140 211624 378192 211676
rect 380900 211624 380952 211676
rect 56692 211148 56744 211200
rect 47676 211080 47728 211132
rect 51356 211080 51408 211132
rect 62120 211080 62172 211132
rect 63500 210196 63552 210248
rect 65616 210196 65668 210248
rect 393320 209924 393372 209976
rect 397552 209924 397604 209976
rect 45100 208360 45152 208412
rect 46388 208360 46440 208412
rect 69664 208360 69716 208412
rect 72424 208292 72476 208344
rect 62120 207612 62172 207664
rect 63500 207612 63552 207664
rect 65524 207000 65576 207052
rect 69664 206932 69716 206984
rect 382924 206252 382976 206304
rect 393320 206252 393372 206304
rect 62764 205640 62816 205692
rect 188344 205640 188396 205692
rect 579988 205640 580040 205692
rect 65524 205572 65576 205624
rect 65616 205436 65668 205488
rect 66904 205436 66956 205488
rect 51356 204892 51408 204944
rect 58624 204892 58676 204944
rect 375748 204620 375800 204672
rect 378048 204620 378100 204672
rect 71044 203532 71096 203584
rect 95148 203532 95200 203584
rect 366364 203532 366416 203584
rect 375748 203532 375800 203584
rect 377128 202988 377180 203040
rect 378784 202988 378836 203040
rect 63500 202172 63552 202224
rect 66260 202172 66312 202224
rect 3148 201492 3200 201544
rect 22836 201492 22888 201544
rect 46388 201424 46440 201476
rect 47584 201424 47636 201476
rect 95148 200744 95200 200796
rect 104900 200744 104952 200796
rect 375380 200744 375432 200796
rect 377128 200744 377180 200796
rect 155960 199384 156012 199436
rect 296720 199384 296772 199436
rect 72424 199180 72476 199232
rect 75276 199180 75328 199232
rect 66260 198704 66312 198756
rect 68192 198704 68244 198756
rect 170404 198704 170456 198756
rect 171784 198704 171836 198756
rect 104900 198500 104952 198552
rect 108304 198500 108356 198552
rect 65524 198092 65576 198144
rect 66260 198092 66312 198144
rect 148968 197956 149020 198008
rect 207020 197956 207072 198008
rect 154488 197412 154540 197464
rect 155960 197412 156012 197464
rect 364984 197344 365036 197396
rect 366364 197344 366416 197396
rect 379520 197344 379572 197396
rect 382924 197344 382976 197396
rect 152740 197276 152792 197328
rect 157984 197276 158036 197328
rect 147956 196732 148008 196784
rect 166264 196732 166316 196784
rect 160836 196664 160888 196716
rect 236644 196664 236696 196716
rect 151176 196596 151228 196648
rect 236000 196596 236052 196648
rect 66904 196460 66956 196512
rect 68284 196460 68336 196512
rect 58624 196256 58676 196308
rect 61384 196256 61436 196308
rect 68192 195984 68244 196036
rect 71044 195916 71096 195968
rect 138664 195916 138716 195968
rect 141424 195916 141476 195968
rect 157524 195916 157576 195968
rect 356060 195916 356112 195968
rect 86960 195848 87012 195900
rect 139400 195848 139452 195900
rect 157432 195848 157484 195900
rect 297364 195848 297416 195900
rect 56600 195780 56652 195832
rect 138112 195780 138164 195832
rect 66260 195440 66312 195492
rect 68376 195440 68428 195492
rect 75276 195440 75328 195492
rect 77944 195440 77996 195492
rect 376024 195168 376076 195220
rect 379520 195168 379572 195220
rect 371240 194352 371292 194404
rect 375288 194352 375340 194404
rect 217324 193808 217376 193860
rect 580172 193808 580224 193860
rect 47584 193128 47636 193180
rect 48964 193128 49016 193180
rect 365076 191768 365128 191820
rect 371240 191836 371292 191888
rect 157340 189864 157392 189916
rect 61384 188300 61436 188352
rect 68928 188300 68980 188352
rect 71044 187892 71096 187944
rect 73160 187892 73212 187944
rect 3148 187688 3200 187740
rect 112444 187688 112496 187740
rect 166172 187620 166224 187672
rect 399576 187620 399628 187672
rect 108304 186600 108356 186652
rect 111064 186600 111116 186652
rect 45652 184832 45704 184884
rect 53104 184832 53156 184884
rect 73160 184832 73212 184884
rect 75184 184832 75236 184884
rect 135260 184152 135312 184204
rect 142436 184220 142488 184272
rect 376116 182792 376168 182844
rect 384304 182792 384356 182844
rect 68928 181432 68980 181484
rect 83464 181432 83516 181484
rect 117320 180140 117372 180192
rect 136364 180140 136416 180192
rect 53104 180072 53156 180124
rect 63500 180072 63552 180124
rect 122104 180072 122156 180124
rect 141240 180344 141292 180396
rect 77944 179392 77996 179444
rect 79324 179392 79376 179444
rect 136364 178780 136416 178832
rect 136732 178780 136784 178832
rect 120724 178644 120776 178696
rect 136456 178644 136508 178696
rect 154396 178168 154448 178220
rect 157800 178168 157852 178220
rect 75184 178100 75236 178152
rect 77208 178100 77260 178152
rect 135996 178100 136048 178152
rect 136548 178100 136600 178152
rect 48964 178032 49016 178084
rect 49700 178032 49752 178084
rect 115756 178032 115808 178084
rect 153936 178032 153988 178084
rect 158628 178032 158680 178084
rect 579988 178032 580040 178084
rect 63500 177284 63552 177336
rect 69756 177284 69808 177336
rect 120080 177284 120132 177336
rect 135996 177284 136048 177336
rect 135720 176128 135772 176180
rect 136548 176128 136600 176180
rect 122840 176060 122892 176112
rect 136456 176060 136508 176112
rect 121460 175924 121512 175976
rect 136364 175924 136416 175976
rect 149980 175516 150032 175568
rect 144460 175448 144512 175500
rect 144092 175380 144144 175432
rect 153936 175380 153988 175432
rect 77208 175244 77260 175296
rect 154396 175244 154448 175296
rect 156512 175244 156564 175296
rect 78680 175176 78732 175228
rect 141700 174700 141752 174752
rect 141792 174700 141844 174752
rect 125600 174496 125652 174548
rect 135720 174496 135772 174548
rect 153476 174564 153528 174616
rect 162492 174496 162544 174548
rect 115664 174292 115716 174344
rect 580448 174292 580500 174344
rect 129740 173884 129792 173936
rect 137284 173884 137336 173936
rect 153476 173884 153528 173936
rect 83464 173136 83516 173188
rect 91560 173136 91612 173188
rect 126980 173136 127032 173188
rect 136640 173136 136692 173188
rect 161480 173136 161532 173188
rect 166540 173136 166592 173188
rect 159456 173000 159508 173052
rect 143448 172932 143500 172984
rect 145656 172932 145708 172984
rect 146484 172932 146536 172984
rect 148600 172932 148652 172984
rect 156512 172932 156564 172984
rect 158444 172932 158496 172984
rect 143540 172864 143592 172916
rect 146668 172864 146720 172916
rect 142436 172796 142488 172848
rect 147588 172796 147640 172848
rect 49700 172456 49752 172508
rect 53104 172456 53156 172508
rect 78680 172456 78732 172508
rect 80612 172456 80664 172508
rect 133880 172116 133932 172168
rect 140780 172116 140832 172168
rect 131120 171912 131172 171964
rect 138664 171912 138716 171964
rect 140780 171776 140832 171828
rect 144920 171776 144972 171828
rect 132500 171504 132552 171556
rect 139676 171504 139728 171556
rect 128360 171096 128412 171148
rect 136732 171096 136784 171148
rect 111064 170688 111116 170740
rect 114468 170688 114520 170740
rect 45560 170348 45612 170400
rect 63500 170348 63552 170400
rect 91560 170348 91612 170400
rect 99380 170348 99432 170400
rect 358544 170348 358596 170400
rect 376116 170348 376168 170400
rect 117412 169736 117464 169788
rect 122104 169736 122156 169788
rect 362960 169056 363012 169108
rect 364984 169056 365036 169108
rect 366364 168988 366416 169040
rect 376024 168988 376076 169040
rect 79324 168716 79376 168768
rect 81532 168716 81584 168768
rect 80612 168444 80664 168496
rect 83464 168444 83516 168496
rect 114468 167628 114520 167680
rect 138664 167628 138716 167680
rect 355324 167016 355376 167068
rect 358544 167016 358596 167068
rect 68376 166404 68428 166456
rect 69848 166404 69900 166456
rect 115112 166268 115164 166320
rect 117412 166268 117464 166320
rect 185584 165588 185636 165640
rect 579804 165588 579856 165640
rect 363604 165112 363656 165164
rect 365076 165112 365128 165164
rect 81532 164160 81584 164212
rect 83556 164160 83608 164212
rect 63500 163548 63552 163600
rect 66260 163548 66312 163600
rect 99380 163480 99432 163532
rect 113732 163480 113784 163532
rect 53104 162936 53156 162988
rect 55864 162936 55916 162988
rect 3148 162868 3200 162920
rect 175280 162868 175332 162920
rect 358452 162800 358504 162852
rect 362960 162868 363012 162920
rect 66260 160692 66312 160744
rect 79324 160692 79376 160744
rect 138664 160692 138716 160744
rect 147680 160692 147732 160744
rect 69664 159196 69716 159248
rect 71688 159196 71740 159248
rect 356060 157360 356112 157412
rect 358452 157360 358504 157412
rect 79324 157292 79376 157344
rect 85304 157292 85356 157344
rect 352564 157292 352616 157344
rect 355324 157292 355376 157344
rect 69848 154504 69900 154556
rect 71228 154504 71280 154556
rect 85304 154504 85356 154556
rect 87604 154504 87656 154556
rect 147680 153824 147732 153876
rect 159364 153824 159416 153876
rect 71780 153620 71832 153672
rect 75920 153620 75972 153672
rect 147496 153144 147548 153196
rect 149244 153144 149296 153196
rect 349804 153144 349856 153196
rect 356060 153212 356112 153264
rect 343640 151036 343692 151088
rect 349804 151036 349856 151088
rect 69756 150900 69808 150952
rect 72148 150900 72200 150952
rect 71228 150424 71280 150476
rect 72424 150424 72476 150476
rect 159364 149744 159416 149796
rect 166264 149744 166316 149796
rect 115572 149676 115624 149728
rect 580540 149676 580592 149728
rect 3148 149064 3200 149116
rect 25504 149064 25556 149116
rect 363696 148792 363748 148844
rect 366364 148792 366416 148844
rect 83464 148316 83516 148368
rect 88248 148316 88300 148368
rect 149244 148316 149296 148368
rect 155224 148316 155276 148368
rect 83556 147636 83608 147688
rect 171784 147636 171836 147688
rect 173164 147636 173216 147688
rect 341524 147636 341576 147688
rect 343640 147636 343692 147688
rect 86224 147568 86276 147620
rect 351184 146888 351236 146940
rect 363604 146888 363656 146940
rect 75920 146276 75972 146328
rect 80704 146208 80756 146260
rect 88340 144848 88392 144900
rect 89996 144848 90048 144900
rect 115480 144168 115532 144220
rect 580632 144168 580684 144220
rect 72148 142808 72200 142860
rect 91744 142808 91796 142860
rect 115940 142808 115992 142860
rect 477500 142808 477552 142860
rect 89996 141380 90048 141432
rect 98000 141380 98052 141432
rect 86224 141108 86276 141160
rect 91100 141108 91152 141160
rect 166264 141108 166316 141160
rect 169760 141108 169812 141160
rect 68284 140768 68336 140820
rect 71412 140700 71464 140752
rect 173164 140292 173216 140344
rect 177304 140292 177356 140344
rect 87604 139884 87656 139936
rect 89904 139884 89956 139936
rect 347044 139408 347096 139460
rect 351184 139408 351236 139460
rect 91744 138660 91796 138712
rect 97172 138660 97224 138712
rect 55864 138524 55916 138576
rect 57888 138524 57940 138576
rect 3424 138320 3476 138372
rect 4068 138320 4120 138372
rect 71412 137980 71464 138032
rect 80704 137980 80756 138032
rect 73160 137912 73212 137964
rect 114468 137980 114520 138032
rect 579620 137980 579672 138032
rect 86224 137912 86276 137964
rect 119344 137912 119396 137964
rect 120724 137912 120776 137964
rect 150532 137912 150584 137964
rect 152188 137912 152240 137964
rect 152464 137912 152516 137964
rect 153752 137912 153804 137964
rect 164516 137912 164568 137964
rect 172520 137912 172572 137964
rect 155224 137640 155276 137692
rect 164700 137640 164752 137692
rect 144460 137572 144512 137624
rect 156880 137572 156932 137624
rect 163504 137572 163556 137624
rect 174084 137572 174136 137624
rect 342260 137572 342312 137624
rect 352564 137572 352616 137624
rect 114192 137504 114244 137556
rect 396908 137504 396960 137556
rect 114284 137436 114336 137488
rect 397092 137436 397144 137488
rect 114376 137368 114428 137420
rect 397184 137368 397236 137420
rect 114100 137300 114152 137352
rect 398104 137300 398156 137352
rect 113916 137232 113968 137284
rect 542360 137232 542412 137284
rect 142436 137028 142488 137080
rect 145932 137028 145984 137080
rect 163596 136824 163648 136876
rect 170956 136824 171008 136876
rect 138112 136756 138164 136808
rect 142528 136756 142580 136808
rect 153476 136756 153528 136808
rect 155316 136756 155368 136808
rect 3424 136620 3476 136672
rect 115204 136620 115256 136672
rect 72424 136552 72476 136604
rect 73804 136552 73856 136604
rect 89904 136552 89956 136604
rect 95884 136552 95936 136604
rect 113732 136552 113784 136604
rect 116584 136552 116636 136604
rect 73160 136484 73212 136536
rect 75184 136484 75236 136536
rect 169760 136484 169812 136536
rect 175924 136484 175976 136536
rect 40040 136416 40092 136468
rect 175464 136416 175516 136468
rect 3976 136348 4028 136400
rect 178776 136348 178828 136400
rect 3792 136280 3844 136332
rect 178040 136280 178092 136332
rect 360844 136280 360896 136332
rect 363696 136280 363748 136332
rect 3884 136212 3936 136264
rect 178408 136212 178460 136264
rect 3700 136144 3752 136196
rect 178684 136144 178736 136196
rect 3240 136076 3292 136128
rect 178868 136076 178920 136128
rect 3332 136008 3384 136060
rect 178500 136008 178552 136060
rect 113824 135940 113876 135992
rect 412640 135940 412692 135992
rect 115388 135872 115440 135924
rect 580816 135872 580868 135924
rect 97172 135192 97224 135244
rect 102784 135192 102836 135244
rect 57888 134716 57940 134768
rect 176568 134716 176620 134768
rect 3608 134648 3660 134700
rect 178316 134648 178368 134700
rect 4068 134580 4120 134632
rect 178132 134580 178184 134632
rect 115296 134512 115348 134564
rect 342260 134512 342312 134564
rect 3792 133900 3844 133952
rect 175372 133900 175424 133952
rect 98000 133832 98052 133884
rect 101404 133832 101456 133884
rect 91100 133084 91152 133136
rect 93860 133084 93912 133136
rect 3424 131112 3476 131164
rect 113732 131112 113784 131164
rect 345664 131112 345716 131164
rect 347044 131112 347096 131164
rect 95884 130364 95936 130416
rect 108304 130364 108356 130416
rect 93860 128596 93912 128648
rect 97264 128596 97316 128648
rect 3608 128324 3660 128376
rect 113732 128324 113784 128376
rect 73804 127576 73856 127628
rect 82084 127576 82136 127628
rect 3700 126964 3752 127016
rect 113640 126964 113692 127016
rect 25504 126896 25556 126948
rect 113732 126896 113784 126948
rect 86224 126828 86276 126880
rect 88340 126828 88392 126880
rect 184204 125604 184256 125656
rect 579712 125604 579764 125656
rect 22836 125536 22888 125588
rect 113548 125536 113600 125588
rect 88340 125468 88392 125520
rect 90364 125468 90416 125520
rect 344284 124176 344336 124228
rect 345664 124176 345716 124228
rect 22744 124108 22796 124160
rect 113732 124108 113784 124160
rect 175924 124108 175976 124160
rect 178224 124108 178276 124160
rect 358084 124108 358136 124160
rect 360844 124108 360896 124160
rect 24124 122748 24176 122800
rect 113364 122748 113416 122800
rect 97264 121796 97316 121848
rect 98736 121796 98788 121848
rect 10324 121388 10376 121440
rect 113732 121388 113784 121440
rect 82084 121320 82136 121372
rect 85856 121320 85908 121372
rect 98736 121320 98788 121372
rect 100024 121320 100076 121372
rect 8944 120028 8996 120080
rect 113732 120028 113784 120080
rect 5080 118600 5132 118652
rect 113640 118600 113692 118652
rect 85856 117376 85908 117428
rect 87604 117376 87656 117428
rect 42064 117240 42116 117292
rect 113732 117240 113784 117292
rect 338764 117240 338816 117292
rect 341524 117240 341576 117292
rect 19984 115880 20036 115932
rect 113732 115880 113784 115932
rect 177304 115880 177356 115932
rect 178040 115880 178092 115932
rect 90364 115812 90416 115864
rect 93492 115812 93544 115864
rect 37924 113092 37976 113144
rect 113732 113092 113784 113144
rect 15844 111732 15896 111784
rect 113732 111732 113784 111784
rect 93492 111664 93544 111716
rect 96528 111664 96580 111716
rect 348424 111052 348476 111104
rect 358084 111052 358136 111104
rect 87604 110916 87656 110968
rect 88708 110916 88760 110968
rect 75184 110508 75236 110560
rect 77944 110508 77996 110560
rect 23480 110372 23532 110424
rect 113732 110372 113784 110424
rect 101404 109216 101456 109268
rect 102140 109216 102192 109268
rect 100024 108944 100076 108996
rect 102232 108944 102284 108996
rect 108304 108944 108356 108996
rect 113732 108944 113784 108996
rect 96528 108604 96580 108656
rect 97908 108604 97960 108656
rect 88708 107584 88760 107636
rect 113548 107584 113600 107636
rect 337016 106768 337068 106820
rect 338764 106768 338816 106820
rect 102232 106224 102284 106276
rect 113732 106224 113784 106276
rect 178040 106224 178092 106276
rect 344284 106224 344336 106276
rect 102140 105204 102192 105256
rect 104624 105204 104676 105256
rect 98000 104796 98052 104848
rect 113364 104796 113416 104848
rect 178040 104796 178092 104848
rect 337016 104796 337068 104848
rect 178040 103436 178092 103488
rect 413284 103436 413336 103488
rect 178040 102076 178092 102128
rect 410524 102076 410576 102128
rect 178040 100648 178092 100700
rect 409144 100648 409196 100700
rect 175924 99356 175976 99408
rect 580172 99356 580224 99408
rect 178040 99288 178092 99340
rect 407764 99288 407816 99340
rect 104624 98948 104676 99000
rect 106556 98948 106608 99000
rect 102784 97928 102836 97980
rect 105544 97928 105596 97980
rect 178040 97928 178092 97980
rect 406384 97928 406436 97980
rect 77944 96636 77996 96688
rect 81900 96568 81952 96620
rect 341524 95888 341576 95940
rect 348424 95888 348476 95940
rect 106556 95140 106608 95192
rect 108396 95140 108448 95192
rect 178040 95140 178092 95192
rect 405004 95140 405056 95192
rect 81900 93780 81952 93832
rect 84844 93780 84896 93832
rect 178040 93780 178092 93832
rect 403624 93780 403676 93832
rect 178040 92420 178092 92472
rect 400864 92420 400916 92472
rect 178040 90992 178092 91044
rect 399484 90992 399536 91044
rect 108396 90108 108448 90160
rect 109776 90108 109828 90160
rect 178040 89632 178092 89684
rect 418804 89632 418856 89684
rect 178040 88272 178092 88324
rect 417424 88272 417476 88324
rect 109776 86912 109828 86964
rect 110972 86912 111024 86964
rect 178040 86912 178092 86964
rect 414664 86912 414716 86964
rect 178684 85552 178736 85604
rect 580172 85552 580224 85604
rect 178040 85484 178092 85536
rect 188344 85484 188396 85536
rect 105544 84804 105596 84856
rect 116768 84804 116820 84856
rect 3332 84192 3384 84244
rect 116676 84192 116728 84244
rect 178040 84124 178092 84176
rect 185584 84124 185636 84176
rect 178040 82764 178092 82816
rect 184204 82764 184256 82816
rect 332600 82084 332652 82136
rect 341524 82084 341576 82136
rect 110972 79976 111024 80028
rect 115848 79976 115900 80028
rect 324320 79296 324372 79348
rect 332600 79296 332652 79348
rect 178040 75896 178092 75948
rect 562324 75896 562376 75948
rect 115940 75624 115992 75676
rect 120356 75624 120408 75676
rect 5264 75216 5316 75268
rect 141792 74876 141844 74928
rect 140964 74808 141016 74860
rect 170404 75624 170456 75676
rect 171324 75420 171376 75472
rect 171416 75420 171468 75472
rect 176568 75420 176620 75472
rect 171140 75352 171192 75404
rect 195980 75284 196032 75336
rect 156144 74876 156196 74928
rect 170496 75216 170548 75268
rect 171140 75148 171192 75200
rect 249800 75148 249852 75200
rect 171324 75080 171376 75132
rect 259460 75080 259512 75132
rect 156144 74740 156196 74792
rect 176384 75012 176436 75064
rect 324320 75012 324372 75064
rect 320180 74944 320232 74996
rect 338120 74876 338172 74928
rect 146484 74536 146536 74588
rect 147864 74604 147916 74656
rect 157524 74740 157576 74792
rect 167552 74808 167604 74860
rect 157524 74604 157576 74656
rect 167736 74740 167788 74792
rect 168564 74808 168616 74860
rect 176384 74808 176436 74860
rect 396816 74808 396868 74860
rect 176568 74740 176620 74792
rect 397000 74740 397052 74792
rect 390560 74672 390612 74724
rect 157800 74536 157852 74588
rect 465172 74604 465224 74656
rect 154764 74468 154816 74520
rect 167552 74536 167604 74588
rect 168196 74536 168248 74588
rect 579620 74536 579672 74588
rect 167092 74468 167144 74520
rect 580540 74468 580592 74520
rect 43444 74400 43496 74452
rect 169760 74400 169812 74452
rect 43536 74332 43588 74384
rect 169852 74332 169904 74384
rect 143724 74264 143776 74316
rect 284300 74264 284352 74316
rect 145104 74196 145156 74248
rect 302240 74196 302292 74248
rect 146760 74128 146812 74180
rect 324320 74128 324372 74180
rect 150624 74060 150676 74112
rect 374000 74060 374052 74112
rect 153384 73992 153436 74044
rect 408500 73992 408552 74044
rect 112444 73924 112496 73976
rect 115204 73856 115256 73908
rect 161664 73856 161716 73908
rect 116676 73720 116728 73772
rect 168380 73924 168432 73976
rect 462320 73924 462372 73976
rect 168288 73856 168340 73908
rect 527180 73856 527232 73908
rect 164424 73788 164476 73840
rect 550640 73788 550692 73840
rect 155500 73652 155552 73704
rect 5172 73584 5224 73636
rect 169944 73720 169996 73772
rect 168196 73652 168248 73704
rect 170496 73652 170548 73704
rect 84844 73516 84896 73568
rect 85580 73516 85632 73568
rect 131672 73380 131724 73432
rect 170128 73584 170180 73636
rect 161664 73516 161716 73568
rect 170036 73516 170088 73568
rect 167184 73448 167236 73500
rect 169576 73380 169628 73432
rect 131396 73244 131448 73296
rect 131672 73244 131724 73296
rect 120908 73108 120960 73160
rect 127900 73108 127952 73160
rect 131396 73108 131448 73160
rect 147864 73176 147916 73228
rect 153384 73176 153436 73228
rect 136824 73108 136876 73160
rect 156144 73108 156196 73160
rect 137652 73040 137704 73092
rect 207020 73176 207072 73228
rect 167920 73108 167972 73160
rect 168288 73108 168340 73160
rect 167828 73040 167880 73092
rect 580724 73040 580776 73092
rect 120724 72972 120776 73024
rect 128176 72972 128228 73024
rect 137744 72972 137796 73024
rect 145104 72972 145156 73024
rect 151820 72972 151872 73024
rect 152004 72972 152056 73024
rect 152740 72972 152792 73024
rect 168012 72972 168064 73024
rect 168472 72972 168524 73024
rect 397460 72972 397512 73024
rect 120816 72904 120868 72956
rect 129280 72904 129332 72956
rect 136272 72904 136324 72956
rect 147864 72904 147916 72956
rect 150256 72904 150308 72956
rect 119344 72836 119396 72888
rect 122748 72836 122800 72888
rect 141608 72836 141660 72888
rect 150624 72836 150676 72888
rect 153384 72904 153436 72956
rect 167920 72904 167972 72956
rect 168288 72904 168340 72956
rect 217324 72904 217376 72956
rect 154764 72836 154816 72888
rect 156604 72836 156656 72888
rect 231124 72836 231176 72888
rect 121092 72768 121144 72820
rect 130384 72768 130436 72820
rect 142712 72768 142764 72820
rect 151820 72768 151872 72820
rect 154396 72768 154448 72820
rect 121000 72700 121052 72752
rect 129832 72700 129884 72752
rect 140504 72700 140556 72752
rect 146760 72700 146812 72752
rect 151912 72700 151964 72752
rect 155500 72700 155552 72752
rect 86224 72632 86276 72684
rect 122380 72632 122432 72684
rect 122748 72632 122800 72684
rect 127348 72632 127400 72684
rect 132316 72632 132368 72684
rect 137744 72632 137796 72684
rect 138848 72632 138900 72684
rect 142712 72632 142764 72684
rect 85580 72564 85632 72616
rect 93952 72564 94004 72616
rect 60740 72496 60792 72548
rect 126336 72496 126388 72548
rect 25504 72428 25556 72480
rect 123116 72428 123168 72480
rect 121368 72360 121420 72412
rect 132684 72564 132736 72616
rect 139216 72564 139268 72616
rect 152924 72632 152976 72684
rect 157432 72768 157484 72820
rect 239220 72768 239272 72820
rect 158260 72700 158312 72752
rect 158628 72700 158680 72752
rect 166632 72700 166684 72752
rect 259368 72700 259420 72752
rect 422300 72632 422352 72684
rect 151268 72564 151320 72616
rect 154120 72564 154172 72616
rect 158628 72564 158680 72616
rect 471980 72564 472032 72616
rect 134708 72496 134760 72548
rect 149980 72496 150032 72548
rect 152004 72496 152056 72548
rect 156604 72496 156656 72548
rect 166724 72496 166776 72548
rect 520924 72496 520976 72548
rect 135720 72428 135772 72480
rect 165252 72428 165304 72480
rect 166908 72428 166960 72480
rect 580264 72428 580316 72480
rect 142160 72360 142212 72412
rect 152924 72360 152976 72412
rect 156052 72360 156104 72412
rect 171784 72360 171836 72412
rect 133972 72292 134024 72344
rect 137652 72292 137704 72344
rect 150808 72292 150860 72344
rect 152832 72292 152884 72344
rect 145472 72224 145524 72276
rect 116676 72156 116728 72208
rect 124864 72156 124916 72208
rect 142712 72156 142764 72208
rect 150164 72156 150216 72208
rect 118148 72088 118200 72140
rect 124312 72088 124364 72140
rect 151820 72224 151872 72276
rect 153016 72224 153068 72276
rect 152188 72156 152240 72208
rect 167644 72292 167696 72344
rect 154948 72224 155000 72276
rect 169024 72224 169076 72276
rect 153844 72156 153896 72208
rect 167736 72156 167788 72208
rect 154304 72088 154356 72140
rect 117964 72020 118016 72072
rect 123760 72020 123812 72072
rect 145104 72020 145156 72072
rect 146024 72020 146076 72072
rect 151360 72020 151412 72072
rect 158444 72020 158496 72072
rect 118056 71952 118108 72004
rect 123024 71952 123076 72004
rect 149152 71952 149204 72004
rect 154396 71952 154448 72004
rect 149704 71884 149756 71936
rect 156880 71884 156932 71936
rect 127716 71816 127768 71868
rect 128084 71816 128136 71868
rect 146760 71816 146812 71868
rect 151636 71816 151688 71868
rect 153292 71816 153344 71868
rect 167368 72088 167420 72140
rect 162768 72020 162820 72072
rect 166724 72020 166776 72072
rect 165068 71816 165120 71868
rect 166632 71816 166684 71868
rect 132500 71748 132552 71800
rect 136180 71748 136232 71800
rect 136640 71748 136692 71800
rect 143264 71748 143316 71800
rect 145840 71748 145892 71800
rect 147312 71748 147364 71800
rect 3516 71680 3568 71732
rect 178592 72020 178644 72072
rect 167276 71952 167328 72004
rect 580172 71952 580224 72004
rect 93952 71612 94004 71664
rect 168656 71612 168708 71664
rect 127624 71544 127676 71596
rect 168748 71544 168800 71596
rect 116768 71068 116820 71120
rect 168932 71476 168984 71528
rect 116584 70932 116636 70984
rect 127624 70932 127676 70984
rect 120356 70864 120408 70916
rect 168840 71408 168892 71460
rect 259368 71000 259420 71052
rect 581092 71000 581144 71052
rect 123024 69912 123076 69964
rect 123576 69912 123628 69964
rect 129096 69912 129148 69964
rect 129648 69912 129700 69964
rect 138756 69912 138808 69964
rect 121920 69844 121972 69896
rect 122564 69844 122616 69896
rect 125784 69844 125836 69896
rect 126612 69844 126664 69896
rect 122380 69776 122432 69828
rect 122656 69776 122708 69828
rect 122932 69776 122984 69828
rect 124128 69776 124180 69828
rect 123116 69708 123168 69760
rect 123852 69708 123904 69760
rect 121736 69640 121788 69692
rect 122196 69640 122248 69692
rect 123208 69640 123260 69692
rect 123760 69640 123812 69692
rect 124956 69776 125008 69828
rect 126060 69708 126112 69760
rect 126612 69708 126664 69760
rect 126336 69640 126388 69692
rect 126796 69640 126848 69692
rect 127716 69640 127768 69692
rect 128176 69640 128228 69692
rect 128544 69640 128596 69692
rect 128820 69640 128872 69692
rect 129004 69640 129056 69692
rect 129188 69640 129240 69692
rect 130476 69844 130528 69896
rect 130108 69776 130160 69828
rect 130568 69776 130620 69828
rect 138112 69776 138164 69828
rect 122104 69572 122156 69624
rect 122564 69572 122616 69624
rect 123392 69572 123444 69624
rect 123944 69572 123996 69624
rect 124588 69572 124640 69624
rect 125692 69572 125744 69624
rect 126888 69572 126940 69624
rect 128636 69572 128688 69624
rect 129740 69572 129792 69624
rect 130016 69572 130068 69624
rect 124496 69504 124548 69556
rect 125324 69504 125376 69556
rect 138756 69640 138808 69692
rect 156604 69640 156656 69692
rect 156972 69640 157024 69692
rect 167552 69640 167604 69692
rect 130200 69572 130252 69624
rect 130568 69572 130620 69624
rect 130936 69572 130988 69624
rect 138664 69572 138716 69624
rect 167276 69572 167328 69624
rect 130476 69504 130528 69556
rect 124864 69436 124916 69488
rect 125416 69436 125468 69488
rect 130108 69436 130160 69488
rect 130844 69436 130896 69488
rect 167552 69436 167604 69488
rect 167920 69436 167972 69488
rect 154764 68824 154816 68876
rect 158352 68824 158404 68876
rect 131396 68280 131448 68332
rect 239220 68280 239272 68332
rect 460940 68280 460992 68332
rect 127440 68144 127492 68196
rect 131304 67940 131356 67992
rect 127348 67872 127400 67924
rect 123300 67804 123352 67856
rect 123668 67804 123720 67856
rect 125968 67804 126020 67856
rect 126244 67804 126296 67856
rect 127440 67804 127492 67856
rect 127900 67804 127952 67856
rect 128728 67804 128780 67856
rect 129096 67804 129148 67856
rect 127256 67736 127308 67788
rect 128268 67736 128320 67788
rect 129004 67736 129056 67788
rect 129556 67736 129608 67788
rect 123668 67668 123720 67720
rect 124036 67668 124088 67720
rect 128728 67668 128780 67720
rect 129464 67668 129516 67720
rect 126060 67532 126112 67584
rect 126428 67532 126480 67584
rect 125968 67464 126020 67516
rect 126704 67464 126756 67516
rect 5540 66852 5592 66904
rect 122012 67192 122064 67244
rect 121644 66852 121696 66904
rect 122288 66852 122340 66904
rect 122196 66784 122248 66836
rect 122748 66784 122800 66836
rect 124772 66172 124824 66224
rect 125048 66172 125100 66224
rect 114376 60664 114428 60716
rect 580172 60664 580224 60716
rect 163504 58624 163556 58676
rect 326344 58624 326396 58676
rect 15200 54476 15252 54528
rect 119344 54476 119396 54528
rect 113180 51076 113232 51128
rect 121092 51076 121144 51128
rect 178684 46860 178736 46912
rect 580172 46860 580224 46912
rect 3516 45500 3568 45552
rect 170220 45500 170272 45552
rect 106280 43392 106332 43444
rect 121000 43392 121052 43444
rect 153108 40672 153160 40724
rect 226340 40672 226392 40724
rect 155500 36660 155552 36712
rect 390652 36660 390704 36712
rect 152464 36592 152516 36644
rect 397460 36592 397512 36644
rect 157800 36524 157852 36576
rect 456800 36524 456852 36576
rect 145564 35844 145616 35896
rect 307760 35844 307812 35896
rect 147312 35776 147364 35828
rect 311900 35776 311952 35828
rect 146392 35708 146444 35760
rect 318800 35708 318852 35760
rect 146668 35640 146720 35692
rect 322940 35640 322992 35692
rect 146944 35572 146996 35624
rect 325700 35572 325752 35624
rect 147772 35504 147824 35556
rect 336740 35504 336792 35556
rect 148600 35436 148652 35488
rect 347780 35436 347832 35488
rect 154488 35368 154540 35420
rect 354680 35368 354732 35420
rect 149428 35300 149480 35352
rect 357440 35300 357492 35352
rect 158352 35232 158404 35284
rect 368480 35232 368532 35284
rect 158444 35164 158496 35216
rect 382280 35164 382332 35216
rect 145288 35096 145340 35148
rect 305000 35096 305052 35148
rect 138664 34416 138716 34468
rect 212540 34416 212592 34468
rect 138388 34348 138440 34400
rect 216680 34348 216732 34400
rect 138848 34280 138900 34332
rect 219440 34280 219492 34332
rect 139768 34212 139820 34264
rect 234620 34212 234672 34264
rect 140872 34144 140924 34196
rect 248420 34144 248472 34196
rect 141424 34076 141476 34128
rect 255320 34076 255372 34128
rect 142528 34008 142580 34060
rect 269120 34008 269172 34060
rect 143080 33940 143132 33992
rect 276020 33940 276072 33992
rect 143632 33872 143684 33924
rect 284392 33872 284444 33924
rect 144184 33804 144236 33856
rect 291200 33804 291252 33856
rect 145012 33736 145064 33788
rect 300860 33736 300912 33788
rect 2872 33056 2924 33108
rect 175556 33056 175608 33108
rect 135352 32920 135404 32972
rect 176660 32920 176712 32972
rect 135628 32852 135680 32904
rect 180800 32852 180852 32904
rect 135904 32784 135956 32836
rect 184940 32784 184992 32836
rect 136732 32716 136784 32768
rect 194600 32716 194652 32768
rect 137008 32648 137060 32700
rect 198740 32648 198792 32700
rect 137560 32580 137612 32632
rect 205640 32580 205692 32632
rect 142252 32512 142304 32564
rect 266360 32512 266412 32564
rect 164332 32444 164384 32496
rect 549260 32444 549312 32496
rect 166264 32376 166316 32428
rect 574100 32376 574152 32428
rect 157616 31696 157668 31748
rect 463700 31696 463752 31748
rect 158168 31628 158220 31680
rect 470600 31628 470652 31680
rect 158720 31560 158772 31612
rect 477500 31560 477552 31612
rect 159088 31492 159140 31544
rect 481640 31492 481692 31544
rect 161020 31424 161072 31476
rect 490012 31424 490064 31476
rect 160192 31356 160244 31408
rect 496820 31356 496872 31408
rect 160744 31288 160796 31340
rect 503720 31288 503772 31340
rect 162584 31220 162636 31272
rect 510620 31220 510672 31272
rect 161848 31152 161900 31204
rect 517520 31152 517572 31204
rect 166724 31084 166776 31136
rect 524420 31084 524472 31136
rect 162124 31016 162176 31068
rect 521660 31016 521712 31068
rect 154304 30268 154356 30320
rect 307852 30268 307904 30320
rect 144920 30200 144972 30252
rect 299480 30200 299532 30252
rect 145196 30132 145248 30184
rect 303620 30132 303672 30184
rect 150716 30064 150768 30116
rect 374092 30064 374144 30116
rect 154212 29996 154264 30048
rect 382372 29996 382424 30048
rect 156972 29928 157024 29980
rect 389180 29928 389232 29980
rect 155132 29860 155184 29912
rect 431960 29860 432012 29912
rect 157064 29792 157116 29844
rect 438860 29792 438912 29844
rect 155960 29724 156012 29776
rect 441620 29724 441672 29776
rect 156236 29656 156288 29708
rect 445760 29656 445812 29708
rect 156788 29588 156840 29640
rect 452660 29588 452712 29640
rect 139400 28908 139452 28960
rect 229100 28908 229152 28960
rect 151544 28840 151596 28892
rect 242900 28840 242952 28892
rect 140228 28772 140280 28824
rect 240140 28772 240192 28824
rect 140780 28704 140832 28756
rect 247040 28704 247092 28756
rect 150624 28636 150676 28688
rect 258080 28636 258132 28688
rect 141056 28568 141108 28620
rect 251180 28568 251232 28620
rect 152924 28500 152976 28552
rect 264980 28500 265032 28552
rect 153016 28432 153068 28484
rect 271880 28432 271932 28484
rect 150440 28364 150492 28416
rect 371240 28364 371292 28416
rect 152832 28296 152884 28348
rect 375380 28296 375432 28348
rect 165988 28228 166040 28280
rect 571340 28228 571392 28280
rect 138296 28160 138348 28212
rect 215300 28160 215352 28212
rect 138112 28092 138164 28144
rect 211160 28092 211212 28144
rect 150164 28024 150216 28076
rect 222200 28024 222252 28076
rect 143264 27548 143316 27600
rect 193220 27548 193272 27600
rect 136088 27480 136140 27532
rect 186320 27480 186372 27532
rect 136916 27412 136968 27464
rect 197360 27412 197412 27464
rect 146024 27344 146076 27396
rect 208400 27344 208452 27396
rect 137192 27276 137244 27328
rect 201500 27276 201552 27328
rect 137468 27208 137520 27260
rect 204260 27208 204312 27260
rect 138572 27140 138624 27192
rect 218060 27140 218112 27192
rect 139676 27072 139728 27124
rect 233240 27072 233292 27124
rect 148324 27004 148376 27056
rect 343640 27004 343692 27056
rect 154580 26936 154632 26988
rect 423680 26936 423732 26988
rect 157984 26868 158036 26920
rect 467840 26868 467892 26920
rect 135812 26188 135864 26240
rect 183560 26188 183612 26240
rect 139952 26120 140004 26172
rect 236000 26120 236052 26172
rect 141884 26052 141936 26104
rect 260840 26052 260892 26104
rect 144368 25984 144420 26036
rect 292580 25984 292632 26036
rect 149336 25916 149388 25968
rect 357532 25916 357584 25968
rect 150532 25848 150584 25900
rect 372620 25848 372672 25900
rect 153752 25780 153804 25832
rect 414020 25780 414072 25832
rect 164792 25712 164844 25764
rect 556160 25712 556212 25764
rect 166632 25644 166684 25696
rect 558920 25644 558972 25696
rect 165620 25576 165672 25628
rect 565820 25576 565872 25628
rect 81440 25508 81492 25560
rect 120908 25508 120960 25560
rect 166172 25508 166224 25560
rect 572720 25508 572772 25560
rect 135536 25440 135588 25492
rect 179420 25440 179472 25492
rect 135260 25372 135312 25424
rect 176752 25372 176804 25424
rect 141332 24760 141384 24812
rect 253940 24760 253992 24812
rect 143540 24692 143592 24744
rect 282920 24692 282972 24744
rect 153200 24624 153252 24676
rect 407212 24624 407264 24676
rect 162860 24556 162912 24608
rect 531320 24556 531372 24608
rect 163136 24488 163188 24540
rect 534080 24488 534132 24540
rect 163412 24420 163464 24472
rect 538220 24420 538272 24472
rect 163688 24352 163740 24404
rect 540980 24352 541032 24404
rect 164240 24284 164292 24336
rect 547880 24284 547932 24336
rect 164516 24216 164568 24268
rect 552020 24216 552072 24268
rect 165712 24148 165764 24200
rect 567200 24148 567252 24200
rect 165896 24080 165948 24132
rect 569960 24080 570012 24132
rect 157340 23400 157392 23452
rect 459560 23400 459612 23452
rect 160100 23332 160152 23384
rect 495440 23332 495492 23384
rect 160376 23264 160428 23316
rect 498292 23264 498344 23316
rect 160652 23196 160704 23248
rect 502340 23196 502392 23248
rect 160928 23128 160980 23180
rect 506480 23128 506532 23180
rect 161480 23060 161532 23112
rect 513380 23060 513432 23112
rect 161756 22992 161808 23044
rect 516140 22992 516192 23044
rect 162032 22924 162084 22976
rect 520280 22924 520332 22976
rect 162308 22856 162360 22908
rect 523040 22856 523092 22908
rect 165160 22788 165212 22840
rect 560300 22788 560352 22840
rect 114468 22720 114520 22772
rect 580172 22720 580224 22772
rect 3516 22652 3568 22704
rect 170312 22652 170364 22704
rect 148048 21972 148100 22024
rect 340880 21972 340932 22024
rect 156880 21904 156932 21956
rect 361580 21904 361632 21956
rect 155040 21836 155092 21888
rect 430580 21836 430632 21888
rect 155224 21768 155276 21820
rect 432052 21768 432104 21820
rect 156328 21700 156380 21752
rect 447140 21700 447192 21752
rect 156420 21632 156472 21684
rect 448520 21632 448572 21684
rect 158996 21564 159048 21616
rect 481732 21564 481784 21616
rect 159272 21496 159324 21548
rect 484400 21496 484452 21548
rect 159548 21428 159600 21480
rect 488540 21428 488592 21480
rect 159824 21360 159876 21412
rect 491300 21360 491352 21412
rect 140044 20408 140096 20460
rect 237380 20408 237432 20460
rect 141700 20340 141752 20392
rect 259552 20340 259604 20392
rect 147220 20272 147272 20324
rect 329840 20272 329892 20324
rect 139492 20204 139544 20256
rect 230480 20204 230532 20256
rect 231124 20204 231176 20256
rect 449900 20204 449952 20256
rect 152280 20136 152332 20188
rect 394700 20136 394752 20188
rect 152556 20068 152608 20120
rect 398840 20068 398892 20120
rect 153660 20000 153712 20052
rect 412640 20000 412692 20052
rect 158076 19932 158128 19984
rect 469220 19932 469272 19984
rect 141148 19048 141200 19100
rect 251272 19048 251324 19100
rect 163780 18980 163832 19032
rect 312544 18980 312596 19032
rect 149520 18912 149572 18964
rect 358820 18912 358872 18964
rect 150900 18844 150952 18896
rect 376760 18844 376812 18896
rect 151176 18776 151228 18828
rect 380900 18776 380952 18828
rect 156696 18708 156748 18760
rect 451280 18708 451332 18760
rect 163228 18640 163280 18692
rect 535460 18640 535512 18692
rect 35900 18572 35952 18624
rect 118148 18572 118200 18624
rect 164608 18572 164660 18624
rect 553400 18572 553452 18624
rect 142804 17620 142856 17672
rect 273260 17620 273312 17672
rect 147036 17552 147088 17604
rect 327080 17552 327132 17604
rect 154856 17484 154908 17536
rect 427820 17484 427872 17536
rect 155316 17416 155368 17468
rect 433340 17416 433392 17468
rect 155408 17348 155460 17400
rect 434720 17348 434772 17400
rect 155592 17280 155644 17332
rect 437480 17280 437532 17332
rect 164884 17212 164936 17264
rect 556252 17212 556304 17264
rect 142896 16396 142948 16448
rect 274824 16396 274876 16448
rect 143908 16328 143960 16380
rect 287336 16328 287388 16380
rect 144000 16260 144052 16312
rect 288992 16260 289044 16312
rect 144276 16192 144328 16244
rect 292672 16192 292724 16244
rect 148508 16124 148560 16176
rect 346952 16124 347004 16176
rect 149060 16056 149112 16108
rect 353576 16056 353628 16108
rect 153936 15988 153988 16040
rect 415492 15988 415544 16040
rect 171784 15920 171836 15972
rect 443368 15920 443420 15972
rect 162952 15852 163004 15904
rect 532056 15852 532108 15904
rect 141240 14900 141292 14952
rect 253480 14900 253532 14952
rect 141516 14832 141568 14884
rect 256700 14832 256752 14884
rect 142344 14764 142396 14816
rect 267740 14764 267792 14816
rect 142620 14696 142672 14748
rect 270776 14696 270828 14748
rect 149612 14628 149664 14680
rect 361120 14628 361172 14680
rect 151452 14560 151504 14612
rect 384304 14560 384356 14612
rect 154672 14492 154724 14544
rect 425704 14492 425756 14544
rect 157892 14424 157944 14476
rect 467472 14424 467524 14476
rect 139584 13404 139636 13456
rect 231860 13404 231912 13456
rect 140136 13336 140188 13388
rect 239312 13336 239364 13388
rect 146852 13268 146904 13320
rect 324412 13268 324464 13320
rect 147128 13200 147180 13252
rect 328736 13200 328788 13252
rect 149796 13132 149848 13184
rect 363512 13132 363564 13184
rect 14280 13064 14332 13116
rect 122104 13064 122156 13116
rect 150992 13064 151044 13116
rect 378416 13064 378468 13116
rect 157708 12248 157760 12300
rect 169116 12248 169168 12300
rect 138204 12180 138256 12232
rect 214472 12180 214524 12232
rect 138480 12112 138532 12164
rect 218152 12112 218204 12164
rect 138756 12044 138808 12096
rect 221096 12044 221148 12096
rect 146576 11976 146628 12028
rect 322112 11976 322164 12028
rect 148232 11908 148284 11960
rect 342904 11908 342956 11960
rect 148416 11840 148468 11892
rect 345296 11840 345348 11892
rect 149244 11772 149296 11824
rect 356336 11772 356388 11824
rect 159364 11704 159416 11756
rect 486424 11704 486476 11756
rect 176660 11636 176712 11688
rect 177856 11636 177908 11688
rect 218060 11636 218112 11688
rect 219256 11636 219308 11688
rect 242900 11636 242952 11688
rect 244096 11636 244148 11688
rect 259460 11636 259512 11688
rect 260656 11636 260708 11688
rect 110512 10956 110564 11008
rect 130476 10956 130528 11008
rect 102140 10888 102192 10940
rect 129004 10888 129056 10940
rect 95792 10820 95844 10872
rect 129188 10820 129240 10872
rect 134800 10820 134852 10872
rect 170312 10820 170364 10872
rect 92480 10752 92532 10804
rect 129096 10752 129148 10804
rect 137100 10752 137152 10804
rect 200304 10752 200356 10804
rect 75000 10684 75052 10736
rect 122196 10684 122248 10736
rect 137376 10684 137428 10736
rect 203432 10684 203484 10736
rect 78128 10616 78180 10668
rect 127808 10616 127860 10668
rect 142988 10616 143040 10668
rect 276112 10616 276164 10668
rect 67640 10548 67692 10600
rect 126336 10548 126388 10600
rect 144460 10548 144512 10600
rect 294880 10548 294932 10600
rect 64328 10480 64380 10532
rect 126428 10480 126480 10532
rect 145932 10480 145984 10532
rect 313832 10480 313884 10532
rect 46664 10412 46716 10464
rect 125048 10412 125100 10464
rect 146300 10412 146352 10464
rect 318064 10412 318116 10464
rect 31944 10344 31996 10396
rect 123668 10344 123720 10396
rect 152648 10344 152700 10396
rect 398932 10344 398984 10396
rect 25320 10276 25372 10328
rect 123576 10276 123628 10328
rect 156512 10276 156564 10328
rect 448612 10276 448664 10328
rect 117320 10208 117372 10260
rect 130384 10208 130436 10260
rect 120632 10140 120684 10192
rect 130568 10140 130620 10192
rect 116400 9596 116452 9648
rect 130200 9596 130252 9648
rect 135444 9596 135496 9648
rect 179052 9596 179104 9648
rect 112812 9528 112864 9580
rect 130292 9528 130344 9580
rect 135996 9528 136048 9580
rect 186136 9528 186188 9580
rect 60832 9460 60884 9512
rect 126152 9460 126204 9512
rect 145380 9460 145432 9512
rect 306748 9460 306800 9512
rect 57244 9392 57296 9444
rect 126244 9392 126296 9444
rect 145656 9392 145708 9444
rect 310244 9392 310296 9444
rect 43076 9324 43128 9376
rect 116676 9324 116728 9376
rect 145748 9324 145800 9376
rect 311440 9324 311492 9376
rect 50160 9256 50212 9308
rect 124864 9256 124916 9308
rect 147956 9256 148008 9308
rect 339868 9256 339920 9308
rect 45468 9188 45520 9240
rect 124772 9188 124824 9240
rect 148140 9188 148192 9240
rect 342168 9188 342220 9240
rect 41880 9120 41932 9172
rect 124956 9120 125008 9172
rect 152096 9120 152148 9172
rect 393044 9120 393096 9172
rect 31300 9052 31352 9104
rect 123392 9052 123444 9104
rect 153476 9052 153528 9104
rect 410800 9052 410852 9104
rect 24216 8984 24268 9036
rect 123484 8984 123536 9036
rect 153568 8984 153620 9036
rect 411904 8984 411956 9036
rect 9956 8916 10008 8968
rect 122012 8916 122064 8968
rect 166080 8916 166132 8968
rect 572720 8916 572772 8968
rect 134892 8848 134944 8900
rect 171968 8848 172020 8900
rect 98644 8236 98696 8288
rect 128912 8236 128964 8288
rect 95148 8168 95200 8220
rect 128820 8168 128872 8220
rect 84476 8100 84528 8152
rect 127716 8100 127768 8152
rect 80888 8032 80940 8084
rect 127440 8032 127492 8084
rect 77392 7964 77444 8016
rect 127624 7964 127676 8016
rect 142436 7964 142488 8016
rect 268844 7964 268896 8016
rect 73804 7896 73856 7948
rect 127532 7896 127584 7948
rect 144092 7896 144144 7948
rect 290188 7896 290240 7948
rect 66720 7828 66772 7880
rect 125968 7828 126020 7880
rect 147680 7828 147732 7880
rect 336280 7828 336332 7880
rect 63224 7760 63276 7812
rect 126060 7760 126112 7812
rect 154028 7760 154080 7812
rect 417884 7760 417936 7812
rect 27712 7692 27764 7744
rect 123300 7692 123352 7744
rect 164700 7692 164752 7744
rect 554964 7692 555016 7744
rect 19432 7624 19484 7676
rect 118056 7624 118108 7676
rect 119896 7624 119948 7676
rect 130108 7624 130160 7676
rect 164976 7624 165028 7676
rect 558552 7624 558604 7676
rect 23020 7556 23072 7608
rect 123208 7556 123260 7608
rect 165804 7556 165856 7608
rect 569132 7556 569184 7608
rect 102232 7488 102284 7540
rect 128728 7488 128780 7540
rect 481640 7488 481692 7540
rect 482468 7488 482520 7540
rect 115204 6808 115256 6860
rect 130016 6808 130068 6860
rect 562324 6808 562376 6860
rect 580172 6808 580224 6860
rect 99840 6740 99892 6792
rect 120816 6740 120868 6792
rect 59636 6672 59688 6724
rect 125876 6672 125928 6724
rect 139860 6672 139912 6724
rect 235816 6672 235868 6724
rect 11152 6604 11204 6656
rect 86224 6604 86276 6656
rect 104532 6604 104584 6656
rect 128636 6604 128688 6656
rect 143816 6604 143868 6656
rect 286600 6604 286652 6656
rect 48964 6536 49016 6588
rect 124496 6536 124548 6588
rect 151084 6536 151136 6588
rect 379980 6536 380032 6588
rect 44272 6468 44324 6520
rect 124588 6468 124640 6520
rect 152372 6468 152424 6520
rect 396540 6468 396592 6520
rect 40684 6400 40736 6452
rect 124680 6400 124732 6452
rect 169024 6400 169076 6452
rect 429660 6400 429712 6452
rect 30104 6332 30156 6384
rect 123116 6332 123168 6384
rect 167184 6332 167236 6384
rect 436744 6332 436796 6384
rect 13544 6264 13596 6316
rect 121920 6264 121972 6316
rect 161572 6264 161624 6316
rect 514760 6264 514812 6316
rect 8760 6196 8812 6248
rect 121736 6196 121788 6248
rect 163596 6196 163648 6248
rect 540796 6196 540848 6248
rect 4068 6128 4120 6180
rect 121828 6128 121880 6180
rect 163872 6128 163924 6180
rect 544384 6128 544436 6180
rect 97448 5448 97500 5500
rect 129648 5448 129700 5500
rect 93952 5380 94004 5432
rect 128544 5380 128596 5432
rect 132592 5380 132644 5432
rect 142436 5380 142488 5432
rect 85672 5312 85724 5364
rect 120724 5312 120776 5364
rect 132776 5312 132828 5364
rect 144736 5312 144788 5364
rect 86868 5244 86920 5296
rect 127256 5244 127308 5296
rect 134524 5244 134576 5296
rect 167184 5244 167236 5296
rect 76196 5176 76248 5228
rect 127348 5176 127400 5228
rect 137284 5176 137336 5228
rect 202696 5176 202748 5228
rect 72608 5108 72660 5160
rect 127164 5108 127216 5160
rect 133052 5108 133104 5160
rect 148324 5108 148376 5160
rect 149888 5108 149940 5160
rect 364616 5108 364668 5160
rect 405004 5108 405056 5160
rect 479340 5108 479392 5160
rect 65524 5040 65576 5092
rect 125784 5040 125836 5092
rect 133144 5040 133196 5092
rect 149520 5040 149572 5092
rect 160468 5040 160520 5092
rect 500592 5040 500644 5092
rect 33600 4972 33652 5024
rect 122932 4972 122984 5024
rect 133420 4972 133472 5024
rect 153016 4972 153068 5024
rect 160560 4972 160612 5024
rect 501788 4972 501840 5024
rect 28908 4904 28960 4956
rect 117964 4904 118016 4956
rect 118792 4904 118844 4956
rect 130844 4904 130896 4956
rect 133328 4904 133380 4956
rect 151820 4904 151872 4956
rect 161940 4904 161992 4956
rect 519544 4904 519596 4956
rect 5264 4836 5316 4888
rect 22744 4836 22796 4888
rect 26516 4836 26568 4888
rect 123024 4836 123076 4888
rect 133880 4836 133932 4888
rect 158904 4836 158956 4888
rect 162216 4836 162268 4888
rect 523040 4836 523092 4888
rect 21824 4768 21876 4820
rect 123760 4768 123812 4820
rect 134248 4768 134300 4820
rect 163688 4768 163740 4820
rect 166908 4768 166960 4820
rect 577412 4768 577464 4820
rect 111616 4700 111668 4752
rect 129924 4700 129976 4752
rect 117228 4632 117280 4684
rect 129372 4632 129424 4684
rect 101036 4088 101088 4140
rect 117228 4088 117280 4140
rect 121368 4088 121420 4140
rect 143540 4088 143592 4140
rect 167552 4088 167604 4140
rect 189724 4088 189776 4140
rect 276020 4088 276072 4140
rect 276756 4088 276808 4140
rect 284300 4088 284352 4140
rect 285036 4088 285088 4140
rect 292580 4088 292632 4140
rect 293316 4088 293368 4140
rect 312544 4088 312596 4140
rect 543188 4088 543240 4140
rect 83280 4020 83332 4072
rect 127992 4020 128044 4072
rect 131856 4020 131908 4072
rect 132960 4020 133012 4072
rect 79692 3952 79744 4004
rect 128084 3952 128136 4004
rect 132868 3952 132920 4004
rect 134064 3952 134116 4004
rect 146944 4020 146996 4072
rect 160100 4020 160152 4072
rect 168104 4020 168156 4072
rect 401324 4020 401376 4072
rect 69112 3884 69164 3936
rect 125692 3884 125744 3936
rect 132040 3884 132092 3936
rect 135260 3884 135312 3936
rect 145932 3952 145984 4004
rect 167368 3952 167420 4004
rect 408408 3952 408460 4004
rect 161296 3884 161348 3936
rect 167644 3884 167696 3936
rect 415400 3884 415452 3936
rect 58440 3816 58492 3868
rect 126612 3816 126664 3868
rect 134156 3816 134208 3868
rect 162492 3816 162544 3868
rect 167276 3816 167328 3868
rect 427268 3816 427320 3868
rect 51356 3748 51408 3800
rect 125508 3748 125560 3800
rect 134340 3748 134392 3800
rect 164884 3748 164936 3800
rect 168196 3748 168248 3800
rect 445024 3748 445076 3800
rect 445116 3748 445168 3800
rect 546684 3748 546736 3800
rect 47860 3680 47912 3732
rect 125324 3680 125376 3732
rect 134432 3680 134484 3732
rect 166080 3680 166132 3732
rect 167736 3680 167788 3732
rect 462780 3680 462832 3732
rect 39580 3612 39632 3664
rect 124312 3612 124364 3664
rect 134616 3612 134668 3664
rect 168380 3612 168432 3664
rect 169116 3612 169168 3664
rect 465172 3612 465224 3664
rect 12348 3544 12400 3596
rect 122656 3544 122708 3596
rect 133052 3544 133104 3596
rect 147128 3544 147180 3596
rect 159180 3544 159232 3596
rect 484032 3544 484084 3596
rect 7656 3476 7708 3528
rect 122564 3476 122616 3528
rect 125876 3476 125928 3528
rect 131212 3476 131264 3528
rect 133236 3476 133288 3528
rect 150624 3476 150676 3528
rect 159456 3476 159508 3528
rect 478052 3476 478104 3528
rect 2872 3408 2924 3460
rect 122196 3408 122248 3460
rect 126980 3408 127032 3460
rect 131580 3408 131632 3460
rect 133512 3408 133564 3460
rect 154212 3408 154264 3460
rect 159732 3408 159784 3460
rect 491116 3408 491168 3460
rect 520924 3408 520976 3460
rect 582196 3408 582248 3460
rect 102140 3340 102192 3392
rect 103336 3340 103388 3392
rect 122288 3340 122340 3392
rect 131028 3340 131080 3392
rect 131948 3340 132000 3392
rect 134156 3340 134208 3392
rect 137744 3340 137796 3392
rect 146944 3340 146996 3392
rect 167460 3340 167512 3392
rect 394240 3340 394292 3392
rect 398932 3340 398984 3392
rect 400128 3340 400180 3392
rect 415492 3340 415544 3392
rect 416688 3340 416740 3392
rect 423680 3340 423732 3392
rect 424968 3340 425020 3392
rect 440332 3340 440384 3392
rect 441528 3340 441580 3392
rect 448612 3340 448664 3392
rect 449808 3340 449860 3392
rect 456800 3340 456852 3392
rect 458088 3340 458140 3392
rect 473360 3340 473412 3392
rect 474188 3340 474240 3392
rect 478052 3340 478104 3392
rect 487620 3340 487672 3392
rect 132132 3272 132184 3324
rect 136456 3272 136508 3324
rect 150072 3272 150124 3324
rect 169576 3272 169628 3324
rect 169668 3272 169720 3324
rect 175464 3272 175516 3324
rect 193220 3272 193272 3324
rect 194416 3272 194468 3324
rect 226340 3272 226392 3324
rect 227536 3272 227588 3324
rect 299480 3272 299532 3324
rect 300768 3272 300820 3324
rect 307760 3272 307812 3324
rect 309048 3272 309100 3324
rect 316040 3272 316092 3324
rect 317328 3272 317380 3324
rect 324412 3272 324464 3324
rect 325608 3272 325660 3324
rect 332600 3272 332652 3324
rect 333888 3272 333940 3324
rect 20628 3204 20680 3256
rect 25504 3204 25556 3256
rect 165252 3204 165304 3256
rect 182548 3204 182600 3256
rect 326436 3204 326488 3256
rect 539600 3272 539652 3324
rect 349160 3204 349212 3256
rect 350448 3204 350500 3256
rect 357440 3204 357492 3256
rect 358728 3204 358780 3256
rect 365720 3204 365772 3256
rect 367008 3204 367060 3256
rect 374092 3204 374144 3256
rect 375288 3204 375340 3256
rect 382280 3204 382332 3256
rect 383568 3204 383620 3256
rect 390560 3204 390612 3256
rect 391848 3204 391900 3256
rect 128176 3068 128228 3120
rect 131396 3068 131448 3120
rect 129372 3000 129424 3052
rect 131488 3000 131540 3052
rect 136180 2932 136232 2984
rect 141240 2932 141292 2984
rect 432052 1776 432104 1828
rect 433248 1776 433300 1828
<< metal2 >>
rect 6932 703582 7972 703610
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3330 566944 3386 566953
rect 3330 566879 3386 566888
rect 3344 565894 3372 566879
rect 3332 565888 3384 565894
rect 3332 565830 3384 565836
rect 2778 553888 2834 553897
rect 2778 553823 2780 553832
rect 2832 553823 2834 553832
rect 2780 553794 2832 553800
rect 3330 514856 3386 514865
rect 3330 514791 3332 514800
rect 3384 514791 3386 514800
rect 3332 514762 3384 514768
rect 2778 501800 2834 501809
rect 2778 501735 2834 501744
rect 2792 501090 2820 501735
rect 2780 501084 2832 501090
rect 2780 501026 2832 501032
rect 2778 462632 2834 462641
rect 2778 462567 2780 462576
rect 2832 462567 2834 462576
rect 2780 462538 2832 462544
rect 2778 449576 2834 449585
rect 2778 449511 2834 449520
rect 2792 448866 2820 449511
rect 2780 448860 2832 448866
rect 2780 448802 2832 448808
rect 3330 410544 3386 410553
rect 3330 410479 3386 410488
rect 3344 409970 3372 410479
rect 3332 409964 3384 409970
rect 3332 409906 3384 409912
rect 2780 397520 2832 397526
rect 2778 397488 2780 397497
rect 2832 397488 2834 397497
rect 2778 397423 2834 397432
rect 3330 358456 3386 358465
rect 3330 358391 3386 358400
rect 3344 357474 3372 358391
rect 3332 357468 3384 357474
rect 3332 357410 3384 357416
rect 2778 345400 2834 345409
rect 2778 345335 2834 345344
rect 2792 345234 2820 345335
rect 2780 345228 2832 345234
rect 2780 345170 2832 345176
rect 3330 319288 3386 319297
rect 3330 319223 3386 319232
rect 3238 306232 3294 306241
rect 3238 306167 3294 306176
rect 3252 305046 3280 306167
rect 3240 305040 3292 305046
rect 3240 304982 3292 304988
rect 3238 293176 3294 293185
rect 3238 293111 3294 293120
rect 3252 292602 3280 293111
rect 3240 292596 3292 292602
rect 3240 292538 3292 292544
rect 3238 267200 3294 267209
rect 3238 267135 3294 267144
rect 3146 254144 3202 254153
rect 3146 254079 3202 254088
rect 3160 253978 3188 254079
rect 3148 253972 3200 253978
rect 3148 253914 3200 253920
rect 3054 241088 3110 241097
rect 3054 241023 3110 241032
rect 3068 240174 3096 241023
rect 3056 240168 3108 240174
rect 3056 240110 3108 240116
rect 3146 214976 3202 214985
rect 3146 214911 3202 214920
rect 3160 213994 3188 214911
rect 3148 213988 3200 213994
rect 3148 213930 3200 213936
rect 3146 201920 3202 201929
rect 3146 201855 3202 201864
rect 3160 201550 3188 201855
rect 3148 201544 3200 201550
rect 3148 201486 3200 201492
rect 3146 188864 3202 188873
rect 3146 188799 3202 188808
rect 3160 187746 3188 188799
rect 3148 187740 3200 187746
rect 3148 187682 3200 187688
rect 3148 162920 3200 162926
rect 3146 162888 3148 162897
rect 3200 162888 3202 162897
rect 3146 162823 3202 162832
rect 3146 149832 3202 149841
rect 3146 149767 3202 149776
rect 3160 149122 3188 149767
rect 3148 149116 3200 149122
rect 3148 149058 3200 149064
rect 3252 136134 3280 267135
rect 3240 136128 3292 136134
rect 3240 136070 3292 136076
rect 3344 136066 3372 319223
rect 3436 138378 3464 684247
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3606 632088 3662 632097
rect 3606 632023 3662 632032
rect 3514 619168 3570 619177
rect 3514 619103 3570 619112
rect 3528 618322 3556 619103
rect 3516 618316 3568 618322
rect 3516 618258 3568 618264
rect 3514 606112 3570 606121
rect 3514 606047 3570 606056
rect 3424 138372 3476 138378
rect 3424 138314 3476 138320
rect 3422 136776 3478 136785
rect 3422 136711 3478 136720
rect 3436 136678 3464 136711
rect 3424 136672 3476 136678
rect 3424 136614 3476 136620
rect 3332 136060 3384 136066
rect 3332 136002 3384 136008
rect 3424 131164 3476 131170
rect 3424 131106 3476 131112
rect 3330 84688 3386 84697
rect 3330 84623 3386 84632
rect 3344 84250 3372 84623
rect 3332 84244 3384 84250
rect 3332 84186 3384 84192
rect 2872 33108 2924 33114
rect 2872 33050 2924 33056
rect 2884 32473 2912 33050
rect 2870 32464 2926 32473
rect 2870 32399 2926 32408
rect 3436 19417 3464 131106
rect 3528 74361 3556 606047
rect 3620 134706 3648 632023
rect 3698 580000 3754 580009
rect 3698 579935 3754 579944
rect 3712 136202 3740 579935
rect 4804 553852 4856 553858
rect 4804 553794 4856 553800
rect 3790 527912 3846 527921
rect 3790 527847 3846 527856
rect 3804 136338 3832 527847
rect 3882 475688 3938 475697
rect 3882 475623 3938 475632
rect 3792 136332 3844 136338
rect 3792 136274 3844 136280
rect 3896 136270 3924 475623
rect 4066 423600 4122 423609
rect 4066 423535 4122 423544
rect 3974 371376 4030 371385
rect 3974 371311 4030 371320
rect 3988 136406 4016 371311
rect 4080 231130 4108 423535
rect 4068 231124 4120 231130
rect 4068 231066 4120 231072
rect 4068 138372 4120 138378
rect 4068 138314 4120 138320
rect 3976 136400 4028 136406
rect 3976 136342 4028 136348
rect 3884 136264 3936 136270
rect 3884 136206 3936 136212
rect 3700 136196 3752 136202
rect 3700 136138 3752 136144
rect 3608 134700 3660 134706
rect 3608 134642 3660 134648
rect 4080 134638 4108 138314
rect 4068 134632 4120 134638
rect 4068 134574 4120 134580
rect 3792 133952 3844 133958
rect 3792 133894 3844 133900
rect 3608 128376 3660 128382
rect 3608 128318 3660 128324
rect 3514 74352 3570 74361
rect 3514 74287 3570 74296
rect 3516 71732 3568 71738
rect 3516 71674 3568 71680
rect 3528 71641 3556 71674
rect 3514 71632 3570 71641
rect 3514 71567 3570 71576
rect 3620 58585 3648 128318
rect 3700 127016 3752 127022
rect 3700 126958 3752 126964
rect 3712 97617 3740 126958
rect 3804 110673 3832 133894
rect 3790 110664 3846 110673
rect 3790 110599 3846 110608
rect 3698 97608 3754 97617
rect 3698 97543 3754 97552
rect 4816 75041 4844 553794
rect 4896 501084 4948 501090
rect 4896 501026 4948 501032
rect 4802 75032 4858 75041
rect 4802 74967 4858 74976
rect 4908 73953 4936 501026
rect 5080 462596 5132 462602
rect 5080 462538 5132 462544
rect 4988 448860 5040 448866
rect 4988 448802 5040 448808
rect 5000 75177 5028 448802
rect 5092 118658 5120 462538
rect 5172 397520 5224 397526
rect 5172 397462 5224 397468
rect 5080 118652 5132 118658
rect 5080 118594 5132 118600
rect 4986 75168 5042 75177
rect 4986 75103 5042 75112
rect 4894 73944 4950 73953
rect 4894 73879 4950 73888
rect 5184 73642 5212 397462
rect 5264 345228 5316 345234
rect 5264 345170 5316 345176
rect 5276 75274 5304 345170
rect 5264 75268 5316 75274
rect 5264 75210 5316 75216
rect 6932 74089 6960 703582
rect 7944 703474 7972 703582
rect 8086 703520 8198 704960
rect 23492 703582 24164 703610
rect 8128 703474 8156 703520
rect 7944 703446 8156 703474
rect 15844 670744 15896 670750
rect 15844 670686 15896 670692
rect 8944 409964 8996 409970
rect 8944 409906 8996 409912
rect 8956 120086 8984 409906
rect 10324 357468 10376 357474
rect 10324 357410 10376 357416
rect 10336 121446 10364 357410
rect 10324 121440 10376 121446
rect 10324 121382 10376 121388
rect 8944 120080 8996 120086
rect 8944 120022 8996 120028
rect 15856 111790 15884 670686
rect 19984 565888 20036 565894
rect 19984 565830 20036 565836
rect 19996 115938 20024 565830
rect 22744 253972 22796 253978
rect 22744 253914 22796 253920
rect 22756 124166 22784 253914
rect 22836 201544 22888 201550
rect 22836 201486 22888 201492
rect 22848 125594 22876 201486
rect 22836 125588 22888 125594
rect 22836 125530 22888 125536
rect 22744 124160 22796 124166
rect 22744 124102 22796 124108
rect 19984 115932 20036 115938
rect 19984 115874 20036 115880
rect 15844 111784 15896 111790
rect 15844 111726 15896 111732
rect 23492 110430 23520 703582
rect 24136 703474 24164 703582
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 24320 703474 24348 703520
rect 24136 703446 24348 703474
rect 37924 618316 37976 618322
rect 37924 618258 37976 618264
rect 24124 305040 24176 305046
rect 24124 304982 24176 304988
rect 24136 122806 24164 304982
rect 25504 149116 25556 149122
rect 25504 149058 25556 149064
rect 25516 126954 25544 149058
rect 25504 126948 25556 126954
rect 25504 126890 25556 126896
rect 24124 122800 24176 122806
rect 24124 122742 24176 122748
rect 37936 113150 37964 618258
rect 40052 136474 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 104912 703582 105308 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 703050 73016 703520
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 62672 537532 62724 537538
rect 62672 537474 62724 537480
rect 62684 533050 62712 537474
rect 61384 533044 61436 533050
rect 61384 532986 61436 532992
rect 62672 533044 62724 533050
rect 62672 532986 62724 532992
rect 42064 514820 42116 514826
rect 42064 514762 42116 514768
rect 40040 136468 40092 136474
rect 40040 136410 40092 136416
rect 42076 117298 42104 514762
rect 58624 474700 58676 474706
rect 58624 474642 58676 474648
rect 58636 466478 58664 474642
rect 55864 466472 55916 466478
rect 55864 466414 55916 466420
rect 58624 466472 58676 466478
rect 58624 466414 58676 466420
rect 55876 451926 55904 466414
rect 46204 451920 46256 451926
rect 46204 451862 46256 451868
rect 55864 451920 55916 451926
rect 55864 451862 55916 451868
rect 46216 428330 46244 451862
rect 45100 428324 45152 428330
rect 45100 428266 45152 428272
rect 46204 428324 46256 428330
rect 46204 428266 46256 428272
rect 43444 292596 43496 292602
rect 43444 292538 43496 292544
rect 42064 117292 42116 117298
rect 42064 117234 42116 117240
rect 37924 113144 37976 113150
rect 37924 113086 37976 113092
rect 23480 110424 23532 110430
rect 23480 110366 23532 110372
rect 43456 74458 43484 292538
rect 45008 274780 45060 274786
rect 45008 274722 45060 274728
rect 44824 243908 44876 243914
rect 44824 243850 44876 243856
rect 43536 240168 43588 240174
rect 43536 240110 43588 240116
rect 43444 74452 43496 74458
rect 43444 74394 43496 74400
rect 43548 74390 43576 240110
rect 44836 233238 44864 243850
rect 44916 240780 44968 240786
rect 44916 240722 44968 240728
rect 44824 233232 44876 233238
rect 44824 233174 44876 233180
rect 44928 231198 44956 240722
rect 44916 231192 44968 231198
rect 44916 231134 44968 231140
rect 45020 220862 45048 274722
rect 45008 220856 45060 220862
rect 45008 220798 45060 220804
rect 45112 208418 45140 428266
rect 61396 376650 61424 532986
rect 69480 509924 69532 509930
rect 69480 509866 69532 509872
rect 69492 504422 69520 509866
rect 61476 504416 61528 504422
rect 61476 504358 61528 504364
rect 69480 504416 69532 504422
rect 69480 504358 69532 504364
rect 61488 474706 61516 504358
rect 61476 474700 61528 474706
rect 61476 474642 61528 474648
rect 58624 376644 58676 376650
rect 58624 376586 58676 376592
rect 61384 376644 61436 376650
rect 61384 376586 61436 376592
rect 58636 346390 58664 376586
rect 69664 356720 69716 356726
rect 69664 356662 69716 356668
rect 56876 346384 56928 346390
rect 56876 346326 56928 346332
rect 58624 346384 58676 346390
rect 58624 346326 58676 346332
rect 56888 338298 56916 346326
rect 69676 339726 69704 356662
rect 68284 339720 68336 339726
rect 68284 339662 68336 339668
rect 69664 339720 69716 339726
rect 69664 339662 69716 339668
rect 55864 338292 55916 338298
rect 55864 338234 55916 338240
rect 56876 338292 56928 338298
rect 56876 338234 56928 338240
rect 55876 323406 55904 338234
rect 53104 323400 53156 323406
rect 53104 323342 53156 323348
rect 55864 323400 55916 323406
rect 55864 323342 55916 323348
rect 53116 305046 53144 323342
rect 62764 313948 62816 313954
rect 62764 313890 62816 313896
rect 51724 305040 51776 305046
rect 51724 304982 51776 304988
rect 53104 305040 53156 305046
rect 53104 304982 53156 304988
rect 49608 287632 49660 287638
rect 49608 287574 49660 287580
rect 49620 284374 49648 287574
rect 46204 284368 46256 284374
rect 46204 284310 46256 284316
rect 49608 284368 49660 284374
rect 49608 284310 49660 284316
rect 46216 274786 46244 284310
rect 46204 274780 46256 274786
rect 46204 274722 46256 274728
rect 51080 266416 51132 266422
rect 51080 266358 51132 266364
rect 50344 262880 50396 262886
rect 50344 262822 50396 262828
rect 47584 260500 47636 260506
rect 47584 260442 47636 260448
rect 47492 256760 47544 256766
rect 47492 256702 47544 256708
rect 47504 253978 47532 256702
rect 45836 253972 45888 253978
rect 45836 253914 45888 253920
rect 47492 253972 47544 253978
rect 47492 253914 47544 253920
rect 45744 243568 45796 243574
rect 45744 243510 45796 243516
rect 45652 241460 45704 241466
rect 45652 241402 45704 241408
rect 45560 241392 45612 241398
rect 45560 241334 45612 241340
rect 45376 240916 45428 240922
rect 45376 240858 45428 240864
rect 45284 240848 45336 240854
rect 45284 240790 45336 240796
rect 45192 238808 45244 238814
rect 45192 238750 45244 238756
rect 45204 232966 45232 238750
rect 45192 232960 45244 232966
rect 45192 232902 45244 232908
rect 45296 232286 45324 240790
rect 45388 232354 45416 240858
rect 45468 240100 45520 240106
rect 45468 240042 45520 240048
rect 45480 232422 45508 240042
rect 45468 232416 45520 232422
rect 45468 232358 45520 232364
rect 45376 232348 45428 232354
rect 45376 232290 45428 232296
rect 45284 232280 45336 232286
rect 45284 232222 45336 232228
rect 45100 208412 45152 208418
rect 45100 208354 45152 208360
rect 45572 170406 45600 241334
rect 45664 184890 45692 241402
rect 45756 232218 45784 243510
rect 45848 238814 45876 253914
rect 46940 249484 46992 249490
rect 46940 249426 46992 249432
rect 46952 248414 46980 249426
rect 46860 248386 46980 248414
rect 46860 243914 46888 248386
rect 46848 243908 46900 243914
rect 46848 243850 46900 243856
rect 47124 241732 47176 241738
rect 47124 241674 47176 241680
rect 47136 240174 47164 241674
rect 47596 241398 47624 260442
rect 49240 259004 49292 259010
rect 49240 258946 49292 258952
rect 49252 256766 49280 258946
rect 49240 256760 49292 256766
rect 49240 256702 49292 256708
rect 50356 252618 50384 262822
rect 50896 261248 50948 261254
rect 50896 261190 50948 261196
rect 50908 259010 50936 261190
rect 51092 260506 51120 266358
rect 51080 260500 51132 260506
rect 51080 260442 51132 260448
rect 50896 259004 50948 259010
rect 50896 258946 50948 258952
rect 48688 252612 48740 252618
rect 48688 252554 48740 252560
rect 50344 252612 50396 252618
rect 50344 252554 50396 252560
rect 47676 251864 47728 251870
rect 47676 251806 47728 251812
rect 47688 241466 47716 251806
rect 48700 249490 48728 252554
rect 48688 249484 48740 249490
rect 48688 249426 48740 249432
rect 51736 247110 51764 304982
rect 57244 301504 57296 301510
rect 57244 301446 57296 301452
rect 51816 300144 51868 300150
rect 51816 300086 51868 300092
rect 51828 287638 51856 300086
rect 57256 288386 57284 301446
rect 62776 301102 62804 313890
rect 67180 303680 67232 303686
rect 67180 303622 67232 303628
rect 61384 301096 61436 301102
rect 61384 301038 61436 301044
rect 62764 301096 62816 301102
rect 62764 301038 62816 301044
rect 55864 288380 55916 288386
rect 55864 288322 55916 288328
rect 57244 288380 57296 288386
rect 57244 288322 57296 288328
rect 51816 287632 51868 287638
rect 51816 287574 51868 287580
rect 55876 272950 55904 288322
rect 61396 280838 61424 301038
rect 66904 300212 66956 300218
rect 66904 300154 66956 300160
rect 60004 280832 60056 280838
rect 60004 280774 60056 280780
rect 61384 280832 61436 280838
rect 61384 280774 61436 280780
rect 60016 274718 60044 280774
rect 57980 274712 58032 274718
rect 57980 274654 58032 274660
rect 60004 274712 60056 274718
rect 60004 274654 60056 274660
rect 54484 272944 54536 272950
rect 54484 272886 54536 272892
rect 55864 272944 55916 272950
rect 55864 272886 55916 272892
rect 52368 269136 52420 269142
rect 52368 269078 52420 269084
rect 52380 261254 52408 269078
rect 54496 266422 54524 272886
rect 57992 270586 58020 274654
rect 57900 270558 58020 270586
rect 57900 269142 57928 270558
rect 65524 270496 65576 270502
rect 65524 270438 65576 270444
rect 57888 269136 57940 269142
rect 57888 269078 57940 269084
rect 63500 266552 63552 266558
rect 63500 266494 63552 266500
rect 54484 266416 54536 266422
rect 54484 266358 54536 266364
rect 63512 262886 63540 266494
rect 63500 262880 63552 262886
rect 63500 262822 63552 262828
rect 52368 261248 52420 261254
rect 52368 261190 52420 261196
rect 65536 259486 65564 270438
rect 66916 266558 66944 300154
rect 67192 300150 67220 303622
rect 68296 300218 68324 339662
rect 69664 311160 69716 311166
rect 69664 311102 69716 311108
rect 69676 303686 69704 311102
rect 69664 303680 69716 303686
rect 69664 303622 69716 303628
rect 68284 300212 68336 300218
rect 68284 300154 68336 300160
rect 67180 300144 67232 300150
rect 67180 300086 67232 300092
rect 69480 279744 69532 279750
rect 69480 279686 69532 279692
rect 69492 270570 69520 279686
rect 69480 270564 69532 270570
rect 69480 270506 69532 270512
rect 66904 266552 66956 266558
rect 66904 266494 66956 266500
rect 65524 259480 65576 259486
rect 65524 259422 65576 259428
rect 60648 259412 60700 259418
rect 60648 259354 60700 259360
rect 60660 251938 60688 259354
rect 57980 251932 58032 251938
rect 57980 251874 58032 251880
rect 60648 251932 60700 251938
rect 60648 251874 60700 251880
rect 57992 249082 58020 251874
rect 71792 251870 71820 702986
rect 89180 702434 89208 703520
rect 88352 702406 89208 702434
rect 83464 537600 83516 537606
rect 83464 537542 83516 537548
rect 83476 512990 83504 537542
rect 80060 512984 80112 512990
rect 80060 512926 80112 512932
rect 83464 512984 83516 512990
rect 83464 512926 83516 512932
rect 80072 509930 80100 512926
rect 80060 509924 80112 509930
rect 80060 509866 80112 509872
rect 87604 336796 87656 336802
rect 87604 336738 87656 336744
rect 87616 323610 87644 336738
rect 81716 323604 81768 323610
rect 81716 323546 81768 323552
rect 87604 323604 87656 323610
rect 87604 323546 87656 323552
rect 81728 316810 81756 323546
rect 88352 318782 88380 702406
rect 94504 543040 94556 543046
rect 94504 542982 94556 542988
rect 94516 537606 94544 542982
rect 94504 537600 94556 537606
rect 94504 537542 94556 537548
rect 102784 412684 102836 412690
rect 102784 412626 102836 412632
rect 102796 392018 102824 412626
rect 101404 392012 101456 392018
rect 101404 391954 101456 391960
rect 102784 392012 102836 392018
rect 102784 391954 102836 391960
rect 101416 368558 101444 391954
rect 101404 368552 101456 368558
rect 101404 368494 101456 368500
rect 98644 368484 98696 368490
rect 98644 368426 98696 368432
rect 94504 348900 94556 348906
rect 94504 348842 94556 348848
rect 94516 336802 94544 348842
rect 98656 338842 98684 368426
rect 99012 354000 99064 354006
rect 99012 353942 99064 353948
rect 99024 348906 99052 353942
rect 99012 348900 99064 348906
rect 99012 348842 99064 348848
rect 97264 338836 97316 338842
rect 97264 338778 97316 338784
rect 98644 338836 98696 338842
rect 98644 338778 98696 338784
rect 94504 336796 94556 336802
rect 94504 336738 94556 336744
rect 97276 329118 97304 338778
rect 95884 329112 95936 329118
rect 95884 329054 95936 329060
rect 97264 329112 97316 329118
rect 97264 329054 97316 329060
rect 95896 321774 95924 329054
rect 94780 321768 94832 321774
rect 94780 321710 94832 321716
rect 95884 321768 95936 321774
rect 95884 321710 95936 321716
rect 94792 319802 94820 321710
rect 91100 319796 91152 319802
rect 91100 319738 91152 319744
rect 94780 319796 94832 319802
rect 94780 319738 94832 319744
rect 85580 318776 85632 318782
rect 85580 318718 85632 318724
rect 88340 318776 88392 318782
rect 88340 318718 88392 318724
rect 79232 316804 79284 316810
rect 79232 316746 79284 316752
rect 81716 316804 81768 316810
rect 81716 316746 81768 316752
rect 79244 311166 79272 316746
rect 85592 313410 85620 318718
rect 91112 317490 91140 319738
rect 91100 317484 91152 317490
rect 91100 317426 91152 317432
rect 88340 317416 88392 317422
rect 88340 317358 88392 317364
rect 79324 313404 79376 313410
rect 79324 313346 79376 313352
rect 85580 313404 85632 313410
rect 85580 313346 85632 313352
rect 79232 311160 79284 311166
rect 79232 311102 79284 311108
rect 79336 301510 79364 313346
rect 88352 311930 88380 317358
rect 104912 313954 104940 703582
rect 105280 703474 105308 703582
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 136652 703582 137692 703610
rect 105464 703474 105492 703520
rect 105280 703446 105492 703474
rect 133696 646876 133748 646882
rect 133696 646818 133748 646824
rect 133708 644502 133736 646818
rect 131764 644496 131816 644502
rect 131764 644438 131816 644444
rect 133696 644496 133748 644502
rect 133696 644438 133748 644444
rect 131776 632126 131804 644438
rect 128360 632120 128412 632126
rect 128360 632062 128412 632068
rect 131764 632120 131816 632126
rect 131764 632062 131816 632068
rect 128372 629746 128400 632062
rect 127624 629740 127676 629746
rect 127624 629682 127676 629688
rect 128360 629740 128412 629746
rect 128360 629682 128412 629688
rect 127636 623830 127664 629682
rect 127624 623824 127676 623830
rect 127624 623766 127676 623772
rect 124220 623756 124272 623762
rect 124220 623698 124272 623704
rect 124232 621042 124260 623698
rect 123484 621036 123536 621042
rect 123484 620978 123536 620984
rect 124220 621036 124272 621042
rect 124220 620978 124272 620984
rect 123496 600370 123524 620978
rect 123484 600364 123536 600370
rect 123484 600306 123536 600312
rect 120724 600296 120776 600302
rect 120724 600238 120776 600244
rect 120736 591326 120764 600238
rect 112444 591320 112496 591326
rect 112444 591262 112496 591268
rect 120724 591320 120776 591326
rect 120724 591262 120776 591268
rect 112456 565894 112484 591262
rect 111064 565888 111116 565894
rect 111064 565830 111116 565836
rect 112444 565888 112496 565894
rect 112444 565830 112496 565836
rect 111076 551342 111104 565830
rect 127624 560992 127676 560998
rect 127624 560934 127676 560940
rect 127636 554062 127664 560934
rect 117228 554056 117280 554062
rect 117228 553998 117280 554004
rect 127624 554056 127676 554062
rect 127624 553998 127676 554004
rect 109684 551336 109736 551342
rect 109684 551278 109736 551284
rect 111064 551336 111116 551342
rect 111064 551278 111116 551284
rect 104992 549908 105044 549914
rect 104992 549850 105044 549856
rect 105004 543046 105032 549850
rect 104992 543040 105044 543046
rect 104992 542982 105044 542988
rect 109696 516186 109724 551278
rect 117240 549914 117268 553998
rect 117228 549908 117280 549914
rect 117228 549850 117280 549856
rect 109684 516180 109736 516186
rect 109684 516122 109736 516128
rect 105544 516112 105596 516118
rect 105544 516054 105596 516060
rect 105556 412690 105584 516054
rect 136652 508570 136680 703582
rect 137664 703474 137692 703582
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 234632 703582 235028 703610
rect 137848 703474 137876 703520
rect 137664 703446 137876 703474
rect 154132 699718 154160 703520
rect 170324 702434 170352 703520
rect 202800 703050 202828 703520
rect 201500 703044 201552 703050
rect 201500 702986 201552 702992
rect 202788 703044 202840 703050
rect 202788 702986 202840 702992
rect 169772 702406 170352 702434
rect 153016 699712 153068 699718
rect 153016 699654 153068 699660
rect 154120 699712 154172 699718
rect 154120 699654 154172 699660
rect 153028 696998 153056 699654
rect 153016 696992 153068 696998
rect 153016 696934 153068 696940
rect 146944 696924 146996 696930
rect 146944 696866 146996 696872
rect 146956 688702 146984 696866
rect 145656 688696 145708 688702
rect 145656 688638 145708 688644
rect 146944 688696 146996 688702
rect 146944 688638 146996 688644
rect 145668 684010 145696 688638
rect 144184 684004 144236 684010
rect 144184 683946 144236 683952
rect 145656 684004 145708 684010
rect 145656 683946 145708 683952
rect 144196 670750 144224 683946
rect 144184 670744 144236 670750
rect 144184 670686 144236 670692
rect 140320 670676 140372 670682
rect 140320 670618 140372 670624
rect 140332 667962 140360 670618
rect 138664 667956 138716 667962
rect 138664 667898 138716 667904
rect 140320 667956 140372 667962
rect 140320 667898 140372 667904
rect 138676 651438 138704 667898
rect 136732 651432 136784 651438
rect 136732 651374 136784 651380
rect 138664 651432 138716 651438
rect 138664 651374 138716 651380
rect 136744 646882 136772 651374
rect 136732 646876 136784 646882
rect 136732 646818 136784 646824
rect 155224 632732 155276 632738
rect 155224 632674 155276 632680
rect 155236 572014 155264 632674
rect 169024 616140 169076 616146
rect 169024 616082 169076 616088
rect 144184 572008 144236 572014
rect 144184 571950 144236 571956
rect 155224 572008 155276 572014
rect 155224 571950 155276 571956
rect 144196 563106 144224 571950
rect 140780 563100 140832 563106
rect 140780 563042 140832 563048
rect 144184 563100 144236 563106
rect 144184 563042 144236 563048
rect 140792 560998 140820 563042
rect 140780 560992 140832 560998
rect 140780 560934 140832 560940
rect 117964 508564 118016 508570
rect 117964 508506 118016 508512
rect 136640 508564 136692 508570
rect 136640 508506 136692 508512
rect 117976 487218 118004 508506
rect 169036 498846 169064 616082
rect 169772 537538 169800 702406
rect 201512 687954 201540 702986
rect 218992 699718 219020 703520
rect 218980 699712 219032 699718
rect 218980 699654 219032 699660
rect 215208 699644 215260 699650
rect 215208 699586 215260 699592
rect 215220 693666 215248 699586
rect 211804 693660 211856 693666
rect 211804 693602 211856 693608
rect 215208 693660 215260 693666
rect 215208 693602 215260 693608
rect 191104 687948 191156 687954
rect 191104 687890 191156 687896
rect 201500 687948 201552 687954
rect 201500 687890 201552 687896
rect 191116 680610 191144 687890
rect 187976 680604 188028 680610
rect 187976 680546 188028 680552
rect 191104 680604 191156 680610
rect 191104 680546 191156 680552
rect 187988 677618 188016 680546
rect 185584 677612 185636 677618
rect 185584 677554 185636 677560
rect 187976 677612 188028 677618
rect 187976 677554 188028 677560
rect 178040 650684 178092 650690
rect 178040 650626 178092 650632
rect 178052 647902 178080 650626
rect 170404 647896 170456 647902
rect 170404 647838 170456 647844
rect 178040 647896 178092 647902
rect 178040 647838 178092 647844
rect 170416 632738 170444 647838
rect 185596 640354 185624 677554
rect 204904 667208 204956 667214
rect 204904 667150 204956 667156
rect 204916 664494 204944 667150
rect 211816 665174 211844 693602
rect 234632 693462 234660 703582
rect 235000 703474 235028 703582
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299492 703582 299980 703610
rect 235184 703474 235212 703520
rect 235000 703446 235212 703474
rect 267660 699718 267688 703520
rect 283852 699718 283880 703520
rect 267648 699712 267700 699718
rect 267648 699654 267700 699660
rect 282184 699712 282236 699718
rect 282184 699654 282236 699660
rect 283840 699712 283892 699718
rect 283840 699654 283892 699660
rect 262864 699644 262916 699650
rect 262864 699586 262916 699592
rect 226984 693456 227036 693462
rect 226984 693398 227036 693404
rect 234620 693456 234672 693462
rect 234620 693398 234672 693404
rect 226996 676802 227024 693398
rect 221464 676796 221516 676802
rect 221464 676738 221516 676744
rect 226984 676796 227036 676802
rect 226984 676738 227036 676744
rect 221476 672110 221504 676738
rect 262876 675034 262904 699586
rect 282196 679046 282224 699654
rect 299492 681222 299520 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 412652 703582 413508 703610
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 332520 699718 332548 703520
rect 348804 699854 348832 703520
rect 348792 699848 348844 699854
rect 348792 699790 348844 699796
rect 351184 699848 351236 699854
rect 351184 699790 351236 699796
rect 332508 699712 332560 699718
rect 332508 699654 332560 699660
rect 336004 699712 336056 699718
rect 336004 699654 336056 699660
rect 336016 684486 336044 699654
rect 351196 690674 351224 699790
rect 364996 698154 365024 703520
rect 364984 698148 365036 698154
rect 364984 698090 365036 698096
rect 369124 698148 369176 698154
rect 369124 698090 369176 698096
rect 351184 690668 351236 690674
rect 351184 690610 351236 690616
rect 359464 690668 359516 690674
rect 359464 690610 359516 690616
rect 336004 684480 336056 684486
rect 336004 684422 336056 684428
rect 341248 684480 341300 684486
rect 341248 684422 341300 684428
rect 299480 681216 299532 681222
rect 299480 681158 299532 681164
rect 305000 681216 305052 681222
rect 305000 681158 305052 681164
rect 280896 679040 280948 679046
rect 280896 678982 280948 678988
rect 282184 679040 282236 679046
rect 282184 678982 282236 678988
rect 280908 677074 280936 678982
rect 279424 677068 279476 677074
rect 279424 677010 279476 677016
rect 280896 677068 280948 677074
rect 280896 677010 280948 677016
rect 259460 675028 259512 675034
rect 259460 674970 259512 674976
rect 262864 675028 262916 675034
rect 262864 674970 262916 674976
rect 259472 672110 259500 674970
rect 215300 672104 215352 672110
rect 215300 672046 215352 672052
rect 221464 672104 221516 672110
rect 221464 672046 221516 672052
rect 259460 672104 259512 672110
rect 259460 672046 259512 672052
rect 215312 667214 215340 672046
rect 255688 672036 255740 672042
rect 255688 671978 255740 671984
rect 255700 669390 255728 671978
rect 253204 669384 253256 669390
rect 253204 669326 253256 669332
rect 255688 669384 255740 669390
rect 255688 669326 255740 669332
rect 215300 667208 215352 667214
rect 215300 667150 215352 667156
rect 210424 665168 210476 665174
rect 210424 665110 210476 665116
rect 211804 665168 211856 665174
rect 211804 665110 211856 665116
rect 197268 664488 197320 664494
rect 197268 664430 197320 664436
rect 204904 664488 204956 664494
rect 204904 664430 204956 664436
rect 197280 661094 197308 664430
rect 191104 661088 191156 661094
rect 191104 661030 191156 661036
rect 197268 661088 197320 661094
rect 197268 661030 197320 661036
rect 191116 650690 191144 661030
rect 191104 650684 191156 650690
rect 191104 650626 191156 650632
rect 181444 640348 181496 640354
rect 181444 640290 181496 640296
rect 185584 640348 185636 640354
rect 185584 640290 185636 640296
rect 170404 632732 170456 632738
rect 170404 632674 170456 632680
rect 181456 622742 181484 640290
rect 210436 636274 210464 665110
rect 207664 636268 207716 636274
rect 207664 636210 207716 636216
rect 210424 636268 210476 636274
rect 210424 636210 210476 636216
rect 207676 625258 207704 636210
rect 204904 625252 204956 625258
rect 204904 625194 204956 625200
rect 207664 625252 207716 625258
rect 207664 625194 207716 625200
rect 175924 622736 175976 622742
rect 175924 622678 175976 622684
rect 181444 622736 181496 622742
rect 181444 622678 181496 622684
rect 175936 616146 175964 622678
rect 175924 616140 175976 616146
rect 175924 616082 175976 616088
rect 204916 609278 204944 625194
rect 203524 609272 203576 609278
rect 203524 609214 203576 609220
rect 204904 609272 204956 609278
rect 204904 609214 204956 609220
rect 203536 558890 203564 609214
rect 253216 601730 253244 669326
rect 279436 662454 279464 677010
rect 305012 675646 305040 681158
rect 341260 679182 341288 684422
rect 359476 679318 359504 690610
rect 369136 690402 369164 698090
rect 369124 690396 369176 690402
rect 369124 690338 369176 690344
rect 371240 690396 371292 690402
rect 371240 690338 371292 690344
rect 371252 687954 371280 690338
rect 371240 687948 371292 687954
rect 371240 687890 371292 687896
rect 377404 687948 377456 687954
rect 377404 687890 377456 687896
rect 359464 679312 359516 679318
rect 359464 679254 359516 679260
rect 362224 679312 362276 679318
rect 362224 679254 362276 679260
rect 341248 679176 341300 679182
rect 341248 679118 341300 679124
rect 344284 679176 344336 679182
rect 344284 679118 344336 679124
rect 305000 675640 305052 675646
rect 305000 675582 305052 675588
rect 307760 675640 307812 675646
rect 307760 675582 307812 675588
rect 307772 672790 307800 675582
rect 307760 672784 307812 672790
rect 307760 672726 307812 672732
rect 319904 672784 319956 672790
rect 319904 672726 319956 672732
rect 319916 665174 319944 672726
rect 344296 669322 344324 679118
rect 362236 670002 362264 679254
rect 377416 678978 377444 687890
rect 377404 678972 377456 678978
rect 377404 678914 377456 678920
rect 385684 678972 385736 678978
rect 385684 678914 385736 678920
rect 362224 669996 362276 670002
rect 362224 669938 362276 669944
rect 383936 669996 383988 670002
rect 383936 669938 383988 669944
rect 344284 669316 344336 669322
rect 344284 669258 344336 669264
rect 346676 669316 346728 669322
rect 346676 669258 346728 669264
rect 319904 665168 319956 665174
rect 319904 665110 319956 665116
rect 324964 665168 325016 665174
rect 324964 665110 325016 665116
rect 277492 662448 277544 662454
rect 277492 662390 277544 662396
rect 279424 662448 279476 662454
rect 279424 662390 279476 662396
rect 277504 660618 277532 662390
rect 276664 660612 276716 660618
rect 276664 660554 276716 660560
rect 277492 660612 277544 660618
rect 277492 660554 277544 660560
rect 276676 640354 276704 660554
rect 276664 640348 276716 640354
rect 276664 640290 276716 640296
rect 272524 640280 272576 640286
rect 272524 640222 272576 640228
rect 272536 614174 272564 640222
rect 324976 635526 325004 665110
rect 346688 664494 346716 669258
rect 383948 665854 383976 669938
rect 383936 665848 383988 665854
rect 383936 665790 383988 665796
rect 385696 665174 385724 678914
rect 395344 665848 395396 665854
rect 395344 665790 395396 665796
rect 385684 665168 385736 665174
rect 385684 665110 385736 665116
rect 389824 665168 389876 665174
rect 389824 665110 389876 665116
rect 346676 664488 346728 664494
rect 346676 664430 346728 664436
rect 364984 664488 365036 664494
rect 364984 664430 365036 664436
rect 324964 635520 325016 635526
rect 324964 635462 325016 635468
rect 329196 635520 329248 635526
rect 329196 635462 329248 635468
rect 329208 629270 329236 635462
rect 329196 629264 329248 629270
rect 329196 629206 329248 629212
rect 331864 629264 331916 629270
rect 331864 629206 331916 629212
rect 270500 614168 270552 614174
rect 270500 614110 270552 614116
rect 272524 614168 272576 614174
rect 272524 614110 272576 614116
rect 270512 609278 270540 614110
rect 331876 611318 331904 629206
rect 364996 626550 365024 664430
rect 389836 656878 389864 665110
rect 389824 656872 389876 656878
rect 389824 656814 389876 656820
rect 392584 656872 392636 656878
rect 392584 656814 392636 656820
rect 392596 646202 392624 656814
rect 392584 646196 392636 646202
rect 392584 646138 392636 646144
rect 364984 626544 365036 626550
rect 364984 626486 365036 626492
rect 369124 626544 369176 626550
rect 369124 626486 369176 626492
rect 331864 611312 331916 611318
rect 331864 611254 331916 611260
rect 337384 611312 337436 611318
rect 337384 611254 337436 611260
rect 263600 609272 263652 609278
rect 263600 609214 263652 609220
rect 270500 609272 270552 609278
rect 270500 609214 270552 609220
rect 263612 606626 263640 609214
rect 262864 606620 262916 606626
rect 262864 606562 262916 606568
rect 263600 606620 263652 606626
rect 263600 606562 263652 606568
rect 251916 601724 251968 601730
rect 251916 601666 251968 601672
rect 253204 601724 253256 601730
rect 253204 601666 253256 601672
rect 251928 596970 251956 601666
rect 262876 598670 262904 606562
rect 261484 598664 261536 598670
rect 261484 598606 261536 598612
rect 262864 598664 262916 598670
rect 262864 598606 262916 598612
rect 250444 596964 250496 596970
rect 250444 596906 250496 596912
rect 251916 596964 251968 596970
rect 251916 596906 251968 596912
rect 250456 586566 250484 596906
rect 250444 586560 250496 586566
rect 250444 586502 250496 586508
rect 246304 586492 246356 586498
rect 246304 586434 246356 586440
rect 246316 564466 246344 586434
rect 243544 564460 243596 564466
rect 243544 564402 243596 564408
rect 246304 564460 246356 564466
rect 246304 564402 246356 564408
rect 202144 558884 202196 558890
rect 202144 558826 202196 558832
rect 203524 558884 203576 558890
rect 203524 558826 203576 558832
rect 169760 537532 169812 537538
rect 169760 537474 169812 537480
rect 202156 502994 202184 558826
rect 243556 520334 243584 564402
rect 261496 563106 261524 598606
rect 337396 592278 337424 611254
rect 337384 592272 337436 592278
rect 337384 592214 337436 592220
rect 339500 592272 339552 592278
rect 339500 592214 339552 592220
rect 339512 590646 339540 592214
rect 339500 590640 339552 590646
rect 339500 590582 339552 590588
rect 343640 590640 343692 590646
rect 343640 590582 343692 590588
rect 343652 587654 343680 590582
rect 343640 587648 343692 587654
rect 343640 587590 343692 587596
rect 347044 587648 347096 587654
rect 347044 587590 347096 587596
rect 260104 563100 260156 563106
rect 260104 563042 260156 563048
rect 261484 563100 261536 563106
rect 261484 563042 261536 563048
rect 260116 528630 260144 563042
rect 347056 562358 347084 587590
rect 369136 582282 369164 626486
rect 369124 582276 369176 582282
rect 369124 582218 369176 582224
rect 373264 582276 373316 582282
rect 373264 582218 373316 582224
rect 373276 563038 373304 582218
rect 373264 563032 373316 563038
rect 373264 562974 373316 562980
rect 376668 563032 376720 563038
rect 376668 562974 376720 562980
rect 347044 562352 347096 562358
rect 347044 562294 347096 562300
rect 349804 562352 349856 562358
rect 349804 562294 349856 562300
rect 349816 555490 349844 562294
rect 376680 559570 376708 562974
rect 376668 559564 376720 559570
rect 376668 559506 376720 559512
rect 383660 559564 383712 559570
rect 383660 559506 383712 559512
rect 383672 556782 383700 559506
rect 383660 556776 383712 556782
rect 383660 556718 383712 556724
rect 389824 556776 389876 556782
rect 389824 556718 389876 556724
rect 349804 555484 349856 555490
rect 349804 555426 349856 555432
rect 368388 555484 368440 555490
rect 368388 555426 368440 555432
rect 368400 549914 368428 555426
rect 368388 549908 368440 549914
rect 368388 549850 368440 549856
rect 382924 549908 382976 549914
rect 382924 549850 382976 549856
rect 257068 528624 257120 528630
rect 257068 528566 257120 528572
rect 260104 528624 260156 528630
rect 260104 528566 260156 528572
rect 257080 522170 257108 528566
rect 382936 528086 382964 549850
rect 389836 538014 389864 556718
rect 389824 538008 389876 538014
rect 389824 537950 389876 537956
rect 395160 538008 395212 538014
rect 395160 537950 395212 537956
rect 395172 534138 395200 537950
rect 395160 534132 395212 534138
rect 395160 534074 395212 534080
rect 382924 528080 382976 528086
rect 382924 528022 382976 528028
rect 386328 528080 386380 528086
rect 386328 528022 386380 528028
rect 386340 522986 386368 528022
rect 386328 522980 386380 522986
rect 386328 522922 386380 522928
rect 391204 522980 391256 522986
rect 391204 522922 391256 522928
rect 255964 522164 256016 522170
rect 255964 522106 256016 522112
rect 257068 522164 257120 522170
rect 257068 522106 257120 522112
rect 243544 520328 243596 520334
rect 243544 520270 243596 520276
rect 239404 520260 239456 520266
rect 239404 520202 239456 520208
rect 200764 502988 200816 502994
rect 200764 502930 200816 502936
rect 202144 502988 202196 502994
rect 202144 502930 202196 502936
rect 158720 498840 158772 498846
rect 158720 498782 158772 498788
rect 169024 498840 169076 498846
rect 169024 498782 169076 498788
rect 158732 490618 158760 498782
rect 150440 490612 150492 490618
rect 150440 490554 150492 490560
rect 158720 490612 158772 490618
rect 158720 490554 158772 490560
rect 150452 487218 150480 490554
rect 116584 487212 116636 487218
rect 116584 487154 116636 487160
rect 117964 487212 118016 487218
rect 117964 487154 118016 487160
rect 146024 487212 146076 487218
rect 146024 487154 146076 487160
rect 150440 487212 150492 487218
rect 150440 487154 150492 487160
rect 116596 473006 116624 487154
rect 146036 484362 146064 487154
rect 142804 484356 142856 484362
rect 142804 484298 142856 484304
rect 146024 484356 146076 484362
rect 146024 484298 146076 484304
rect 142816 479534 142844 484298
rect 135168 479528 135220 479534
rect 135168 479470 135220 479476
rect 142804 479528 142856 479534
rect 142804 479470 142856 479476
rect 135180 476338 135208 479470
rect 129740 476332 129792 476338
rect 129740 476274 129792 476280
rect 135168 476332 135220 476338
rect 135168 476274 135220 476280
rect 115204 473000 115256 473006
rect 115204 472942 115256 472948
rect 116584 473000 116636 473006
rect 116584 472942 116636 472948
rect 111064 427100 111116 427106
rect 111064 427042 111116 427048
rect 105544 412684 105596 412690
rect 105544 412626 105596 412632
rect 111076 390590 111104 427042
rect 108304 390584 108356 390590
rect 108304 390526 108356 390532
rect 111064 390584 111116 390590
rect 111064 390526 111116 390532
rect 108316 354006 108344 390526
rect 115216 356726 115244 472942
rect 129752 471306 129780 476274
rect 200776 472054 200804 502930
rect 239416 486538 239444 520202
rect 255976 511970 256004 522106
rect 253204 511964 253256 511970
rect 253204 511906 253256 511912
rect 255964 511964 256016 511970
rect 255964 511906 256016 511912
rect 253216 494086 253244 511906
rect 391216 498438 391244 522922
rect 391204 498432 391256 498438
rect 391204 498374 391256 498380
rect 393964 498432 394016 498438
rect 393964 498374 394016 498380
rect 253204 494080 253256 494086
rect 253204 494022 253256 494028
rect 250444 494012 250496 494018
rect 250444 493954 250496 493960
rect 237380 486532 237432 486538
rect 237380 486474 237432 486480
rect 239404 486532 239456 486538
rect 239404 486474 239456 486480
rect 237392 482594 237420 486474
rect 236644 482588 236696 482594
rect 236644 482530 236696 482536
rect 237380 482588 237432 482594
rect 237380 482530 237432 482536
rect 199384 472048 199436 472054
rect 199384 471990 199436 471996
rect 200764 472048 200816 472054
rect 200764 471990 200816 471996
rect 120724 471300 120776 471306
rect 120724 471242 120776 471248
rect 129740 471300 129792 471306
rect 129740 471242 129792 471248
rect 120736 449954 120764 471242
rect 199396 469266 199424 471990
rect 198004 469260 198056 469266
rect 198004 469202 198056 469208
rect 199384 469260 199436 469266
rect 199384 469202 199436 469208
rect 198016 456822 198044 469202
rect 198004 456816 198056 456822
rect 198004 456758 198056 456764
rect 193864 456748 193916 456754
rect 193864 456690 193916 456696
rect 117964 449948 118016 449954
rect 117964 449890 118016 449896
rect 120724 449948 120776 449954
rect 120724 449890 120776 449896
rect 117976 427106 118004 449890
rect 117964 427100 118016 427106
rect 117964 427042 118016 427048
rect 193876 425746 193904 456690
rect 192484 425740 192536 425746
rect 192484 425682 192536 425688
rect 193864 425740 193916 425746
rect 193864 425682 193916 425688
rect 192496 392018 192524 425682
rect 236656 394670 236684 482530
rect 250456 478922 250484 493954
rect 249432 478916 249484 478922
rect 249432 478858 249484 478864
rect 250444 478916 250496 478922
rect 250444 478858 250496 478864
rect 249444 474434 249472 478858
rect 393976 475454 394004 498374
rect 393964 475448 394016 475454
rect 393964 475390 394016 475396
rect 247684 474428 247736 474434
rect 247684 474370 247736 474376
rect 249432 474428 249484 474434
rect 249432 474370 249484 474376
rect 247696 419558 247724 474370
rect 247684 419552 247736 419558
rect 247684 419494 247736 419500
rect 244924 419484 244976 419490
rect 244924 419426 244976 419432
rect 244936 404326 244964 419426
rect 243544 404320 243596 404326
rect 243544 404262 243596 404268
rect 244924 404320 244976 404326
rect 244924 404262 244976 404268
rect 235264 394664 235316 394670
rect 235264 394606 235316 394612
rect 236644 394664 236696 394670
rect 236644 394606 236696 394612
rect 189724 392012 189776 392018
rect 189724 391954 189776 391960
rect 192484 392012 192536 392018
rect 192484 391954 192536 391960
rect 189736 369918 189764 391954
rect 188436 369912 188488 369918
rect 188436 369854 188488 369860
rect 189724 369912 189776 369918
rect 189724 369854 189776 369860
rect 188448 365566 188476 369854
rect 186964 365560 187016 365566
rect 186964 365502 187016 365508
rect 188436 365560 188488 365566
rect 188436 365502 188488 365508
rect 115204 356720 115256 356726
rect 115204 356662 115256 356668
rect 108304 354000 108356 354006
rect 108304 353942 108356 353948
rect 186976 353326 187004 365502
rect 235276 360262 235304 394606
rect 243556 371278 243584 404262
rect 239404 371272 239456 371278
rect 239404 371214 239456 371220
rect 243544 371272 243596 371278
rect 243544 371214 243596 371220
rect 232504 360256 232556 360262
rect 232504 360198 232556 360204
rect 235264 360256 235316 360262
rect 235264 360198 235316 360204
rect 185584 353320 185636 353326
rect 185584 353262 185636 353268
rect 186964 353320 187016 353326
rect 186964 353262 187016 353268
rect 185596 320822 185624 353262
rect 232516 348838 232544 360198
rect 239416 352102 239444 371214
rect 235264 352096 235316 352102
rect 235264 352038 235316 352044
rect 239404 352096 239456 352102
rect 239404 352038 239456 352044
rect 229744 348832 229796 348838
rect 229744 348774 229796 348780
rect 232504 348832 232556 348838
rect 232504 348774 232556 348780
rect 229756 335374 229784 348774
rect 235276 342310 235304 352038
rect 233976 342304 234028 342310
rect 233976 342246 234028 342252
rect 235264 342304 235316 342310
rect 235264 342246 235316 342252
rect 233988 340066 234016 342246
rect 232504 340060 232556 340066
rect 232504 340002 232556 340008
rect 233976 340060 234028 340066
rect 233976 340002 234028 340008
rect 229744 335368 229796 335374
rect 229744 335310 229796 335316
rect 225328 335300 225380 335306
rect 225328 335242 225380 335248
rect 225340 329050 225368 335242
rect 232516 334014 232544 340002
rect 231216 334008 231268 334014
rect 231216 333950 231268 333956
rect 232504 334008 232556 334014
rect 232504 333950 232556 333956
rect 224224 329044 224276 329050
rect 224224 328986 224276 328992
rect 225328 329044 225380 329050
rect 225328 328986 225380 328992
rect 224236 322998 224264 328986
rect 231228 326330 231256 333950
rect 229836 326324 229888 326330
rect 229836 326266 229888 326272
rect 231216 326324 231268 326330
rect 231216 326266 231268 326272
rect 229848 323610 229876 326266
rect 227720 323604 227772 323610
rect 227720 323546 227772 323552
rect 229836 323604 229888 323610
rect 229836 323546 229888 323552
rect 221464 322992 221516 322998
rect 221464 322934 221516 322940
rect 224224 322992 224276 322998
rect 224224 322934 224276 322940
rect 182456 320816 182508 320822
rect 182456 320758 182508 320764
rect 185584 320816 185636 320822
rect 185584 320758 185636 320764
rect 182468 318714 182496 320758
rect 180800 318708 180852 318714
rect 180800 318650 180852 318656
rect 182456 318708 182508 318714
rect 182456 318650 182508 318656
rect 104900 313948 104952 313954
rect 104900 313890 104952 313896
rect 180812 313682 180840 318650
rect 178684 313676 178736 313682
rect 178684 313618 178736 313624
rect 180800 313676 180852 313682
rect 180800 313618 180852 313624
rect 88260 311902 88380 311930
rect 88260 309466 88288 311902
rect 85396 309460 85448 309466
rect 85396 309402 85448 309408
rect 88248 309460 88300 309466
rect 88248 309402 88300 309408
rect 85408 307834 85436 309402
rect 81348 307828 81400 307834
rect 81348 307770 81400 307776
rect 85396 307828 85448 307834
rect 85396 307770 85448 307776
rect 79324 301504 79376 301510
rect 79324 301446 79376 301452
rect 81360 300354 81388 307770
rect 79324 300348 79376 300354
rect 79324 300290 79376 300296
rect 81348 300348 81400 300354
rect 81348 300290 81400 300296
rect 79336 292602 79364 300290
rect 76564 292596 76616 292602
rect 76564 292538 76616 292544
rect 79324 292596 79376 292602
rect 79324 292538 79376 292544
rect 76576 281994 76604 292538
rect 72056 281988 72108 281994
rect 72056 281930 72108 281936
rect 76564 281988 76616 281994
rect 76564 281930 76616 281936
rect 72068 279750 72096 281930
rect 72056 279744 72108 279750
rect 72056 279686 72108 279692
rect 178696 276078 178724 313618
rect 221476 313342 221504 322934
rect 227732 318306 227760 323546
rect 223120 318300 223172 318306
rect 223120 318242 223172 318248
rect 227720 318300 227772 318306
rect 227720 318242 227772 318248
rect 220084 313336 220136 313342
rect 220084 313278 220136 313284
rect 221464 313336 221516 313342
rect 221464 313278 221516 313284
rect 218060 292596 218112 292602
rect 218060 292538 218112 292544
rect 218072 289882 218100 292538
rect 215944 289876 215996 289882
rect 215944 289818 215996 289824
rect 218060 289876 218112 289882
rect 218060 289818 218112 289824
rect 215956 280022 215984 289818
rect 213920 280016 213972 280022
rect 213920 279958 213972 279964
rect 215944 280016 215996 280022
rect 215944 279958 215996 279964
rect 175924 276072 175976 276078
rect 175924 276014 175976 276020
rect 178684 276072 178736 276078
rect 178684 276014 178736 276020
rect 175936 260846 175964 276014
rect 213932 275330 213960 279958
rect 220096 276078 220124 313278
rect 223132 311914 223160 318242
rect 220176 311908 220228 311914
rect 220176 311850 220228 311856
rect 223120 311908 223172 311914
rect 223120 311850 223172 311856
rect 220188 292602 220216 311850
rect 220176 292596 220228 292602
rect 220176 292538 220228 292544
rect 218060 276072 218112 276078
rect 218060 276014 218112 276020
rect 220084 276072 220136 276078
rect 220084 276014 220136 276020
rect 204168 275324 204220 275330
rect 204168 275266 204220 275272
rect 213920 275324 213972 275330
rect 213920 275266 213972 275272
rect 204180 271930 204208 275266
rect 218072 273306 218100 276014
rect 217980 273278 218100 273306
rect 202144 271924 202196 271930
rect 202144 271866 202196 271872
rect 204168 271924 204220 271930
rect 204168 271866 204220 271872
rect 202156 266422 202184 271866
rect 217980 270570 218008 273278
rect 217968 270564 218020 270570
rect 217968 270506 218020 270512
rect 213368 270496 213420 270502
rect 213368 270438 213420 270444
rect 202144 266416 202196 266422
rect 202144 266358 202196 266364
rect 197728 266348 197780 266354
rect 197728 266290 197780 266296
rect 197740 261866 197768 266290
rect 213380 264246 213408 270438
rect 208400 264240 208452 264246
rect 208400 264182 208452 264188
rect 213368 264240 213420 264246
rect 213368 264182 213420 264188
rect 208412 262290 208440 264182
rect 208320 262262 208440 262290
rect 195244 261860 195296 261866
rect 195244 261802 195296 261808
rect 197728 261860 197780 261866
rect 197728 261802 197780 261808
rect 189080 261520 189132 261526
rect 189080 261462 189132 261468
rect 174268 260840 174320 260846
rect 174268 260782 174320 260788
rect 175924 260840 175976 260846
rect 175924 260782 175976 260788
rect 174280 252550 174308 260782
rect 189092 259486 189120 261462
rect 189080 259480 189132 259486
rect 189080 259422 189132 259428
rect 185584 259412 185636 259418
rect 185584 259354 185636 259360
rect 173164 252544 173216 252550
rect 173164 252486 173216 252492
rect 174268 252544 174320 252550
rect 174268 252486 174320 252492
rect 71780 251864 71832 251870
rect 71780 251806 71832 251812
rect 52460 249076 52512 249082
rect 52460 249018 52512 249024
rect 57980 249076 58032 249082
rect 57980 249018 58032 249024
rect 49700 247104 49752 247110
rect 49700 247046 49752 247052
rect 51724 247104 51776 247110
rect 51724 247046 51776 247052
rect 49712 243574 49740 247046
rect 52472 244338 52500 249018
rect 173176 247110 173204 252486
rect 185596 247110 185624 259354
rect 195256 256766 195284 261802
rect 208320 261526 208348 262262
rect 208308 261520 208360 261526
rect 208308 261462 208360 261468
rect 193864 256760 193916 256766
rect 193864 256702 193916 256708
rect 195244 256760 195296 256766
rect 195244 256702 195296 256708
rect 173164 247104 173216 247110
rect 173164 247046 173216 247052
rect 185584 247104 185636 247110
rect 185584 247046 185636 247052
rect 166264 247036 166316 247042
rect 166264 246978 166316 246984
rect 182916 247036 182968 247042
rect 182916 246978 182968 246984
rect 52380 244310 52500 244338
rect 49700 243568 49752 243574
rect 49700 243510 49752 243516
rect 52380 241738 52408 244310
rect 52368 241732 52420 241738
rect 52368 241674 52420 241680
rect 47676 241460 47728 241466
rect 47676 241402 47728 241408
rect 47584 241392 47636 241398
rect 47584 241334 47636 241340
rect 166276 240922 166304 246978
rect 166264 240916 166316 240922
rect 166264 240858 166316 240864
rect 182928 240854 182956 246978
rect 182916 240848 182968 240854
rect 182916 240790 182968 240796
rect 193876 240786 193904 256702
rect 193864 240780 193916 240786
rect 193864 240722 193916 240728
rect 47124 240168 47176 240174
rect 47124 240110 47176 240116
rect 395356 240009 395384 665790
rect 395528 646196 395580 646202
rect 395528 646138 395580 646144
rect 395436 475448 395488 475454
rect 395436 475390 395488 475396
rect 395448 240106 395476 475390
rect 395540 240145 395568 646138
rect 396724 378208 396776 378214
rect 396724 378150 396776 378156
rect 395526 240136 395582 240145
rect 395436 240100 395488 240106
rect 395526 240071 395582 240080
rect 396540 240100 396592 240106
rect 395436 240042 395488 240048
rect 396540 240042 396592 240048
rect 395342 240000 395398 240009
rect 395342 239935 395398 239944
rect 396552 238882 396580 240042
rect 396540 238876 396592 238882
rect 396540 238818 396592 238824
rect 45836 238808 45888 238814
rect 45836 238750 45888 238756
rect 396540 238740 396592 238746
rect 396540 238682 396592 238688
rect 45836 233232 45888 233238
rect 45836 233174 45888 233180
rect 45744 232212 45796 232218
rect 45744 232154 45796 232160
rect 45848 230382 45876 233174
rect 86316 232416 86368 232422
rect 86316 232358 86368 232364
rect 46848 232348 46900 232354
rect 46848 232290 46900 232296
rect 46940 232348 46992 232354
rect 46940 232290 46992 232296
rect 46204 232280 46256 232286
rect 46204 232222 46256 232228
rect 46216 230450 46244 232222
rect 46204 230444 46256 230450
rect 46204 230386 46256 230392
rect 45836 230376 45888 230382
rect 45836 230318 45888 230324
rect 46860 229094 46888 232290
rect 46952 230314 46980 232290
rect 53196 232212 53248 232218
rect 53196 232154 53248 232160
rect 52368 231192 52420 231198
rect 52368 231134 52420 231140
rect 48964 230444 49016 230450
rect 48964 230386 49016 230392
rect 47584 230376 47636 230382
rect 47584 230318 47636 230324
rect 46940 230308 46992 230314
rect 46940 230250 46992 230256
rect 46860 229066 46980 229094
rect 46952 228342 46980 229066
rect 46940 228336 46992 228342
rect 46940 228278 46992 228284
rect 47596 217462 47624 230318
rect 48976 220862 49004 230386
rect 52380 228138 52408 231134
rect 52460 230308 52512 230314
rect 52460 230250 52512 230256
rect 52368 228132 52420 228138
rect 52368 228074 52420 228080
rect 52472 223582 52500 230250
rect 52552 228336 52604 228342
rect 52552 228278 52604 228284
rect 52564 227050 52592 228278
rect 53208 227594 53236 232154
rect 86328 231198 86356 232358
rect 396552 232150 396580 238682
rect 394700 232144 394752 232150
rect 394606 232112 394662 232121
rect 394700 232086 394752 232092
rect 396540 232144 396592 232150
rect 396540 232086 396592 232092
rect 394606 232047 394662 232056
rect 86316 231192 86368 231198
rect 86316 231134 86368 231140
rect 153200 231192 153252 231198
rect 153200 231134 153252 231140
rect 390374 231160 390430 231169
rect 53840 228132 53892 228138
rect 53840 228074 53892 228080
rect 53196 227588 53248 227594
rect 53196 227530 53248 227536
rect 52552 227044 52604 227050
rect 52552 226986 52604 226992
rect 53852 226370 53880 228074
rect 53840 226364 53892 226370
rect 53840 226306 53892 226312
rect 52460 223576 52512 223582
rect 52460 223518 52512 223524
rect 55772 223576 55824 223582
rect 55772 223518 55824 223524
rect 47676 220856 47728 220862
rect 47676 220798 47728 220804
rect 48964 220856 49016 220862
rect 48964 220798 49016 220804
rect 47584 217456 47636 217462
rect 47584 217398 47636 217404
rect 47688 211138 47716 220798
rect 55784 220794 55812 223518
rect 53932 220788 53984 220794
rect 53932 220730 53984 220736
rect 55772 220788 55824 220794
rect 55772 220730 55824 220736
rect 53840 217456 53892 217462
rect 53840 217398 53892 217404
rect 53852 215354 53880 217398
rect 53944 215966 53972 220730
rect 53932 215960 53984 215966
rect 53932 215902 53984 215908
rect 53840 215348 53892 215354
rect 53840 215290 53892 215296
rect 47676 211132 47728 211138
rect 47676 211074 47728 211080
rect 51356 211132 51408 211138
rect 51356 211074 51408 211080
rect 46388 208412 46440 208418
rect 46388 208354 46440 208360
rect 46400 201482 46428 208354
rect 51368 204950 51396 211074
rect 51356 204944 51408 204950
rect 51356 204886 51408 204892
rect 46388 201476 46440 201482
rect 46388 201418 46440 201424
rect 47584 201476 47636 201482
rect 47584 201418 47636 201424
rect 47596 193186 47624 201418
rect 56612 195838 56640 230588
rect 57244 227588 57296 227594
rect 57244 227530 57296 227536
rect 56968 226296 57020 226302
rect 56968 226238 57020 226244
rect 56980 222902 57008 226238
rect 56968 222896 57020 222902
rect 56968 222838 57020 222844
rect 56692 215280 56744 215286
rect 56692 215222 56744 215228
rect 56704 211206 56732 215222
rect 57256 213246 57284 227530
rect 59268 227044 59320 227050
rect 59268 226986 59320 226992
rect 59280 223650 59308 226986
rect 59268 223644 59320 223650
rect 59268 223586 59320 223592
rect 66996 223576 67048 223582
rect 66996 223518 67048 223524
rect 58624 222896 58676 222902
rect 58624 222838 58676 222844
rect 58636 216714 58664 222838
rect 67008 220794 67036 223518
rect 62764 220788 62816 220794
rect 62764 220730 62816 220736
rect 66996 220788 67048 220794
rect 66996 220730 67048 220736
rect 69664 220788 69716 220794
rect 69664 220730 69716 220736
rect 58624 216708 58676 216714
rect 58624 216650 58676 216656
rect 57244 213240 57296 213246
rect 57244 213182 57296 213188
rect 56692 211200 56744 211206
rect 56692 211142 56744 211148
rect 62120 211132 62172 211138
rect 62120 211074 62172 211080
rect 62132 207670 62160 211074
rect 62120 207664 62172 207670
rect 62120 207606 62172 207612
rect 62776 205698 62804 220730
rect 65524 216640 65576 216646
rect 65524 216582 65576 216588
rect 63408 215960 63460 215966
rect 63408 215902 63460 215908
rect 63420 215234 63448 215902
rect 63420 215206 63540 215234
rect 63512 210254 63540 215206
rect 63500 210248 63552 210254
rect 63500 210190 63552 210196
rect 63500 207664 63552 207670
rect 63500 207606 63552 207612
rect 62764 205692 62816 205698
rect 62764 205634 62816 205640
rect 58624 204944 58676 204950
rect 58624 204886 58676 204892
rect 58636 196314 58664 204886
rect 63512 202230 63540 207606
rect 65536 207058 65564 216582
rect 65616 210248 65668 210254
rect 65616 210190 65668 210196
rect 65524 207052 65576 207058
rect 65524 206994 65576 207000
rect 65524 205624 65576 205630
rect 65524 205566 65576 205572
rect 63500 202224 63552 202230
rect 63500 202166 63552 202172
rect 65536 198150 65564 205566
rect 65628 205494 65656 210190
rect 69676 208418 69704 220730
rect 71044 213240 71096 213246
rect 71044 213182 71096 213188
rect 69664 208412 69716 208418
rect 69664 208354 69716 208360
rect 69664 206984 69716 206990
rect 69664 206926 69716 206932
rect 65616 205488 65668 205494
rect 65616 205430 65668 205436
rect 66904 205488 66956 205494
rect 66904 205430 66956 205436
rect 66260 202224 66312 202230
rect 66260 202166 66312 202172
rect 66272 198762 66300 202166
rect 66260 198756 66312 198762
rect 66260 198698 66312 198704
rect 65524 198144 65576 198150
rect 65524 198086 65576 198092
rect 66260 198144 66312 198150
rect 66260 198086 66312 198092
rect 58624 196308 58676 196314
rect 58624 196250 58676 196256
rect 61384 196308 61436 196314
rect 61384 196250 61436 196256
rect 56600 195832 56652 195838
rect 56600 195774 56652 195780
rect 47584 193180 47636 193186
rect 47584 193122 47636 193128
rect 48964 193180 49016 193186
rect 48964 193122 49016 193128
rect 45652 184884 45704 184890
rect 45652 184826 45704 184832
rect 48976 178090 49004 193122
rect 61396 188358 61424 196250
rect 66272 195498 66300 198086
rect 66916 196518 66944 205430
rect 68192 198756 68244 198762
rect 68192 198698 68244 198704
rect 66904 196512 66956 196518
rect 66904 196454 66956 196460
rect 68204 196042 68232 198698
rect 68284 196512 68336 196518
rect 68284 196454 68336 196460
rect 68192 196036 68244 196042
rect 68192 195978 68244 195984
rect 66260 195492 66312 195498
rect 66260 195434 66312 195440
rect 61384 188352 61436 188358
rect 61384 188294 61436 188300
rect 53104 184884 53156 184890
rect 53104 184826 53156 184832
rect 53116 180130 53144 184826
rect 53104 180124 53156 180130
rect 53104 180066 53156 180072
rect 63500 180124 63552 180130
rect 63500 180066 63552 180072
rect 48964 178084 49016 178090
rect 48964 178026 49016 178032
rect 49700 178084 49752 178090
rect 49700 178026 49752 178032
rect 49712 172514 49740 178026
rect 63512 177342 63540 180066
rect 63500 177336 63552 177342
rect 63500 177278 63552 177284
rect 49700 172508 49752 172514
rect 49700 172450 49752 172456
rect 53104 172508 53156 172514
rect 53104 172450 53156 172456
rect 45560 170400 45612 170406
rect 45560 170342 45612 170348
rect 53116 162994 53144 172450
rect 63500 170400 63552 170406
rect 63500 170342 63552 170348
rect 63512 163606 63540 170342
rect 63500 163600 63552 163606
rect 63500 163542 63552 163548
rect 66260 163600 66312 163606
rect 66260 163542 66312 163548
rect 53104 162988 53156 162994
rect 53104 162930 53156 162936
rect 55864 162988 55916 162994
rect 55864 162930 55916 162936
rect 55876 138582 55904 162930
rect 66272 160750 66300 163542
rect 66260 160744 66312 160750
rect 66260 160686 66312 160692
rect 68296 140826 68324 196454
rect 68376 195492 68428 195498
rect 68376 195434 68428 195440
rect 68388 166462 68416 195434
rect 68928 188352 68980 188358
rect 68928 188294 68980 188300
rect 68940 181490 68968 188294
rect 68928 181484 68980 181490
rect 68928 181426 68980 181432
rect 68376 166456 68428 166462
rect 68376 166398 68428 166404
rect 69676 159254 69704 206926
rect 71056 203590 71084 213182
rect 72424 208344 72476 208350
rect 72424 208286 72476 208292
rect 71044 203584 71096 203590
rect 71044 203526 71096 203532
rect 72436 199238 72464 208286
rect 72424 199232 72476 199238
rect 72424 199174 72476 199180
rect 75276 199232 75328 199238
rect 75276 199174 75328 199180
rect 71044 195968 71096 195974
rect 71044 195910 71096 195916
rect 71056 187950 71084 195910
rect 75288 195498 75316 199174
rect 86972 195906 87000 230588
rect 117240 228410 117268 230588
rect 146312 230574 146510 230602
rect 117228 228404 117280 228410
rect 117228 228346 117280 228352
rect 138664 228404 138716 228410
rect 138664 228346 138716 228352
rect 115848 218068 115900 218074
rect 115848 218010 115900 218016
rect 95148 203584 95200 203590
rect 95148 203526 95200 203532
rect 95160 200802 95188 203526
rect 95148 200796 95200 200802
rect 95148 200738 95200 200744
rect 104900 200796 104952 200802
rect 104900 200738 104952 200744
rect 104912 198558 104940 200738
rect 104900 198552 104952 198558
rect 104900 198494 104952 198500
rect 108304 198552 108356 198558
rect 108304 198494 108356 198500
rect 86960 195900 87012 195906
rect 86960 195842 87012 195848
rect 75276 195492 75328 195498
rect 75276 195434 75328 195440
rect 77944 195492 77996 195498
rect 77944 195434 77996 195440
rect 71044 187944 71096 187950
rect 71044 187886 71096 187892
rect 73160 187944 73212 187950
rect 73160 187886 73212 187892
rect 73172 184890 73200 187886
rect 73160 184884 73212 184890
rect 73160 184826 73212 184832
rect 75184 184884 75236 184890
rect 75184 184826 75236 184832
rect 75196 178158 75224 184826
rect 77956 179450 77984 195434
rect 108316 186658 108344 198494
rect 112444 187740 112496 187746
rect 112444 187682 112496 187688
rect 108304 186652 108356 186658
rect 108304 186594 108356 186600
rect 111064 186652 111116 186658
rect 111064 186594 111116 186600
rect 83464 181484 83516 181490
rect 83464 181426 83516 181432
rect 77944 179444 77996 179450
rect 77944 179386 77996 179392
rect 79324 179444 79376 179450
rect 79324 179386 79376 179392
rect 75184 178152 75236 178158
rect 75184 178094 75236 178100
rect 77208 178152 77260 178158
rect 77208 178094 77260 178100
rect 69756 177336 69808 177342
rect 69756 177278 69808 177284
rect 69664 159248 69716 159254
rect 69664 159190 69716 159196
rect 69768 150958 69796 177278
rect 77220 175302 77248 178094
rect 77208 175296 77260 175302
rect 77208 175238 77260 175244
rect 78680 175228 78732 175234
rect 78680 175170 78732 175176
rect 78692 172514 78720 175170
rect 78680 172508 78732 172514
rect 78680 172450 78732 172456
rect 79336 168774 79364 179386
rect 83476 173194 83504 181426
rect 83464 173188 83516 173194
rect 83464 173130 83516 173136
rect 91560 173188 91612 173194
rect 91560 173130 91612 173136
rect 80612 172508 80664 172514
rect 80612 172450 80664 172456
rect 79324 168768 79376 168774
rect 79324 168710 79376 168716
rect 80624 168502 80652 172450
rect 91572 170406 91600 173130
rect 111076 170746 111104 186594
rect 111064 170740 111116 170746
rect 111064 170682 111116 170688
rect 91560 170400 91612 170406
rect 91560 170342 91612 170348
rect 99380 170400 99432 170406
rect 99380 170342 99432 170348
rect 81532 168768 81584 168774
rect 81532 168710 81584 168716
rect 80612 168496 80664 168502
rect 80612 168438 80664 168444
rect 69848 166456 69900 166462
rect 69848 166398 69900 166404
rect 69860 154562 69888 166398
rect 81544 164218 81572 168710
rect 83464 168496 83516 168502
rect 83464 168438 83516 168444
rect 81532 164212 81584 164218
rect 81532 164154 81584 164160
rect 79324 160744 79376 160750
rect 79324 160686 79376 160692
rect 71688 159248 71740 159254
rect 71688 159190 71740 159196
rect 71700 157298 71728 159190
rect 79336 157350 79364 160686
rect 79324 157344 79376 157350
rect 71700 157270 71820 157298
rect 79324 157286 79376 157292
rect 69848 154556 69900 154562
rect 69848 154498 69900 154504
rect 71228 154556 71280 154562
rect 71228 154498 71280 154504
rect 69756 150952 69808 150958
rect 69756 150894 69808 150900
rect 71240 150482 71268 154498
rect 71792 153678 71820 157270
rect 71780 153672 71832 153678
rect 71780 153614 71832 153620
rect 75920 153672 75972 153678
rect 75920 153614 75972 153620
rect 72148 150952 72200 150958
rect 72148 150894 72200 150900
rect 71228 150476 71280 150482
rect 71228 150418 71280 150424
rect 72160 142866 72188 150894
rect 72424 150476 72476 150482
rect 72424 150418 72476 150424
rect 72148 142860 72200 142866
rect 72148 142802 72200 142808
rect 68284 140820 68336 140826
rect 68284 140762 68336 140768
rect 71412 140752 71464 140758
rect 71412 140694 71464 140700
rect 55864 138576 55916 138582
rect 55864 138518 55916 138524
rect 57888 138576 57940 138582
rect 57888 138518 57940 138524
rect 57900 134774 57928 138518
rect 71424 138038 71452 140694
rect 71412 138032 71464 138038
rect 71412 137974 71464 137980
rect 72436 136610 72464 150418
rect 75932 146334 75960 153614
rect 83476 148374 83504 168438
rect 83556 164212 83608 164218
rect 83556 164154 83608 164160
rect 83464 148368 83516 148374
rect 83464 148310 83516 148316
rect 83568 147694 83596 164154
rect 99392 163538 99420 170342
rect 99380 163532 99432 163538
rect 99380 163474 99432 163480
rect 85304 157344 85356 157350
rect 85304 157286 85356 157292
rect 85316 154562 85344 157286
rect 85304 154556 85356 154562
rect 85304 154498 85356 154504
rect 87604 154556 87656 154562
rect 87604 154498 87656 154504
rect 83556 147688 83608 147694
rect 83556 147630 83608 147636
rect 86224 147620 86276 147626
rect 86224 147562 86276 147568
rect 75920 146328 75972 146334
rect 75920 146270 75972 146276
rect 80704 146260 80756 146266
rect 80704 146202 80756 146208
rect 80716 138038 80744 146202
rect 86236 141166 86264 147562
rect 86224 141160 86276 141166
rect 86224 141102 86276 141108
rect 87616 139942 87644 154498
rect 88248 148368 88300 148374
rect 88248 148310 88300 148316
rect 88260 147642 88288 148310
rect 88260 147614 88380 147642
rect 88352 144906 88380 147614
rect 88340 144900 88392 144906
rect 88340 144842 88392 144848
rect 89996 144900 90048 144906
rect 89996 144842 90048 144848
rect 90008 141438 90036 144842
rect 91744 142860 91796 142866
rect 91744 142802 91796 142808
rect 89996 141432 90048 141438
rect 89996 141374 90048 141380
rect 91100 141160 91152 141166
rect 91100 141102 91152 141108
rect 87604 139936 87656 139942
rect 87604 139878 87656 139884
rect 89904 139936 89956 139942
rect 89904 139878 89956 139884
rect 80704 138032 80756 138038
rect 80704 137974 80756 137980
rect 73160 137964 73212 137970
rect 73160 137906 73212 137912
rect 86224 137964 86276 137970
rect 86224 137906 86276 137912
rect 72424 136604 72476 136610
rect 72424 136546 72476 136552
rect 73172 136542 73200 137906
rect 73804 136604 73856 136610
rect 73804 136546 73856 136552
rect 73160 136536 73212 136542
rect 73160 136478 73212 136484
rect 57888 134768 57940 134774
rect 57888 134710 57940 134716
rect 73816 127634 73844 136546
rect 75184 136536 75236 136542
rect 75184 136478 75236 136484
rect 73804 127628 73856 127634
rect 73804 127570 73856 127576
rect 75196 110566 75224 136478
rect 82084 127628 82136 127634
rect 82084 127570 82136 127576
rect 82096 121378 82124 127570
rect 86236 126886 86264 137906
rect 89916 136610 89944 139878
rect 89904 136604 89956 136610
rect 89904 136546 89956 136552
rect 91112 133142 91140 141102
rect 91756 138718 91784 142802
rect 98000 141432 98052 141438
rect 98000 141374 98052 141380
rect 91744 138712 91796 138718
rect 91744 138654 91796 138660
rect 97172 138712 97224 138718
rect 97172 138654 97224 138660
rect 95884 136604 95936 136610
rect 95884 136546 95936 136552
rect 91100 133136 91152 133142
rect 91100 133078 91152 133084
rect 93860 133136 93912 133142
rect 93860 133078 93912 133084
rect 93872 128654 93900 133078
rect 95896 130422 95924 136546
rect 97184 135250 97212 138654
rect 97172 135244 97224 135250
rect 97172 135186 97224 135192
rect 98012 133890 98040 141374
rect 102784 135244 102836 135250
rect 102784 135186 102836 135192
rect 98000 133884 98052 133890
rect 98000 133826 98052 133832
rect 101404 133884 101456 133890
rect 101404 133826 101456 133832
rect 95884 130416 95936 130422
rect 95884 130358 95936 130364
rect 93860 128648 93912 128654
rect 93860 128590 93912 128596
rect 97264 128648 97316 128654
rect 97264 128590 97316 128596
rect 86224 126880 86276 126886
rect 86224 126822 86276 126828
rect 88340 126880 88392 126886
rect 88340 126822 88392 126828
rect 88352 125526 88380 126822
rect 88340 125520 88392 125526
rect 88340 125462 88392 125468
rect 90364 125520 90416 125526
rect 90364 125462 90416 125468
rect 82084 121372 82136 121378
rect 82084 121314 82136 121320
rect 85856 121372 85908 121378
rect 85856 121314 85908 121320
rect 85868 117434 85896 121314
rect 85856 117428 85908 117434
rect 85856 117370 85908 117376
rect 87604 117428 87656 117434
rect 87604 117370 87656 117376
rect 87616 110974 87644 117370
rect 90376 115870 90404 125462
rect 97276 121854 97304 128590
rect 97264 121848 97316 121854
rect 97264 121790 97316 121796
rect 98736 121848 98788 121854
rect 98736 121790 98788 121796
rect 98748 121378 98776 121790
rect 98736 121372 98788 121378
rect 98736 121314 98788 121320
rect 100024 121372 100076 121378
rect 100024 121314 100076 121320
rect 90364 115864 90416 115870
rect 90364 115806 90416 115812
rect 93492 115864 93544 115870
rect 93492 115806 93544 115812
rect 93504 111722 93532 115806
rect 93492 111716 93544 111722
rect 93492 111658 93544 111664
rect 96528 111716 96580 111722
rect 96528 111658 96580 111664
rect 87604 110968 87656 110974
rect 87604 110910 87656 110916
rect 88708 110968 88760 110974
rect 88708 110910 88760 110916
rect 75184 110560 75236 110566
rect 75184 110502 75236 110508
rect 77944 110560 77996 110566
rect 77944 110502 77996 110508
rect 77956 96694 77984 110502
rect 88720 107642 88748 110910
rect 96540 108662 96568 111658
rect 100036 109002 100064 121314
rect 101416 109274 101444 133826
rect 101404 109268 101456 109274
rect 101404 109210 101456 109216
rect 102140 109268 102192 109274
rect 102140 109210 102192 109216
rect 100024 108996 100076 109002
rect 100024 108938 100076 108944
rect 96528 108656 96580 108662
rect 96528 108598 96580 108604
rect 97908 108656 97960 108662
rect 97908 108598 97960 108604
rect 88708 107636 88760 107642
rect 88708 107578 88760 107584
rect 97920 107522 97948 108598
rect 97920 107494 98040 107522
rect 98012 104854 98040 107494
rect 102152 105262 102180 109210
rect 102232 108996 102284 109002
rect 102232 108938 102284 108944
rect 102244 106282 102272 108938
rect 102232 106276 102284 106282
rect 102232 106218 102284 106224
rect 102140 105256 102192 105262
rect 102140 105198 102192 105204
rect 98000 104848 98052 104854
rect 98000 104790 98052 104796
rect 102796 97986 102824 135186
rect 108304 130416 108356 130422
rect 108304 130358 108356 130364
rect 108316 109002 108344 130358
rect 108304 108996 108356 109002
rect 108304 108938 108356 108944
rect 104624 105256 104676 105262
rect 104624 105198 104676 105204
rect 104636 99006 104664 105198
rect 104624 99000 104676 99006
rect 104624 98942 104676 98948
rect 106556 99000 106608 99006
rect 106556 98942 106608 98948
rect 102784 97980 102836 97986
rect 102784 97922 102836 97928
rect 105544 97980 105596 97986
rect 105544 97922 105596 97928
rect 77944 96688 77996 96694
rect 77944 96630 77996 96636
rect 81900 96620 81952 96626
rect 81900 96562 81952 96568
rect 81912 93838 81940 96562
rect 81900 93832 81952 93838
rect 81900 93774 81952 93780
rect 84844 93832 84896 93838
rect 84844 93774 84896 93780
rect 43536 74384 43588 74390
rect 43536 74326 43588 74332
rect 6918 74080 6974 74089
rect 6918 74015 6974 74024
rect 5172 73636 5224 73642
rect 5172 73578 5224 73584
rect 84856 73574 84884 93774
rect 105556 84862 105584 97922
rect 106568 95198 106596 98942
rect 106556 95192 106608 95198
rect 106556 95134 106608 95140
rect 108396 95192 108448 95198
rect 108396 95134 108448 95140
rect 108408 90166 108436 95134
rect 108396 90160 108448 90166
rect 108396 90102 108448 90108
rect 109776 90160 109828 90166
rect 109776 90102 109828 90108
rect 109788 86970 109816 90102
rect 109776 86964 109828 86970
rect 109776 86906 109828 86912
rect 110972 86964 111024 86970
rect 110972 86906 111024 86912
rect 105544 84856 105596 84862
rect 105544 84798 105596 84804
rect 110984 80034 111012 86906
rect 110972 80028 111024 80034
rect 110972 79970 111024 79976
rect 112456 73982 112484 187682
rect 115756 178084 115808 178090
rect 115756 178026 115808 178032
rect 115664 174344 115716 174350
rect 115664 174286 115716 174292
rect 114468 170740 114520 170746
rect 114468 170682 114520 170688
rect 114480 167686 114508 170682
rect 114468 167680 114520 167686
rect 114468 167622 114520 167628
rect 115112 166320 115164 166326
rect 115112 166262 115164 166268
rect 113732 163532 113784 163538
rect 113732 163474 113784 163480
rect 113744 136610 113772 163474
rect 114468 138032 114520 138038
rect 114468 137974 114520 137980
rect 114192 137556 114244 137562
rect 114192 137498 114244 137504
rect 114100 137352 114152 137358
rect 114006 137320 114062 137329
rect 113916 137284 113968 137290
rect 114100 137294 114152 137300
rect 114006 137255 114062 137264
rect 113916 137226 113968 137232
rect 113732 136604 113784 136610
rect 113732 136546 113784 136552
rect 113824 135992 113876 135998
rect 113824 135934 113876 135940
rect 113730 131200 113786 131209
rect 113730 131135 113732 131144
rect 113784 131135 113786 131144
rect 113732 131106 113784 131112
rect 113730 129024 113786 129033
rect 113730 128959 113786 128968
rect 113744 128382 113772 128959
rect 113732 128376 113784 128382
rect 113732 128318 113784 128324
rect 113638 127528 113694 127537
rect 113638 127463 113694 127472
rect 113652 127022 113680 127463
rect 113640 127016 113692 127022
rect 113640 126958 113692 126964
rect 113732 126948 113784 126954
rect 113732 126890 113784 126896
rect 113744 126857 113772 126890
rect 113730 126848 113786 126857
rect 113730 126783 113786 126792
rect 113548 125588 113600 125594
rect 113548 125530 113600 125536
rect 113560 125361 113588 125530
rect 113546 125352 113602 125361
rect 113546 125287 113602 125296
rect 113732 124160 113784 124166
rect 113732 124102 113784 124108
rect 113744 123865 113772 124102
rect 113730 123856 113786 123865
rect 113730 123791 113786 123800
rect 113364 122800 113416 122806
rect 113362 122768 113364 122777
rect 113416 122768 113418 122777
rect 113362 122703 113418 122712
rect 113732 121440 113784 121446
rect 113732 121382 113784 121388
rect 113744 121281 113772 121382
rect 113730 121272 113786 121281
rect 113730 121207 113786 121216
rect 113732 120080 113784 120086
rect 113732 120022 113784 120028
rect 113744 119785 113772 120022
rect 113730 119776 113786 119785
rect 113730 119711 113786 119720
rect 113640 118652 113692 118658
rect 113640 118594 113692 118600
rect 113652 118289 113680 118594
rect 113638 118280 113694 118289
rect 113638 118215 113694 118224
rect 113732 117292 113784 117298
rect 113732 117234 113784 117240
rect 113744 116793 113772 117234
rect 113730 116784 113786 116793
rect 113730 116719 113786 116728
rect 113732 115932 113784 115938
rect 113732 115874 113784 115880
rect 113744 115297 113772 115874
rect 113730 115288 113786 115297
rect 113730 115223 113786 115232
rect 113732 113144 113784 113150
rect 113730 113112 113732 113121
rect 113784 113112 113786 113121
rect 113730 113047 113786 113056
rect 113732 111784 113784 111790
rect 113730 111752 113732 111761
rect 113784 111752 113786 111761
rect 113730 111687 113786 111696
rect 113732 110424 113784 110430
rect 113730 110392 113732 110401
rect 113784 110392 113786 110401
rect 113730 110327 113786 110336
rect 113732 108996 113784 109002
rect 113732 108938 113784 108944
rect 113744 108905 113772 108938
rect 113730 108896 113786 108905
rect 113730 108831 113786 108840
rect 113548 107636 113600 107642
rect 113548 107578 113600 107584
rect 113560 107409 113588 107578
rect 113546 107400 113602 107409
rect 113546 107335 113602 107344
rect 113732 106276 113784 106282
rect 113732 106218 113784 106224
rect 113744 106185 113772 106218
rect 113730 106176 113786 106185
rect 113730 106111 113786 106120
rect 113364 104848 113416 104854
rect 113362 104816 113364 104825
rect 113416 104816 113418 104825
rect 113362 104751 113418 104760
rect 113836 101833 113864 135934
rect 113822 101824 113878 101833
rect 113822 101759 113878 101768
rect 113928 98841 113956 137226
rect 113914 98832 113970 98841
rect 113914 98767 113970 98776
rect 114020 91089 114048 137255
rect 114006 91080 114062 91089
rect 114006 91015 114062 91024
rect 114112 89729 114140 137294
rect 114098 89720 114154 89729
rect 114098 89655 114154 89664
rect 114204 88233 114232 137498
rect 114284 137488 114336 137494
rect 114284 137430 114336 137436
rect 114190 88224 114246 88233
rect 114190 88159 114246 88168
rect 114296 86873 114324 137430
rect 114376 137420 114428 137426
rect 114376 137362 114428 137368
rect 114282 86864 114338 86873
rect 114282 86799 114338 86808
rect 114388 85377 114416 137362
rect 114374 85368 114430 85377
rect 114374 85303 114430 85312
rect 114480 80889 114508 137974
rect 115124 133249 115152 166262
rect 115572 149728 115624 149734
rect 115572 149670 115624 149676
rect 115480 144220 115532 144226
rect 115480 144162 115532 144168
rect 115204 136672 115256 136678
rect 115204 136614 115256 136620
rect 115110 133240 115166 133249
rect 115110 133175 115166 133184
rect 114466 80880 114522 80889
rect 114466 80815 114522 80824
rect 114374 76664 114430 76673
rect 114374 76599 114430 76608
rect 112444 73976 112496 73982
rect 112444 73918 112496 73924
rect 84844 73568 84896 73574
rect 84844 73510 84896 73516
rect 85580 73568 85632 73574
rect 85580 73510 85632 73516
rect 85592 72622 85620 73510
rect 86224 72684 86276 72690
rect 86224 72626 86276 72632
rect 85580 72616 85632 72622
rect 22742 72584 22798 72593
rect 85580 72558 85632 72564
rect 22742 72519 22798 72528
rect 60740 72548 60792 72554
rect 5540 66904 5592 66910
rect 5540 66846 5592 66852
rect 3606 58576 3662 58585
rect 3606 58511 3662 58520
rect 3516 45552 3568 45558
rect 3514 45520 3516 45529
rect 3568 45520 3570 45529
rect 3514 45455 3570 45464
rect 3516 22704 3568 22710
rect 3516 22646 3568 22652
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 3528 6497 3556 22646
rect 5552 16574 5580 66846
rect 15200 54528 15252 54534
rect 15200 54470 15252 54476
rect 15212 16574 15240 54470
rect 5552 16546 6040 16574
rect 15212 16546 15976 16574
rect 3514 6488 3570 6497
rect 3514 6423 3570 6432
rect 4068 6180 4120 6186
rect 4068 6122 4120 6128
rect 1674 3496 1730 3505
rect 1674 3431 1730 3440
rect 2872 3460 2924 3466
rect 570 3360 626 3369
rect 570 3295 626 3304
rect 584 480 612 3295
rect 1688 480 1716 3431
rect 2872 3402 2924 3408
rect 2884 480 2912 3402
rect 4080 480 4108 6122
rect 5264 4888 5316 4894
rect 5264 4830 5316 4836
rect 5276 480 5304 4830
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6012 354 6040 16546
rect 14280 13116 14332 13122
rect 14280 13058 14332 13064
rect 9956 8968 10008 8974
rect 9956 8910 10008 8916
rect 8760 6248 8812 6254
rect 8760 6190 8812 6196
rect 7656 3528 7708 3534
rect 7656 3470 7708 3476
rect 7668 480 7696 3470
rect 8772 480 8800 6190
rect 9968 480 9996 8910
rect 11152 6656 11204 6662
rect 11152 6598 11204 6604
rect 11164 480 11192 6598
rect 13544 6316 13596 6322
rect 13544 6258 13596 6264
rect 12348 3596 12400 3602
rect 12348 3538 12400 3544
rect 12360 480 12388 3538
rect 13556 480 13584 6258
rect 6430 354 6542 480
rect 6012 326 6542 354
rect 6430 -960 6542 326
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14292 354 14320 13058
rect 15948 480 15976 16546
rect 19432 7676 19484 7682
rect 19432 7618 19484 7624
rect 18234 6216 18290 6225
rect 18234 6151 18290 6160
rect 17038 3632 17094 3641
rect 17038 3567 17094 3576
rect 17052 480 17080 3567
rect 18248 480 18276 6151
rect 19444 480 19472 7618
rect 22756 4894 22784 72519
rect 60740 72490 60792 72496
rect 25504 72480 25556 72486
rect 25504 72422 25556 72428
rect 25320 10328 25372 10334
rect 25320 10270 25372 10276
rect 24216 9036 24268 9042
rect 24216 8978 24268 8984
rect 23020 7608 23072 7614
rect 23020 7550 23072 7556
rect 22744 4888 22796 4894
rect 22744 4830 22796 4836
rect 21824 4820 21876 4826
rect 21824 4762 21876 4768
rect 20628 3256 20680 3262
rect 20628 3198 20680 3204
rect 20640 480 20668 3198
rect 21836 480 21864 4762
rect 23032 480 23060 7550
rect 24228 480 24256 8978
rect 25332 480 25360 10270
rect 25516 3262 25544 72422
rect 35900 18624 35952 18630
rect 35900 18566 35952 18572
rect 35912 16574 35940 18566
rect 60752 16574 60780 72490
rect 81440 25560 81492 25566
rect 81440 25502 81492 25508
rect 81452 16574 81480 25502
rect 35912 16546 36032 16574
rect 60752 16546 61608 16574
rect 81452 16546 81664 16574
rect 31944 10396 31996 10402
rect 31944 10338 31996 10344
rect 31300 9104 31352 9110
rect 31300 9046 31352 9052
rect 27712 7744 27764 7750
rect 27712 7686 27764 7692
rect 26516 4888 26568 4894
rect 26516 4830 26568 4836
rect 25504 3256 25556 3262
rect 25504 3198 25556 3204
rect 26528 480 26556 4830
rect 27724 480 27752 7686
rect 30104 6384 30156 6390
rect 30104 6326 30156 6332
rect 28908 4956 28960 4962
rect 28908 4898 28960 4904
rect 28920 480 28948 4898
rect 30116 480 30144 6326
rect 31312 480 31340 9046
rect 14710 354 14822 480
rect 14292 326 14822 354
rect 14710 -960 14822 326
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 31956 354 31984 10338
rect 34794 8936 34850 8945
rect 34794 8871 34850 8880
rect 33600 5024 33652 5030
rect 33600 4966 33652 4972
rect 33612 480 33640 4966
rect 34808 480 34836 8871
rect 36004 480 36032 16546
rect 46664 10464 46716 10470
rect 46664 10406 46716 10412
rect 43076 9376 43128 9382
rect 43076 9318 43128 9324
rect 41880 9172 41932 9178
rect 41880 9114 41932 9120
rect 38382 9072 38438 9081
rect 38382 9007 38438 9016
rect 37186 4856 37242 4865
rect 37186 4791 37242 4800
rect 37200 480 37228 4791
rect 38396 480 38424 9007
rect 40684 6452 40736 6458
rect 40684 6394 40736 6400
rect 39580 3664 39632 3670
rect 39580 3606 39632 3612
rect 39592 480 39620 3606
rect 40696 480 40724 6394
rect 41892 480 41920 9114
rect 43088 480 43116 9318
rect 45468 9240 45520 9246
rect 45468 9182 45520 9188
rect 44272 6520 44324 6526
rect 44272 6462 44324 6468
rect 44284 480 44312 6462
rect 45480 480 45508 9182
rect 46676 480 46704 10406
rect 60832 9512 60884 9518
rect 60832 9454 60884 9460
rect 57244 9444 57296 9450
rect 57244 9386 57296 9392
rect 50160 9308 50212 9314
rect 50160 9250 50212 9256
rect 48964 6588 49016 6594
rect 48964 6530 49016 6536
rect 47860 3732 47912 3738
rect 47860 3674 47912 3680
rect 47872 480 47900 3674
rect 48976 480 49004 6530
rect 50172 480 50200 9250
rect 53746 9208 53802 9217
rect 53746 9143 53802 9152
rect 52550 6352 52606 6361
rect 52550 6287 52606 6296
rect 51356 3800 51408 3806
rect 51356 3742 51408 3748
rect 51368 480 51396 3742
rect 52564 480 52592 6287
rect 53760 480 53788 9143
rect 56046 6488 56102 6497
rect 56046 6423 56102 6432
rect 54942 3768 54998 3777
rect 54942 3703 54998 3712
rect 54956 480 54984 3703
rect 56060 480 56088 6423
rect 57256 480 57284 9386
rect 59636 6724 59688 6730
rect 59636 6666 59688 6672
rect 58440 3868 58492 3874
rect 58440 3810 58492 3816
rect 58452 480 58480 3810
rect 59648 480 59676 6666
rect 60844 480 60872 9454
rect 32374 354 32486 480
rect 31956 326 32486 354
rect 32374 -960 32486 326
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61580 354 61608 16546
rect 75000 10736 75052 10742
rect 75000 10678 75052 10684
rect 67640 10600 67692 10606
rect 67640 10542 67692 10548
rect 64328 10532 64380 10538
rect 64328 10474 64380 10480
rect 63224 7812 63276 7818
rect 63224 7754 63276 7760
rect 63236 480 63264 7754
rect 64340 480 64368 10474
rect 66720 7880 66772 7886
rect 66720 7822 66772 7828
rect 65524 5092 65576 5098
rect 65524 5034 65576 5040
rect 65536 480 65564 5034
rect 66732 480 66760 7822
rect 61998 354 62110 480
rect 61580 326 62110 354
rect 61998 -960 62110 326
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67652 354 67680 10542
rect 71502 10296 71558 10305
rect 71502 10231 71558 10240
rect 70306 7576 70362 7585
rect 70306 7511 70362 7520
rect 69112 3936 69164 3942
rect 69112 3878 69164 3884
rect 69124 480 69152 3878
rect 70320 480 70348 7511
rect 71516 480 71544 10231
rect 73804 7948 73856 7954
rect 73804 7890 73856 7896
rect 72608 5160 72660 5166
rect 72608 5102 72660 5108
rect 72620 480 72648 5102
rect 73816 480 73844 7890
rect 75012 480 75040 10678
rect 78128 10668 78180 10674
rect 78128 10610 78180 10616
rect 77392 8016 77444 8022
rect 77392 7958 77444 7964
rect 76196 5228 76248 5234
rect 76196 5170 76248 5176
rect 76208 480 76236 5170
rect 77404 480 77432 7958
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78140 354 78168 10610
rect 80888 8084 80940 8090
rect 80888 8026 80940 8032
rect 79692 4004 79744 4010
rect 79692 3946 79744 3952
rect 79704 480 79732 3946
rect 80900 480 80928 8026
rect 78558 354 78670 480
rect 78140 326 78670 354
rect 78558 -960 78670 326
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 81636 354 81664 16546
rect 84476 8152 84528 8158
rect 84476 8094 84528 8100
rect 83280 4072 83332 4078
rect 83280 4014 83332 4020
rect 83292 480 83320 4014
rect 84488 480 84516 8094
rect 86236 6662 86264 72626
rect 93952 72616 94004 72622
rect 93952 72558 94004 72564
rect 93964 71670 93992 72558
rect 93952 71664 94004 71670
rect 93952 71606 94004 71612
rect 114388 60722 114416 76599
rect 114466 75440 114522 75449
rect 114466 75375 114522 75384
rect 114376 60716 114428 60722
rect 114376 60658 114428 60664
rect 113180 51128 113232 51134
rect 113180 51070 113232 51076
rect 106280 43444 106332 43450
rect 106280 43386 106332 43392
rect 106292 16574 106320 43386
rect 113192 16574 113220 51070
rect 114480 22778 114508 75375
rect 115216 73914 115244 136614
rect 115388 135924 115440 135930
rect 115388 135866 115440 135872
rect 115296 134564 115348 134570
rect 115296 134506 115348 134512
rect 115308 103193 115336 134506
rect 115294 103184 115350 103193
rect 115294 103119 115350 103128
rect 115400 92449 115428 135866
rect 115492 93809 115520 144162
rect 115584 95169 115612 149670
rect 115676 96733 115704 174286
rect 115662 96724 115718 96733
rect 115662 96659 115718 96668
rect 115570 95160 115626 95169
rect 115570 95095 115626 95104
rect 115478 93800 115534 93809
rect 115478 93735 115534 93744
rect 115386 92440 115442 92449
rect 115386 92375 115442 92384
rect 115768 81773 115796 178026
rect 115860 83269 115888 218010
rect 138676 195974 138704 228346
rect 146312 197418 146340 230574
rect 153212 228410 153240 231134
rect 177856 231124 177908 231130
rect 390374 231095 390430 231104
rect 177856 231066 177908 231072
rect 176672 229770 176700 230588
rect 166264 229764 166316 229770
rect 166264 229706 166316 229712
rect 176660 229764 176712 229770
rect 176660 229706 176712 229712
rect 157984 228472 158036 228478
rect 157984 228414 158036 228420
rect 153200 228404 153252 228410
rect 153200 228346 153252 228352
rect 155960 199436 156012 199442
rect 155960 199378 156012 199384
rect 148968 198008 149020 198014
rect 148968 197950 149020 197956
rect 146142 197390 146340 197418
rect 148980 197404 149008 197950
rect 155972 197470 156000 199378
rect 154488 197464 154540 197470
rect 154146 197412 154488 197418
rect 154146 197406 154540 197412
rect 155960 197464 156012 197470
rect 155960 197406 156012 197412
rect 154146 197390 154528 197406
rect 157996 197334 158024 228414
rect 165068 228404 165120 228410
rect 165068 228346 165120 228352
rect 165080 227254 165108 228346
rect 165068 227248 165120 227254
rect 165068 227190 165120 227196
rect 152740 197328 152792 197334
rect 152582 197276 152740 197282
rect 152582 197270 152792 197276
rect 157984 197328 158036 197334
rect 157984 197270 158036 197276
rect 152582 197254 152780 197270
rect 166276 196790 166304 229706
rect 170404 227248 170456 227254
rect 170404 227190 170456 227196
rect 170416 198762 170444 227190
rect 175372 213988 175424 213994
rect 175372 213930 175424 213936
rect 170404 198756 170456 198762
rect 170404 198698 170456 198704
rect 171784 198756 171836 198762
rect 171784 198698 171836 198704
rect 147956 196784 148008 196790
rect 147798 196732 147956 196738
rect 147798 196726 148008 196732
rect 166264 196784 166316 196790
rect 166264 196726 166316 196732
rect 147798 196710 147996 196726
rect 160836 196716 160888 196722
rect 160836 196658 160888 196664
rect 151176 196648 151228 196654
rect 150926 196596 151176 196602
rect 150926 196590 151228 196596
rect 150926 196574 151216 196590
rect 140424 196030 140530 196058
rect 157366 196030 157564 196058
rect 138664 195968 138716 195974
rect 138110 195936 138166 195945
rect 140424 195945 140452 196030
rect 157536 195974 157564 196030
rect 141424 195968 141476 195974
rect 138664 195910 138716 195916
rect 140410 195936 140466 195945
rect 138110 195871 138166 195880
rect 139400 195900 139452 195906
rect 138124 195838 138152 195871
rect 140410 195871 140466 195880
rect 141422 195936 141424 195945
rect 157524 195968 157576 195974
rect 141476 195936 141478 195945
rect 158916 195937 158944 196044
rect 160848 195945 160876 196658
rect 157524 195910 157576 195916
rect 158902 195928 158958 195937
rect 141422 195871 141478 195880
rect 157432 195900 157484 195906
rect 139400 195842 139452 195848
rect 158902 195863 158958 195872
rect 160834 195936 160890 195945
rect 160834 195871 160890 195880
rect 157432 195842 157484 195848
rect 138112 195832 138164 195838
rect 138112 195774 138164 195780
rect 139412 195537 139440 195842
rect 157154 195664 157210 195673
rect 157444 195650 157472 195842
rect 157210 195622 157472 195650
rect 157154 195599 157210 195608
rect 139398 195528 139454 195537
rect 139398 195463 139454 195472
rect 140870 191856 140926 191865
rect 140870 191791 140926 191800
rect 140778 191720 140834 191729
rect 140778 191655 140834 191664
rect 140792 184249 140820 191655
rect 140778 184240 140834 184249
rect 135260 184204 135312 184210
rect 140778 184175 140834 184184
rect 135260 184146 135312 184152
rect 117320 180192 117372 180198
rect 117320 180134 117372 180140
rect 115940 142860 115992 142866
rect 115940 142802 115992 142808
rect 115952 100337 115980 142802
rect 116584 136604 116636 136610
rect 116584 136546 116636 136552
rect 115938 100328 115994 100337
rect 115938 100263 115994 100272
rect 115846 83260 115902 83269
rect 115846 83195 115902 83204
rect 115754 81764 115810 81773
rect 115754 81699 115810 81708
rect 115848 80028 115900 80034
rect 115848 79970 115900 79976
rect 115860 77262 115888 79970
rect 116490 78432 116546 78441
rect 116490 78367 116546 78376
rect 115860 77234 115980 77262
rect 115952 75682 115980 77234
rect 115940 75676 115992 75682
rect 115940 75618 115992 75624
rect 116504 75585 116532 78367
rect 116490 75576 116546 75585
rect 116490 75511 116546 75520
rect 115204 73908 115256 73914
rect 115204 73850 115256 73856
rect 116596 70990 116624 136546
rect 117332 134994 117360 180134
rect 122104 180124 122156 180130
rect 122104 180066 122156 180072
rect 120724 178696 120776 178702
rect 120724 178638 120776 178644
rect 120080 177336 120132 177342
rect 120080 177278 120132 177284
rect 117412 169788 117464 169794
rect 117412 169730 117464 169736
rect 117424 166326 117452 169730
rect 117412 166320 117464 166326
rect 117412 166262 117464 166268
rect 120092 151814 120120 177278
rect 120092 151786 120488 151814
rect 119344 137964 119396 137970
rect 119344 137906 119396 137912
rect 117332 134966 117806 134994
rect 119356 134980 119384 137906
rect 120460 134994 120488 151786
rect 120736 137970 120764 178638
rect 121460 175976 121512 175982
rect 121460 175918 121512 175924
rect 121472 151814 121500 175918
rect 122116 169794 122144 180066
rect 122840 176112 122892 176118
rect 122840 176054 122892 176060
rect 122104 169788 122156 169794
rect 122104 169730 122156 169736
rect 122852 151814 122880 176054
rect 125600 174548 125652 174554
rect 125600 174490 125652 174496
rect 121472 151786 122144 151814
rect 122852 151786 123616 151814
rect 120724 137964 120776 137970
rect 120724 137906 120776 137912
rect 122116 134994 122144 151786
rect 123588 134994 123616 151786
rect 120460 134966 120934 134994
rect 122116 134966 122498 134994
rect 123588 134966 124062 134994
rect 125612 134980 125640 174490
rect 129740 173936 129792 173942
rect 129740 173878 129792 173884
rect 126980 173188 127032 173194
rect 126980 173130 127032 173136
rect 126992 134994 127020 173130
rect 128360 171148 128412 171154
rect 128360 171090 128412 171096
rect 128372 134994 128400 171090
rect 129752 151814 129780 173878
rect 133880 172168 133932 172174
rect 133880 172110 133932 172116
rect 131120 171964 131172 171970
rect 131120 171906 131172 171912
rect 131132 151814 131160 171906
rect 132500 171556 132552 171562
rect 132500 171498 132552 171504
rect 132512 151814 132540 171498
rect 133892 151814 133920 172110
rect 135272 151814 135300 184146
rect 140884 184113 140912 191791
rect 144366 191040 144422 191049
rect 144288 190998 144366 191026
rect 140962 190904 141018 190913
rect 140962 190839 141018 190848
rect 140976 184385 141004 190839
rect 140962 184376 141018 184385
rect 140962 184311 141018 184320
rect 142436 184272 142488 184278
rect 142436 184214 142488 184220
rect 142448 184212 142476 184214
rect 140870 184104 140926 184113
rect 140870 184039 140926 184048
rect 144288 183526 144316 190998
rect 144366 190975 144422 190984
rect 157340 189916 157392 189922
rect 157340 189858 157392 189864
rect 145838 189816 145894 189825
rect 145894 189774 145958 189802
rect 145838 189751 145894 189760
rect 144826 189272 144882 189281
rect 144826 189207 144882 189216
rect 136376 182158 136758 182186
rect 136376 180198 136404 182158
rect 144840 182050 144868 189207
rect 157352 189009 157380 189858
rect 166106 189366 166212 189394
rect 157338 189000 157394 189009
rect 157338 188935 157394 188944
rect 166184 187678 166212 189366
rect 166172 187672 166224 187678
rect 166172 187614 166224 187620
rect 144918 182064 144974 182073
rect 144840 182022 144918 182050
rect 144918 181999 144974 182008
rect 141238 181112 141294 181121
rect 141238 181047 141294 181056
rect 136468 180934 136758 180962
rect 136364 180192 136416 180198
rect 136364 180134 136416 180140
rect 136364 178832 136416 178838
rect 136364 178774 136416 178780
rect 135996 178152 136048 178158
rect 135996 178094 136048 178100
rect 136008 177342 136036 178094
rect 135996 177336 136048 177342
rect 135996 177278 136048 177284
rect 135720 176180 135772 176186
rect 135720 176122 135772 176128
rect 135732 174554 135760 176122
rect 136376 175982 136404 178774
rect 136468 178702 136496 180934
rect 141252 180402 141280 181047
rect 144642 180976 144698 180985
rect 144578 180934 144642 180962
rect 144642 180911 144698 180920
rect 141240 180396 141292 180402
rect 141240 180338 141292 180344
rect 136560 179982 136758 180010
rect 136456 178696 136508 178702
rect 136456 178638 136508 178644
rect 136560 178158 136588 179982
rect 142666 179072 142722 179081
rect 136744 178838 136772 179044
rect 142666 179007 142722 179016
rect 144090 178936 144146 178945
rect 144090 178871 144146 178880
rect 136732 178832 136784 178838
rect 136732 178774 136784 178780
rect 141698 178800 141754 178809
rect 141698 178735 141754 178744
rect 136548 178152 136600 178158
rect 136548 178094 136600 178100
rect 136468 177942 136758 177970
rect 136468 176118 136496 177942
rect 136560 176990 136758 177018
rect 136560 176186 136588 176990
rect 136548 176180 136600 176186
rect 136548 176122 136600 176128
rect 136456 176112 136508 176118
rect 136456 176054 136508 176060
rect 136560 176038 136758 176066
rect 136364 175976 136416 175982
rect 136364 175918 136416 175924
rect 135720 174548 135772 174554
rect 135720 174490 135772 174496
rect 136560 173894 136588 176038
rect 136560 173866 136680 173894
rect 136652 173194 136680 173866
rect 136640 173188 136692 173194
rect 136640 173130 136692 173136
rect 136744 171154 136772 174964
rect 141712 174758 141740 178735
rect 141790 178664 141846 178673
rect 141790 178599 141846 178608
rect 141804 174758 141832 178599
rect 144104 175438 144132 178871
rect 154396 178220 154448 178226
rect 154396 178162 154448 178168
rect 157800 178220 157852 178226
rect 157800 178162 157852 178168
rect 154408 178106 154436 178162
rect 157812 178129 157840 178162
rect 153948 178090 154436 178106
rect 153936 178084 154436 178090
rect 153988 178078 154436 178084
rect 157798 178120 157854 178129
rect 157798 178055 157854 178064
rect 158534 178120 158590 178129
rect 158590 178090 158668 178106
rect 158590 178084 158680 178090
rect 158590 178078 158628 178084
rect 158534 178055 158590 178064
rect 153936 178026 153988 178032
rect 158628 178026 158680 178032
rect 149980 175568 150032 175574
rect 149980 175510 150032 175516
rect 149992 175508 150020 175510
rect 144460 175500 144512 175506
rect 144460 175442 144512 175448
rect 144092 175432 144144 175438
rect 144092 175374 144144 175380
rect 141700 174752 141752 174758
rect 141700 174694 141752 174700
rect 141792 174752 141844 174758
rect 141792 174694 141844 174700
rect 137284 173936 137336 173942
rect 137336 173884 137586 173890
rect 137284 173878 137586 173884
rect 137296 173862 137586 173878
rect 138676 171970 138704 173196
rect 138664 171964 138716 171970
rect 138664 171906 138716 171912
rect 139688 171562 139716 173196
rect 140792 172174 140820 173196
rect 142436 172848 142488 172854
rect 142436 172790 142488 172796
rect 140780 172168 140832 172174
rect 140780 172110 140832 172116
rect 140780 171828 140832 171834
rect 140780 171770 140832 171776
rect 139676 171556 139728 171562
rect 139676 171498 139728 171504
rect 136732 171148 136784 171154
rect 136732 171090 136784 171096
rect 138664 167680 138716 167686
rect 138664 167622 138716 167628
rect 138676 160750 138704 167622
rect 138664 160744 138716 160750
rect 138664 160686 138716 160692
rect 140792 151814 140820 171770
rect 129752 151786 129872 151814
rect 131132 151786 131528 151814
rect 132512 151786 133000 151814
rect 133892 151786 134656 151814
rect 135272 151786 136128 151814
rect 140792 151786 140912 151814
rect 129844 134994 129872 151786
rect 131500 134994 131528 151786
rect 132972 134994 133000 151786
rect 134628 134994 134656 151786
rect 136100 134994 136128 151786
rect 139674 138000 139730 138009
rect 139674 137935 139730 137944
rect 138112 136808 138164 136814
rect 138112 136750 138164 136756
rect 126992 134966 127190 134994
rect 128372 134966 128754 134994
rect 129844 134966 130318 134994
rect 131500 134966 131882 134994
rect 132972 134966 133446 134994
rect 134628 134966 135010 134994
rect 136100 134966 136574 134994
rect 138124 134980 138152 136750
rect 139688 134980 139716 137935
rect 140884 134994 140912 151786
rect 142448 137086 142476 172790
rect 142632 161474 142660 173196
rect 143448 172984 143500 172990
rect 143448 172926 143500 172932
rect 142540 161446 142660 161474
rect 142436 137080 142488 137086
rect 142436 137022 142488 137028
rect 142540 136814 142568 161446
rect 143460 142154 143488 172926
rect 143540 172916 143592 172922
rect 143540 172858 143592 172864
rect 143552 151814 143580 172858
rect 143552 151786 144040 151814
rect 143184 142126 143488 142154
rect 142528 136808 142580 136814
rect 142528 136750 142580 136756
rect 143184 134994 143212 142126
rect 140884 134966 141266 134994
rect 142830 134966 143212 134994
rect 144012 134994 144040 151786
rect 144472 137630 144500 175442
rect 153936 175432 153988 175438
rect 153988 175380 154436 175386
rect 153936 175374 154436 175380
rect 153948 175358 154436 175374
rect 154408 175302 154436 175358
rect 154396 175296 154448 175302
rect 154396 175238 154448 175244
rect 156512 175296 156564 175302
rect 156512 175238 156564 175244
rect 153476 174616 153528 174622
rect 147494 174584 147550 174593
rect 153476 174558 153528 174564
rect 147494 174519 147550 174528
rect 144932 171834 144960 173196
rect 145668 172990 145696 173196
rect 145656 172984 145708 172990
rect 145656 172926 145708 172932
rect 146484 172984 146536 172990
rect 146484 172926 146536 172932
rect 144920 171828 144972 171834
rect 144920 171770 144972 171776
rect 146496 151814 146524 172926
rect 146680 172922 146708 173196
rect 146668 172916 146720 172922
rect 146668 172858 146720 172864
rect 147508 153202 147536 174519
rect 153488 173942 153516 174558
rect 153476 173936 153528 173942
rect 153476 173878 153528 173884
rect 147600 172854 147628 173196
rect 148612 172990 148640 173196
rect 148600 172984 148652 172990
rect 148600 172926 148652 172932
rect 147588 172848 147640 172854
rect 147588 172790 147640 172796
rect 149624 161474 149652 173196
rect 150636 166994 150664 173196
rect 149532 161446 149652 161474
rect 150452 166966 150664 166994
rect 147680 160744 147732 160750
rect 147680 160686 147732 160692
rect 147692 153882 147720 160686
rect 147680 153876 147732 153882
rect 147680 153818 147732 153824
rect 147496 153196 147548 153202
rect 147496 153138 147548 153144
rect 149244 153196 149296 153202
rect 149244 153138 149296 153144
rect 146496 151786 147168 151814
rect 144460 137624 144512 137630
rect 144460 137566 144512 137572
rect 145932 137080 145984 137086
rect 145932 137022 145984 137028
rect 144012 134966 144394 134994
rect 145944 134980 145972 137022
rect 147140 134994 147168 151786
rect 149256 148374 149284 153138
rect 149244 148368 149296 148374
rect 149244 148310 149296 148316
rect 149532 142154 149560 161446
rect 149440 142126 149560 142154
rect 149440 134994 149468 142126
rect 147140 134966 147522 134994
rect 149086 134966 149468 134994
rect 150452 134994 150480 166966
rect 151648 161474 151676 173196
rect 152660 161474 152688 173196
rect 150544 161446 151676 161474
rect 152476 161446 152688 161474
rect 153488 173182 153686 173210
rect 150544 137970 150572 161446
rect 152476 137970 152504 161446
rect 150532 137964 150584 137970
rect 150532 137906 150584 137912
rect 152188 137964 152240 137970
rect 152188 137906 152240 137912
rect 152464 137964 152516 137970
rect 152464 137906 152516 137912
rect 150452 134966 150650 134994
rect 152200 134980 152228 137906
rect 153488 136814 153516 173182
rect 156524 172990 156552 175238
rect 162492 174548 162544 174554
rect 162492 174490 162544 174496
rect 161414 173194 161520 173210
rect 161414 173188 161532 173194
rect 161414 173182 161480 173188
rect 161480 173130 161532 173136
rect 159456 173052 159508 173058
rect 159456 172994 159508 173000
rect 156512 172984 156564 172990
rect 156512 172926 156564 172932
rect 158444 172984 158496 172990
rect 158444 172926 158496 172932
rect 155224 148368 155276 148374
rect 155224 148310 155276 148316
rect 153752 137964 153804 137970
rect 153752 137906 153804 137912
rect 153476 136808 153528 136814
rect 153476 136750 153528 136756
rect 153764 134980 153792 137906
rect 155236 137698 155264 148310
rect 155224 137692 155276 137698
rect 155224 137634 155276 137640
rect 156880 137624 156932 137630
rect 156880 137566 156932 137572
rect 155316 136808 155368 136814
rect 155316 136750 155368 136756
rect 155328 134980 155356 136750
rect 156892 134980 156920 137566
rect 158456 134980 158484 172926
rect 159364 153876 159416 153882
rect 159364 153818 159416 153824
rect 159376 149802 159404 153818
rect 159468 151814 159496 172994
rect 162504 151814 162532 174490
rect 159468 151786 159680 151814
rect 162504 151786 162808 151814
rect 159364 149796 159416 149802
rect 159364 149738 159416 149744
rect 159652 134994 159680 151786
rect 161570 137728 161626 137737
rect 161570 137663 161626 137672
rect 159652 134966 160034 134994
rect 161584 134980 161612 137663
rect 162780 137034 162808 151786
rect 163516 137630 163544 175100
rect 163504 137624 163556 137630
rect 163504 137566 163556 137572
rect 162780 137006 162900 137034
rect 162872 134994 162900 137006
rect 163608 136882 163636 173196
rect 164528 173182 164634 173210
rect 166540 173188 166592 173194
rect 164528 137970 164556 173182
rect 166540 173130 166592 173136
rect 166552 161474 166580 173130
rect 166460 161446 166580 161474
rect 166264 149796 166316 149802
rect 166264 149738 166316 149744
rect 166276 141166 166304 149738
rect 166264 141160 166316 141166
rect 166264 141102 166316 141108
rect 164516 137964 164568 137970
rect 164516 137906 164568 137912
rect 164700 137692 164752 137698
rect 164700 137634 164752 137640
rect 163596 136876 163648 136882
rect 163596 136818 163648 136824
rect 162872 134966 163162 134994
rect 164712 134980 164740 137634
rect 166460 134994 166488 161446
rect 171796 147694 171824 198698
rect 175280 162920 175332 162926
rect 175280 162862 175332 162868
rect 171784 147688 171836 147694
rect 171784 147630 171836 147636
rect 173164 147688 173216 147694
rect 173164 147630 173216 147636
rect 169760 141160 169812 141166
rect 169760 141102 169812 141108
rect 167826 137592 167882 137601
rect 167826 137527 167882 137536
rect 166290 134966 166488 134994
rect 167840 134980 167868 137527
rect 169390 137456 169446 137465
rect 169390 137391 169446 137400
rect 169404 134980 169432 137391
rect 169772 136542 169800 141102
rect 173176 140350 173204 147630
rect 173164 140344 173216 140350
rect 173164 140286 173216 140292
rect 172520 137964 172572 137970
rect 172520 137906 172572 137912
rect 170956 136876 171008 136882
rect 170956 136818 171008 136824
rect 169760 136536 169812 136542
rect 169760 136478 169812 136484
rect 170968 134980 170996 136818
rect 172532 134980 172560 137906
rect 174084 137624 174136 137630
rect 174084 137566 174136 137572
rect 174096 134980 174124 137566
rect 175292 128330 175320 162862
rect 175384 151814 175412 213930
rect 175384 151786 175596 151814
rect 175464 136468 175516 136474
rect 175464 136410 175516 136416
rect 175372 133952 175424 133958
rect 175372 133894 175424 133900
rect 175384 129985 175412 133894
rect 175370 129976 175426 129985
rect 175370 129911 175426 129920
rect 175370 128344 175426 128353
rect 175292 128302 175370 128330
rect 175370 128279 175426 128288
rect 175476 111897 175504 136410
rect 175568 132494 175596 151786
rect 177304 140344 177356 140350
rect 177304 140286 177356 140292
rect 175924 136536 175976 136542
rect 175924 136478 175976 136484
rect 175568 132466 175688 132494
rect 175554 132424 175610 132433
rect 175554 132359 175610 132368
rect 175462 111888 175518 111897
rect 175462 111823 175518 111832
rect 116768 84856 116820 84862
rect 116768 84798 116820 84804
rect 116676 84244 116728 84250
rect 116676 84186 116728 84192
rect 116688 73778 116716 84186
rect 116676 73772 116728 73778
rect 116676 73714 116728 73720
rect 116676 72208 116728 72214
rect 116676 72150 116728 72156
rect 116584 70984 116636 70990
rect 116584 70926 116636 70932
rect 114468 22772 114520 22778
rect 114468 22714 114520 22720
rect 106292 16546 106504 16574
rect 113192 16546 114048 16574
rect 102140 10940 102192 10946
rect 102140 10882 102192 10888
rect 95792 10872 95844 10878
rect 95792 10814 95844 10820
rect 92480 10804 92532 10810
rect 92480 10746 92532 10752
rect 89166 10432 89222 10441
rect 89166 10367 89222 10376
rect 87970 7712 88026 7721
rect 87970 7647 88026 7656
rect 86224 6656 86276 6662
rect 86224 6598 86276 6604
rect 85672 5364 85724 5370
rect 85672 5306 85724 5312
rect 85684 480 85712 5306
rect 86868 5296 86920 5302
rect 86868 5238 86920 5244
rect 86880 480 86908 5238
rect 87984 480 88012 7647
rect 89180 480 89208 10367
rect 91558 7848 91614 7857
rect 91558 7783 91614 7792
rect 90362 4992 90418 5001
rect 90362 4927 90418 4936
rect 90376 480 90404 4927
rect 91572 480 91600 7783
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92492 354 92520 10746
rect 95148 8220 95200 8226
rect 95148 8162 95200 8168
rect 93952 5432 94004 5438
rect 93952 5374 94004 5380
rect 93964 480 93992 5374
rect 95160 480 95188 8162
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 95804 354 95832 10814
rect 98644 8288 98696 8294
rect 98644 8230 98696 8236
rect 97448 5500 97500 5506
rect 97448 5442 97500 5448
rect 97460 480 97488 5442
rect 98656 480 98684 8230
rect 99840 6792 99892 6798
rect 99840 6734 99892 6740
rect 99852 480 99880 6734
rect 101036 4140 101088 4146
rect 101036 4082 101088 4088
rect 101048 480 101076 4082
rect 102152 3398 102180 10882
rect 105726 9344 105782 9353
rect 105726 9279 105782 9288
rect 102232 7540 102284 7546
rect 102232 7482 102284 7488
rect 102140 3392 102192 3398
rect 102140 3334 102192 3340
rect 102244 480 102272 7482
rect 104532 6656 104584 6662
rect 104532 6598 104584 6604
rect 103336 3392 103388 3398
rect 103336 3334 103388 3340
rect 103348 480 103376 3334
rect 104544 480 104572 6598
rect 105740 480 105768 9279
rect 96222 354 96334 480
rect 95804 326 96334 354
rect 96222 -960 96334 326
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106476 354 106504 16546
rect 110512 11008 110564 11014
rect 110512 10950 110564 10956
rect 109314 9480 109370 9489
rect 109314 9415 109370 9424
rect 108118 6624 108174 6633
rect 108118 6559 108174 6568
rect 108132 480 108160 6559
rect 109328 480 109356 9415
rect 110524 480 110552 10950
rect 112812 9580 112864 9586
rect 112812 9522 112864 9528
rect 111616 4752 111668 4758
rect 111616 4694 111668 4700
rect 111628 480 111656 4694
rect 112824 480 112852 9522
rect 114020 480 114048 16546
rect 116400 9648 116452 9654
rect 116400 9590 116452 9596
rect 115204 6860 115256 6866
rect 115204 6802 115256 6808
rect 115216 480 115244 6802
rect 116412 480 116440 9590
rect 116688 9382 116716 72150
rect 116780 71126 116808 84798
rect 120356 75676 120408 75682
rect 120356 75618 120408 75624
rect 170404 75676 170456 75682
rect 170404 75618 170456 75624
rect 119344 72888 119396 72894
rect 119344 72830 119396 72836
rect 118148 72140 118200 72146
rect 118148 72082 118200 72088
rect 117964 72072 118016 72078
rect 117964 72014 118016 72020
rect 116768 71120 116820 71126
rect 116768 71062 116820 71068
rect 117320 10260 117372 10266
rect 117320 10202 117372 10208
rect 116676 9376 116728 9382
rect 116676 9318 116728 9324
rect 117228 4684 117280 4690
rect 117228 4626 117280 4632
rect 117240 4146 117268 4626
rect 117228 4140 117280 4146
rect 117228 4082 117280 4088
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117332 354 117360 10202
rect 117976 4962 118004 72014
rect 118056 72004 118108 72010
rect 118056 71946 118108 71952
rect 118068 7682 118096 71946
rect 118160 18630 118188 72082
rect 119356 54534 119384 72830
rect 120368 70922 120396 75618
rect 120908 73160 120960 73166
rect 120908 73102 120960 73108
rect 120724 73024 120776 73030
rect 120724 72966 120776 72972
rect 120356 70916 120408 70922
rect 120356 70858 120408 70864
rect 119344 54528 119396 54534
rect 119344 54470 119396 54476
rect 118148 18624 118200 18630
rect 118148 18566 118200 18572
rect 120632 10192 120684 10198
rect 120632 10134 120684 10140
rect 118056 7676 118108 7682
rect 118056 7618 118108 7624
rect 119896 7676 119948 7682
rect 119896 7618 119948 7624
rect 117964 4956 118016 4962
rect 117964 4898 118016 4904
rect 118792 4956 118844 4962
rect 118792 4898 118844 4904
rect 118804 480 118832 4898
rect 119908 480 119936 7618
rect 117566 354 117678 480
rect 117332 326 117678 354
rect 117566 -960 117678 326
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 120644 354 120672 10134
rect 120736 5370 120764 72966
rect 120816 72956 120868 72962
rect 120816 72898 120868 72904
rect 120828 6798 120856 72898
rect 120920 25566 120948 73102
rect 121092 72820 121144 72826
rect 121092 72762 121144 72768
rect 121000 72752 121052 72758
rect 121000 72694 121052 72700
rect 121012 43450 121040 72694
rect 121104 51134 121132 72762
rect 121368 72412 121420 72418
rect 121368 72354 121420 72360
rect 121092 51128 121144 51134
rect 121092 51070 121144 51076
rect 121000 43444 121052 43450
rect 121000 43386 121052 43392
rect 120908 25560 120960 25566
rect 120908 25502 120960 25508
rect 120816 6792 120868 6798
rect 120816 6734 120868 6740
rect 120724 5364 120776 5370
rect 120724 5306 120776 5312
rect 121380 4146 121408 72354
rect 121564 71913 121592 75140
rect 121656 72049 121684 75140
rect 121642 72040 121698 72049
rect 121642 71975 121698 71984
rect 121550 71904 121606 71913
rect 121550 71839 121606 71848
rect 121748 69850 121776 75140
rect 121656 69822 121776 69850
rect 121656 66910 121684 69822
rect 121736 69692 121788 69698
rect 121736 69634 121788 69640
rect 121644 66904 121696 66910
rect 121644 66846 121696 66852
rect 121748 6254 121776 69634
rect 121736 6248 121788 6254
rect 121736 6190 121788 6196
rect 121840 6186 121868 75140
rect 121932 72593 121960 75140
rect 121918 72584 121974 72593
rect 121918 72519 121974 72528
rect 121920 69896 121972 69902
rect 121920 69838 121972 69844
rect 121932 6322 121960 69838
rect 122024 67250 122052 75140
rect 122116 69630 122144 75140
rect 122208 69698 122236 75140
rect 122196 69692 122248 69698
rect 122196 69634 122248 69640
rect 122104 69624 122156 69630
rect 122104 69566 122156 69572
rect 122012 67244 122064 67250
rect 122012 67186 122064 67192
rect 122300 67130 122328 75140
rect 122392 72690 122420 75140
rect 122380 72684 122432 72690
rect 122380 72626 122432 72632
rect 122380 69828 122432 69834
rect 122380 69770 122432 69776
rect 122024 67102 122328 67130
rect 122024 8974 122052 67102
rect 122392 66994 122420 69770
rect 122484 69714 122512 75140
rect 122576 69902 122604 75140
rect 122564 69896 122616 69902
rect 122564 69838 122616 69844
rect 122668 69834 122696 75140
rect 122760 72894 122788 75140
rect 122748 72888 122800 72894
rect 122748 72830 122800 72836
rect 122748 72684 122800 72690
rect 122748 72626 122800 72632
rect 122656 69828 122708 69834
rect 122656 69770 122708 69776
rect 122484 69686 122696 69714
rect 122564 69624 122616 69630
rect 122564 69566 122616 69572
rect 122116 66966 122420 66994
rect 122116 13122 122144 66966
rect 122288 66904 122340 66910
rect 122288 66846 122340 66852
rect 122196 66836 122248 66842
rect 122196 66778 122248 66784
rect 122104 13116 122156 13122
rect 122104 13058 122156 13064
rect 122208 10742 122236 66778
rect 122196 10736 122248 10742
rect 122196 10678 122248 10684
rect 122012 8968 122064 8974
rect 122012 8910 122064 8916
rect 122300 6914 122328 66846
rect 122208 6886 122328 6914
rect 121920 6316 121972 6322
rect 121920 6258 121972 6264
rect 121828 6180 121880 6186
rect 121828 6122 121880 6128
rect 121368 4140 121420 4146
rect 121368 4082 121420 4088
rect 122208 3466 122236 6886
rect 122576 3534 122604 69566
rect 122668 3602 122696 69686
rect 122760 66842 122788 72626
rect 122852 72049 122880 75140
rect 122838 72040 122894 72049
rect 122838 71975 122894 71984
rect 122944 71913 122972 75140
rect 123036 72010 123064 75140
rect 123128 72486 123156 75140
rect 123116 72480 123168 72486
rect 123116 72422 123168 72428
rect 123024 72004 123076 72010
rect 123024 71946 123076 71952
rect 122930 71904 122986 71913
rect 122930 71839 122986 71848
rect 123024 69964 123076 69970
rect 123024 69906 123076 69912
rect 122932 69828 122984 69834
rect 122932 69770 122984 69776
rect 122748 66836 122800 66842
rect 122748 66778 122800 66784
rect 122944 5030 122972 69770
rect 122932 5024 122984 5030
rect 122932 4966 122984 4972
rect 123036 4894 123064 69906
rect 123116 69760 123168 69766
rect 123116 69702 123168 69708
rect 123128 6390 123156 69702
rect 123220 69698 123248 75140
rect 123208 69692 123260 69698
rect 123208 69634 123260 69640
rect 123312 67946 123340 75140
rect 123404 69714 123432 75140
rect 123496 69816 123524 75140
rect 123588 69970 123616 75140
rect 123576 69964 123628 69970
rect 123576 69906 123628 69912
rect 123496 69788 123616 69816
rect 123404 69686 123524 69714
rect 123392 69624 123444 69630
rect 123392 69566 123444 69572
rect 123220 67918 123340 67946
rect 123220 7614 123248 67918
rect 123300 67856 123352 67862
rect 123300 67798 123352 67804
rect 123312 7750 123340 67798
rect 123404 9110 123432 69566
rect 123392 9104 123444 9110
rect 123392 9046 123444 9052
rect 123496 9042 123524 69686
rect 123588 10334 123616 69788
rect 123680 67862 123708 75140
rect 123772 72078 123800 75140
rect 123760 72072 123812 72078
rect 123760 72014 123812 72020
rect 123864 69766 123892 75140
rect 123852 69760 123904 69766
rect 123852 69702 123904 69708
rect 123760 69692 123812 69698
rect 123760 69634 123812 69640
rect 123668 67856 123720 67862
rect 123668 67798 123720 67804
rect 123668 67720 123720 67726
rect 123668 67662 123720 67668
rect 123680 10402 123708 67662
rect 123668 10396 123720 10402
rect 123668 10338 123720 10344
rect 123576 10328 123628 10334
rect 123576 10270 123628 10276
rect 123484 9036 123536 9042
rect 123484 8978 123536 8984
rect 123300 7744 123352 7750
rect 123300 7686 123352 7692
rect 123208 7608 123260 7614
rect 123208 7550 123260 7556
rect 123116 6384 123168 6390
rect 123116 6326 123168 6332
rect 123024 4888 123076 4894
rect 123024 4830 123076 4836
rect 123772 4826 123800 69634
rect 123956 69630 123984 75140
rect 123944 69624 123996 69630
rect 123944 69566 123996 69572
rect 124048 67726 124076 75140
rect 124140 69834 124168 75140
rect 124232 72185 124260 75140
rect 124218 72176 124274 72185
rect 124324 72146 124352 75140
rect 124218 72111 124274 72120
rect 124312 72140 124364 72146
rect 124312 72082 124364 72088
rect 124416 72049 124444 75140
rect 124402 72040 124458 72049
rect 124402 71975 124458 71984
rect 124508 71913 124536 75140
rect 124494 71904 124550 71913
rect 124494 71839 124550 71848
rect 124128 69828 124180 69834
rect 124128 69770 124180 69776
rect 124600 69714 124628 75140
rect 124324 69686 124628 69714
rect 124036 67720 124088 67726
rect 124036 67662 124088 67668
rect 123760 4820 123812 4826
rect 123760 4762 123812 4768
rect 124324 3670 124352 69686
rect 124588 69624 124640 69630
rect 124588 69566 124640 69572
rect 124496 69556 124548 69562
rect 124496 69498 124548 69504
rect 124508 6594 124536 69498
rect 124496 6588 124548 6594
rect 124496 6530 124548 6536
rect 124600 6526 124628 69566
rect 124588 6520 124640 6526
rect 124588 6462 124640 6468
rect 124692 6458 124720 75140
rect 124784 69578 124812 75140
rect 124876 72214 124904 75140
rect 124864 72208 124916 72214
rect 124864 72150 124916 72156
rect 124968 69834 124996 75140
rect 124956 69828 125008 69834
rect 124956 69770 125008 69776
rect 124784 69550 124996 69578
rect 124864 69488 124916 69494
rect 124864 69430 124916 69436
rect 124772 66224 124824 66230
rect 124772 66166 124824 66172
rect 124784 9246 124812 66166
rect 124876 9314 124904 69430
rect 124864 9308 124916 9314
rect 124864 9250 124916 9256
rect 124772 9240 124824 9246
rect 124772 9182 124824 9188
rect 124968 9178 124996 69550
rect 125060 66230 125088 75140
rect 125048 66224 125100 66230
rect 125048 66166 125100 66172
rect 125152 64874 125180 75140
rect 125060 64846 125180 64874
rect 125244 64874 125272 75140
rect 125336 69562 125364 75140
rect 125324 69556 125376 69562
rect 125324 69498 125376 69504
rect 125428 69494 125456 75140
rect 125416 69488 125468 69494
rect 125416 69430 125468 69436
rect 125244 64846 125364 64874
rect 125060 10470 125088 64846
rect 125048 10464 125100 10470
rect 125048 10406 125100 10412
rect 124956 9172 125008 9178
rect 124956 9114 125008 9120
rect 124680 6452 124732 6458
rect 124680 6394 124732 6400
rect 125336 3738 125364 64846
rect 125520 3806 125548 75140
rect 125612 72049 125640 75140
rect 125704 72321 125732 75140
rect 125690 72312 125746 72321
rect 125690 72247 125746 72256
rect 125796 72185 125824 75140
rect 125782 72176 125838 72185
rect 125782 72111 125838 72120
rect 125598 72040 125654 72049
rect 125598 71975 125654 71984
rect 125888 71913 125916 75140
rect 125874 71904 125930 71913
rect 125874 71839 125930 71848
rect 125784 69896 125836 69902
rect 125784 69838 125836 69844
rect 125692 69624 125744 69630
rect 125692 69566 125744 69572
rect 125704 3942 125732 69566
rect 125796 5098 125824 69838
rect 125980 67862 126008 75140
rect 126072 69766 126100 75140
rect 126060 69760 126112 69766
rect 126060 69702 126112 69708
rect 126164 68082 126192 75140
rect 126072 68054 126192 68082
rect 125968 67856 126020 67862
rect 125968 67798 126020 67804
rect 126072 67674 126100 68054
rect 126256 67946 126284 75140
rect 126348 72554 126376 75140
rect 126336 72548 126388 72554
rect 126336 72490 126388 72496
rect 126336 69692 126388 69698
rect 126336 69634 126388 69640
rect 125888 67646 126100 67674
rect 126164 67918 126284 67946
rect 125888 6730 125916 67646
rect 126060 67584 126112 67590
rect 126060 67526 126112 67532
rect 125968 67516 126020 67522
rect 125968 67458 126020 67464
rect 125980 7886 126008 67458
rect 125968 7880 126020 7886
rect 125968 7822 126020 7828
rect 126072 7818 126100 67526
rect 126164 9518 126192 67918
rect 126244 67856 126296 67862
rect 126244 67798 126296 67804
rect 126152 9512 126204 9518
rect 126152 9454 126204 9460
rect 126256 9450 126284 67798
rect 126348 10606 126376 69634
rect 126440 67590 126468 75140
rect 126428 67584 126480 67590
rect 126428 67526 126480 67532
rect 126532 64874 126560 75140
rect 126624 69902 126652 75140
rect 126612 69896 126664 69902
rect 126612 69838 126664 69844
rect 126612 69760 126664 69766
rect 126612 69702 126664 69708
rect 126440 64846 126560 64874
rect 126336 10600 126388 10606
rect 126336 10542 126388 10548
rect 126440 10538 126468 64846
rect 126428 10532 126480 10538
rect 126428 10474 126480 10480
rect 126244 9444 126296 9450
rect 126244 9386 126296 9392
rect 126060 7812 126112 7818
rect 126060 7754 126112 7760
rect 125876 6724 125928 6730
rect 125876 6666 125928 6672
rect 125784 5092 125836 5098
rect 125784 5034 125836 5040
rect 125692 3936 125744 3942
rect 125692 3878 125744 3884
rect 126624 3874 126652 69702
rect 126716 67522 126744 75140
rect 126808 69698 126836 75140
rect 126796 69692 126848 69698
rect 126796 69634 126848 69640
rect 126900 69630 126928 75140
rect 126992 71913 127020 75140
rect 127084 72049 127112 75140
rect 127070 72040 127126 72049
rect 127070 71975 127126 71984
rect 126978 71904 127034 71913
rect 126978 71839 127034 71848
rect 126888 69624 126940 69630
rect 126888 69566 126940 69572
rect 126704 67516 126756 67522
rect 126704 67458 126756 67464
rect 127176 5166 127204 75140
rect 127268 68082 127296 75140
rect 127360 72690 127388 75140
rect 127348 72684 127400 72690
rect 127348 72626 127400 72632
rect 127452 68202 127480 75140
rect 127544 69714 127572 75140
rect 127636 71754 127664 75140
rect 127728 71874 127756 75140
rect 127820 71890 127848 75140
rect 127912 73166 127940 75140
rect 127900 73160 127952 73166
rect 127900 73102 127952 73108
rect 127716 71868 127768 71874
rect 127820 71862 127940 71890
rect 127716 71810 127768 71816
rect 127636 71726 127848 71754
rect 127624 71596 127676 71602
rect 127624 71538 127676 71544
rect 127636 70990 127664 71538
rect 127624 70984 127676 70990
rect 127624 70926 127676 70932
rect 127544 69686 127664 69714
rect 127440 68196 127492 68202
rect 127440 68138 127492 68144
rect 127268 68054 127480 68082
rect 127452 67946 127480 68054
rect 127348 67924 127400 67930
rect 127452 67918 127572 67946
rect 127348 67866 127400 67872
rect 127256 67788 127308 67794
rect 127256 67730 127308 67736
rect 127268 5302 127296 67730
rect 127256 5296 127308 5302
rect 127256 5238 127308 5244
rect 127360 5234 127388 67866
rect 127440 67856 127492 67862
rect 127440 67798 127492 67804
rect 127452 8090 127480 67798
rect 127440 8084 127492 8090
rect 127440 8026 127492 8032
rect 127544 7954 127572 67918
rect 127636 8022 127664 69686
rect 127716 69692 127768 69698
rect 127716 69634 127768 69640
rect 127728 8158 127756 69634
rect 127820 10674 127848 71726
rect 127912 67862 127940 71862
rect 127900 67856 127952 67862
rect 127900 67798 127952 67804
rect 127808 10668 127860 10674
rect 127808 10610 127860 10616
rect 127716 8152 127768 8158
rect 127716 8094 127768 8100
rect 127624 8016 127676 8022
rect 127624 7958 127676 7964
rect 127532 7948 127584 7954
rect 127532 7890 127584 7896
rect 127348 5228 127400 5234
rect 127348 5170 127400 5176
rect 127164 5160 127216 5166
rect 127164 5102 127216 5108
rect 128004 4078 128032 75140
rect 128096 72026 128124 75140
rect 128188 73030 128216 75140
rect 128176 73024 128228 73030
rect 128176 72966 128228 72972
rect 128096 71998 128216 72026
rect 128084 71868 128136 71874
rect 128084 71810 128136 71816
rect 127992 4072 128044 4078
rect 127992 4014 128044 4020
rect 128096 4010 128124 71810
rect 128188 69698 128216 71998
rect 128176 69692 128228 69698
rect 128176 69634 128228 69640
rect 128280 67794 128308 75140
rect 128372 72049 128400 75140
rect 128464 72185 128492 75140
rect 128556 73137 128584 75140
rect 128542 73128 128598 73137
rect 128542 73063 128598 73072
rect 128450 72176 128506 72185
rect 128450 72111 128506 72120
rect 128358 72040 128414 72049
rect 128358 71975 128414 71984
rect 128648 71913 128676 75140
rect 128634 71904 128690 71913
rect 128634 71839 128690 71848
rect 128544 69692 128596 69698
rect 128544 69634 128596 69640
rect 128268 67788 128320 67794
rect 128268 67730 128320 67736
rect 128556 5438 128584 69634
rect 128636 69624 128688 69630
rect 128636 69566 128688 69572
rect 128648 6662 128676 69566
rect 128740 67862 128768 75140
rect 128832 69698 128860 75140
rect 128820 69692 128872 69698
rect 128820 69634 128872 69640
rect 128924 68082 128952 75140
rect 129016 69698 129044 75140
rect 129108 69970 129136 75140
rect 129096 69964 129148 69970
rect 129096 69906 129148 69912
rect 129200 69816 129228 75140
rect 129292 72962 129320 75140
rect 129280 72956 129332 72962
rect 129280 72898 129332 72904
rect 129108 69788 129228 69816
rect 129004 69692 129056 69698
rect 129004 69634 129056 69640
rect 128832 68054 128952 68082
rect 128728 67856 128780 67862
rect 128728 67798 128780 67804
rect 128728 67720 128780 67726
rect 128728 67662 128780 67668
rect 128740 7546 128768 67662
rect 128832 8226 128860 68054
rect 129108 67946 129136 69788
rect 129188 69692 129240 69698
rect 129188 69634 129240 69640
rect 128924 67918 129136 67946
rect 128924 8294 128952 67918
rect 129096 67856 129148 67862
rect 129096 67798 129148 67804
rect 129004 67788 129056 67794
rect 129004 67730 129056 67736
rect 129016 10946 129044 67730
rect 129004 10940 129056 10946
rect 129004 10882 129056 10888
rect 129108 10810 129136 67798
rect 129200 10878 129228 69634
rect 129188 10872 129240 10878
rect 129188 10814 129240 10820
rect 129096 10804 129148 10810
rect 129096 10746 129148 10752
rect 128912 8288 128964 8294
rect 128912 8230 128964 8236
rect 128820 8220 128872 8226
rect 128820 8162 128872 8168
rect 128728 7540 128780 7546
rect 128728 7482 128780 7488
rect 128636 6656 128688 6662
rect 128636 6598 128688 6604
rect 128544 5432 128596 5438
rect 128544 5374 128596 5380
rect 129384 4690 129412 75140
rect 129476 67726 129504 75140
rect 129568 67794 129596 75140
rect 129660 70122 129688 75140
rect 129752 72185 129780 75140
rect 129844 72758 129872 75140
rect 129832 72752 129884 72758
rect 129832 72694 129884 72700
rect 129738 72176 129794 72185
rect 129738 72111 129794 72120
rect 129936 71913 129964 75140
rect 130028 72049 130056 75140
rect 130014 72040 130070 72049
rect 130014 71975 130070 71984
rect 129922 71904 129978 71913
rect 129922 71839 129978 71848
rect 129660 70094 129780 70122
rect 129648 69964 129700 69970
rect 129648 69906 129700 69912
rect 129556 67788 129608 67794
rect 129556 67730 129608 67736
rect 129464 67720 129516 67726
rect 129464 67662 129516 67668
rect 129660 5506 129688 69906
rect 129752 69630 129780 70094
rect 130120 69834 130148 75140
rect 130108 69828 130160 69834
rect 130108 69770 130160 69776
rect 130212 69714 130240 75140
rect 129936 69686 130240 69714
rect 129740 69624 129792 69630
rect 129740 69566 129792 69572
rect 129648 5500 129700 5506
rect 129648 5442 129700 5448
rect 129936 4758 129964 69686
rect 130016 69624 130068 69630
rect 130016 69566 130068 69572
rect 130200 69624 130252 69630
rect 130200 69566 130252 69572
rect 130028 6866 130056 69566
rect 130108 69488 130160 69494
rect 130108 69430 130160 69436
rect 130120 7682 130148 69430
rect 130212 9654 130240 69566
rect 130200 9648 130252 9654
rect 130200 9590 130252 9596
rect 130304 9586 130332 75140
rect 130396 72826 130424 75140
rect 130384 72820 130436 72826
rect 130384 72762 130436 72768
rect 130488 69902 130516 75140
rect 130476 69896 130528 69902
rect 130476 69838 130528 69844
rect 130580 69834 130608 75140
rect 130568 69828 130620 69834
rect 130568 69770 130620 69776
rect 130672 69714 130700 75140
rect 130396 69686 130700 69714
rect 130396 10266 130424 69686
rect 130568 69624 130620 69630
rect 130568 69566 130620 69572
rect 130476 69556 130528 69562
rect 130476 69498 130528 69504
rect 130488 11014 130516 69498
rect 130476 11008 130528 11014
rect 130476 10950 130528 10956
rect 130384 10260 130436 10266
rect 130384 10202 130436 10208
rect 130580 10198 130608 69566
rect 130764 64874 130792 75140
rect 130856 69494 130884 75140
rect 130948 69630 130976 75140
rect 130936 69624 130988 69630
rect 130936 69566 130988 69572
rect 130844 69488 130896 69494
rect 130844 69430 130896 69436
rect 130764 64846 130884 64874
rect 130568 10192 130620 10198
rect 130568 10134 130620 10140
rect 130292 9580 130344 9586
rect 130292 9522 130344 9528
rect 130108 7676 130160 7682
rect 130108 7618 130160 7624
rect 130016 6860 130068 6866
rect 130016 6802 130068 6808
rect 130856 4962 130884 64846
rect 130844 4956 130896 4962
rect 130844 4898 130896 4904
rect 129924 4752 129976 4758
rect 129924 4694 129976 4700
rect 129372 4684 129424 4690
rect 129372 4626 129424 4632
rect 128084 4004 128136 4010
rect 128084 3946 128136 3952
rect 126612 3868 126664 3874
rect 126612 3810 126664 3816
rect 125508 3800 125560 3806
rect 125508 3742 125560 3748
rect 125324 3732 125376 3738
rect 125324 3674 125376 3680
rect 124312 3664 124364 3670
rect 123482 3632 123538 3641
rect 122656 3596 122708 3602
rect 124312 3606 124364 3612
rect 123482 3567 123538 3576
rect 122656 3538 122708 3544
rect 122564 3528 122616 3534
rect 122564 3470 122616 3476
rect 122196 3460 122248 3466
rect 122196 3402 122248 3408
rect 122288 3392 122340 3398
rect 122288 3334 122340 3340
rect 122300 480 122328 3334
rect 123496 480 123524 3567
rect 125876 3528 125928 3534
rect 124678 3496 124734 3505
rect 125876 3470 125928 3476
rect 124678 3431 124734 3440
rect 124692 480 124720 3431
rect 125888 480 125916 3470
rect 126980 3460 127032 3466
rect 126980 3402 127032 3408
rect 126992 480 127020 3402
rect 131040 3398 131068 75140
rect 131132 71913 131160 75140
rect 131224 72049 131252 75140
rect 131210 72040 131266 72049
rect 131210 71975 131266 71984
rect 131118 71904 131174 71913
rect 131118 71839 131174 71848
rect 131316 68082 131344 75140
rect 131408 73302 131436 75140
rect 131396 73296 131448 73302
rect 131396 73238 131448 73244
rect 131396 73160 131448 73166
rect 131396 73102 131448 73108
rect 131408 68338 131436 73102
rect 131396 68332 131448 68338
rect 131396 68274 131448 68280
rect 131500 68218 131528 75140
rect 131224 68054 131344 68082
rect 131408 68190 131528 68218
rect 131224 3534 131252 68054
rect 131304 67992 131356 67998
rect 131304 67934 131356 67940
rect 131212 3528 131264 3534
rect 131212 3470 131264 3476
rect 131028 3392 131080 3398
rect 131028 3334 131080 3340
rect 128176 3120 128228 3126
rect 128176 3062 128228 3068
rect 128188 480 128216 3062
rect 129372 3052 129424 3058
rect 129372 2994 129424 3000
rect 129384 480 129412 2994
rect 131316 2802 131344 67934
rect 131408 3126 131436 68190
rect 131592 67946 131620 75140
rect 131684 73438 131712 75140
rect 131672 73432 131724 73438
rect 131672 73374 131724 73380
rect 131672 73296 131724 73302
rect 131672 73238 131724 73244
rect 131500 67918 131620 67946
rect 131396 3120 131448 3126
rect 131396 3062 131448 3068
rect 131500 3058 131528 67918
rect 131684 64874 131712 73238
rect 131592 64846 131712 64874
rect 131592 3466 131620 64846
rect 131580 3460 131632 3466
rect 131580 3402 131632 3408
rect 131488 3052 131540 3058
rect 131488 2994 131540 3000
rect 131040 2774 131344 2802
rect 121062 354 121174 480
rect 120644 326 121174 354
rect 121062 -960 121174 326
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 354 130650 480
rect 131040 354 131068 2774
rect 131776 480 131804 75140
rect 131868 4078 131896 75140
rect 131856 4072 131908 4078
rect 131856 4014 131908 4020
rect 131960 3398 131988 75140
rect 132052 3942 132080 75140
rect 132040 3936 132092 3942
rect 132040 3878 132092 3884
rect 131948 3392 132000 3398
rect 131948 3334 132000 3340
rect 132144 3330 132172 75140
rect 132236 72049 132264 75140
rect 132328 72690 132356 75140
rect 132316 72684 132368 72690
rect 132316 72626 132368 72632
rect 132222 72040 132278 72049
rect 132222 71975 132278 71984
rect 132420 71913 132448 75140
rect 132406 71904 132462 71913
rect 132406 71839 132462 71848
rect 132512 71806 132540 75140
rect 132500 71800 132552 71806
rect 132500 71742 132552 71748
rect 132604 5438 132632 75140
rect 132696 72622 132724 75140
rect 132684 72616 132736 72622
rect 132684 72558 132736 72564
rect 132592 5432 132644 5438
rect 132592 5374 132644 5380
rect 132788 5370 132816 75140
rect 132776 5364 132828 5370
rect 132776 5306 132828 5312
rect 132880 4010 132908 75140
rect 132972 4978 133000 75140
rect 133064 5166 133092 75140
rect 133052 5160 133104 5166
rect 133052 5102 133104 5108
rect 133156 5098 133184 75140
rect 133144 5092 133196 5098
rect 133144 5034 133196 5040
rect 132972 4950 133092 4978
rect 132960 4072 133012 4078
rect 132960 4014 133012 4020
rect 132868 4004 132920 4010
rect 132868 3946 132920 3952
rect 132132 3324 132184 3330
rect 132132 3266 132184 3272
rect 132972 480 133000 4014
rect 133064 3602 133092 4950
rect 133052 3596 133104 3602
rect 133052 3538 133104 3544
rect 133248 3534 133276 75140
rect 133340 4962 133368 75140
rect 133432 5030 133460 75140
rect 133420 5024 133472 5030
rect 133420 4966 133472 4972
rect 133328 4956 133380 4962
rect 133328 4898 133380 4904
rect 133236 3528 133288 3534
rect 133236 3470 133288 3476
rect 133524 3466 133552 75140
rect 133616 72185 133644 75140
rect 133602 72176 133658 72185
rect 133602 72111 133658 72120
rect 133708 72049 133736 75140
rect 133694 72040 133750 72049
rect 133694 71975 133750 71984
rect 133800 71913 133828 75140
rect 133786 71904 133842 71913
rect 133786 71839 133842 71848
rect 133892 4894 133920 75140
rect 133984 72350 134012 75140
rect 133972 72344 134024 72350
rect 133972 72286 134024 72292
rect 133880 4888 133932 4894
rect 133880 4830 133932 4836
rect 134076 4010 134104 75140
rect 134064 4004 134116 4010
rect 134064 3946 134116 3952
rect 134168 3874 134196 75140
rect 134260 4826 134288 75140
rect 134248 4820 134300 4826
rect 134248 4762 134300 4768
rect 134156 3868 134208 3874
rect 134156 3810 134208 3816
rect 134352 3806 134380 75140
rect 134340 3800 134392 3806
rect 134340 3742 134392 3748
rect 134444 3738 134472 75140
rect 134536 5302 134564 75140
rect 134524 5296 134576 5302
rect 134524 5238 134576 5244
rect 134432 3732 134484 3738
rect 134432 3674 134484 3680
rect 134628 3670 134656 75140
rect 134720 72554 134748 75140
rect 134708 72548 134760 72554
rect 134708 72490 134760 72496
rect 134812 10878 134840 75140
rect 134800 10872 134852 10878
rect 134800 10814 134852 10820
rect 134904 8906 134932 75140
rect 134996 72049 135024 75140
rect 135088 72185 135116 75140
rect 135074 72176 135130 72185
rect 135074 72111 135130 72120
rect 134982 72040 135038 72049
rect 134982 71975 135038 71984
rect 135180 71913 135208 75140
rect 135166 71904 135222 71913
rect 135166 71839 135222 71848
rect 135272 25430 135300 75140
rect 135364 32978 135392 75140
rect 135352 32972 135404 32978
rect 135352 32914 135404 32920
rect 135260 25424 135312 25430
rect 135260 25366 135312 25372
rect 135456 9654 135484 75140
rect 135548 25498 135576 75140
rect 135640 32910 135668 75140
rect 135732 72486 135760 75140
rect 135720 72480 135772 72486
rect 135720 72422 135772 72428
rect 135628 32904 135680 32910
rect 135628 32846 135680 32852
rect 135824 26246 135852 75140
rect 135916 32842 135944 75140
rect 135904 32836 135956 32842
rect 135904 32778 135956 32784
rect 135812 26240 135864 26246
rect 135812 26182 135864 26188
rect 135536 25492 135588 25498
rect 135536 25434 135588 25440
rect 135444 9648 135496 9654
rect 135444 9590 135496 9596
rect 136008 9586 136036 75140
rect 136100 27538 136128 75140
rect 136192 71913 136220 75140
rect 136284 72962 136312 75140
rect 136272 72956 136324 72962
rect 136272 72898 136324 72904
rect 136376 72049 136404 75140
rect 136468 72185 136496 75140
rect 136454 72176 136510 72185
rect 136454 72111 136510 72120
rect 136362 72040 136418 72049
rect 136362 71975 136418 71984
rect 136560 71913 136588 75140
rect 136178 71904 136234 71913
rect 136178 71839 136234 71848
rect 136546 71904 136602 71913
rect 136546 71839 136602 71848
rect 136652 71806 136680 75140
rect 136180 71800 136232 71806
rect 136180 71742 136232 71748
rect 136640 71800 136692 71806
rect 136640 71742 136692 71748
rect 136088 27532 136140 27538
rect 136088 27474 136140 27480
rect 135996 9580 136048 9586
rect 135996 9522 136048 9528
rect 134892 8900 134944 8906
rect 134892 8842 134944 8848
rect 135260 3936 135312 3942
rect 135260 3878 135312 3884
rect 134616 3664 134668 3670
rect 134616 3606 134668 3612
rect 133512 3460 133564 3466
rect 133512 3402 133564 3408
rect 134156 3392 134208 3398
rect 134156 3334 134208 3340
rect 134168 480 134196 3334
rect 135272 480 135300 3878
rect 136192 2990 136220 71742
rect 136744 32774 136772 75140
rect 136836 73166 136864 75140
rect 136824 73160 136876 73166
rect 136824 73102 136876 73108
rect 136732 32768 136784 32774
rect 136732 32710 136784 32716
rect 136928 27470 136956 75140
rect 137020 32706 137048 75140
rect 137008 32700 137060 32706
rect 137008 32642 137060 32648
rect 136916 27464 136968 27470
rect 136916 27406 136968 27412
rect 137112 10810 137140 75140
rect 137204 27334 137232 75140
rect 137192 27328 137244 27334
rect 137192 27270 137244 27276
rect 137100 10804 137152 10810
rect 137100 10746 137152 10752
rect 137296 5234 137324 75140
rect 137388 10742 137416 75140
rect 137480 27266 137508 75140
rect 137572 32638 137600 75140
rect 137664 73098 137692 75140
rect 137652 73092 137704 73098
rect 137652 73034 137704 73040
rect 137756 73030 137784 75140
rect 137744 73024 137796 73030
rect 137744 72966 137796 72972
rect 137744 72684 137796 72690
rect 137744 72626 137796 72632
rect 137652 72344 137704 72350
rect 137652 72286 137704 72292
rect 137560 32632 137612 32638
rect 137560 32574 137612 32580
rect 137468 27260 137520 27266
rect 137468 27202 137520 27208
rect 137664 16574 137692 72286
rect 137756 69578 137784 72626
rect 137848 72049 137876 75140
rect 137834 72040 137890 72049
rect 137834 71975 137890 71984
rect 137940 71913 137968 75140
rect 137926 71904 137982 71913
rect 137926 71839 137982 71848
rect 138032 69714 138060 75140
rect 138124 69834 138152 75140
rect 138112 69828 138164 69834
rect 138112 69770 138164 69776
rect 138032 69686 138152 69714
rect 137756 69550 138060 69578
rect 137664 16546 137784 16574
rect 137376 10736 137428 10742
rect 137376 10678 137428 10684
rect 137284 5228 137336 5234
rect 137284 5170 137336 5176
rect 137650 3632 137706 3641
rect 137650 3567 137706 3576
rect 136456 3324 136508 3330
rect 136456 3266 136508 3272
rect 136180 2984 136232 2990
rect 136180 2926 136232 2932
rect 136468 480 136496 3266
rect 137664 480 137692 3567
rect 137756 3398 137784 16546
rect 138032 6914 138060 69550
rect 138124 28150 138152 69686
rect 138112 28144 138164 28150
rect 138112 28086 138164 28092
rect 138216 12238 138244 75140
rect 138308 28218 138336 75140
rect 138400 34406 138428 75140
rect 138388 34400 138440 34406
rect 138388 34342 138440 34348
rect 138296 28212 138348 28218
rect 138296 28154 138348 28160
rect 138204 12232 138256 12238
rect 138204 12174 138256 12180
rect 138492 12170 138520 75140
rect 138584 27198 138612 75140
rect 138676 69850 138704 75140
rect 138768 69970 138796 75140
rect 138860 72690 138888 75140
rect 138848 72684 138900 72690
rect 138848 72626 138900 72632
rect 138952 71913 138980 75140
rect 139044 72049 139072 75140
rect 139030 72040 139086 72049
rect 139030 71975 139086 71984
rect 139136 71913 139164 75140
rect 139228 72622 139256 75140
rect 139216 72616 139268 72622
rect 139216 72558 139268 72564
rect 139320 72185 139348 75140
rect 139306 72176 139362 72185
rect 139306 72111 139362 72120
rect 138938 71904 138994 71913
rect 138938 71839 138994 71848
rect 139122 71904 139178 71913
rect 139122 71839 139178 71848
rect 138756 69964 138808 69970
rect 138756 69906 138808 69912
rect 138676 69822 138888 69850
rect 138756 69692 138808 69698
rect 138756 69634 138808 69640
rect 138664 69624 138716 69630
rect 138664 69566 138716 69572
rect 138676 34474 138704 69566
rect 138664 34468 138716 34474
rect 138664 34410 138716 34416
rect 138572 27192 138624 27198
rect 138572 27134 138624 27140
rect 138480 12164 138532 12170
rect 138480 12106 138532 12112
rect 138768 12102 138796 69634
rect 138860 34338 138888 69822
rect 138848 34332 138900 34338
rect 138848 34274 138900 34280
rect 139412 28966 139440 75140
rect 139400 28960 139452 28966
rect 139400 28902 139452 28908
rect 139504 20262 139532 75140
rect 139492 20256 139544 20262
rect 139492 20198 139544 20204
rect 139596 13462 139624 75140
rect 139688 27130 139716 75140
rect 139780 34270 139808 75140
rect 139768 34264 139820 34270
rect 139768 34206 139820 34212
rect 139676 27124 139728 27130
rect 139676 27066 139728 27072
rect 139584 13456 139636 13462
rect 139584 13398 139636 13404
rect 138756 12096 138808 12102
rect 138756 12038 138808 12044
rect 138032 6886 138888 6914
rect 137744 3392 137796 3398
rect 137744 3334 137796 3340
rect 138860 480 138888 6886
rect 139872 6730 139900 75140
rect 139964 26178 139992 75140
rect 139952 26172 140004 26178
rect 139952 26114 140004 26120
rect 140056 20466 140084 75140
rect 140044 20460 140096 20466
rect 140044 20402 140096 20408
rect 140148 13394 140176 75140
rect 140240 28830 140268 75140
rect 140332 72185 140360 75140
rect 140318 72176 140374 72185
rect 140318 72111 140374 72120
rect 140424 71913 140452 75140
rect 140516 72758 140544 75140
rect 140504 72752 140556 72758
rect 140504 72694 140556 72700
rect 140608 72049 140636 75140
rect 140594 72040 140650 72049
rect 140594 71975 140650 71984
rect 140700 71913 140728 75140
rect 140410 71904 140466 71913
rect 140410 71839 140466 71848
rect 140686 71904 140742 71913
rect 140686 71839 140742 71848
rect 140228 28824 140280 28830
rect 140228 28766 140280 28772
rect 140792 28762 140820 75140
rect 140884 34202 140912 75140
rect 140976 74866 141004 75140
rect 140964 74860 141016 74866
rect 140964 74802 141016 74808
rect 140872 34196 140924 34202
rect 140872 34138 140924 34144
rect 140780 28756 140832 28762
rect 140780 28698 140832 28704
rect 141068 28626 141096 75140
rect 141056 28620 141108 28626
rect 141056 28562 141108 28568
rect 141160 19106 141188 75140
rect 141148 19100 141200 19106
rect 141148 19042 141200 19048
rect 141252 14958 141280 75140
rect 141344 24818 141372 75140
rect 141436 34134 141464 75140
rect 141424 34128 141476 34134
rect 141424 34070 141476 34076
rect 141332 24812 141384 24818
rect 141332 24754 141384 24760
rect 141240 14952 141292 14958
rect 141240 14894 141292 14900
rect 141528 14890 141556 75140
rect 141620 72894 141648 75140
rect 141608 72888 141660 72894
rect 141608 72830 141660 72836
rect 141712 20398 141740 75140
rect 141804 74934 141832 75140
rect 141792 74928 141844 74934
rect 141792 74870 141844 74876
rect 141896 26110 141924 75140
rect 141988 72049 142016 75140
rect 141974 72040 142030 72049
rect 141974 71975 142030 71984
rect 142080 71913 142108 75140
rect 142172 72418 142200 75140
rect 142160 72412 142212 72418
rect 142160 72354 142212 72360
rect 142066 71904 142122 71913
rect 142066 71839 142122 71848
rect 142264 32570 142292 75140
rect 142252 32564 142304 32570
rect 142252 32506 142304 32512
rect 141884 26104 141936 26110
rect 141884 26046 141936 26052
rect 141700 20392 141752 20398
rect 141700 20334 141752 20340
rect 141516 14884 141568 14890
rect 141516 14826 141568 14832
rect 142356 14822 142384 75140
rect 142344 14816 142396 14822
rect 142344 14758 142396 14764
rect 140136 13388 140188 13394
rect 140136 13330 140188 13336
rect 142448 8022 142476 75140
rect 142540 34066 142568 75140
rect 142528 34060 142580 34066
rect 142528 34002 142580 34008
rect 142632 14754 142660 75140
rect 142724 72826 142752 75140
rect 142712 72820 142764 72826
rect 142712 72762 142764 72768
rect 142712 72684 142764 72690
rect 142712 72626 142764 72632
rect 142724 72214 142752 72626
rect 142712 72208 142764 72214
rect 142712 72150 142764 72156
rect 142816 17678 142844 75140
rect 142804 17672 142856 17678
rect 142804 17614 142856 17620
rect 142908 16454 142936 75140
rect 142896 16448 142948 16454
rect 142896 16390 142948 16396
rect 142620 14748 142672 14754
rect 142620 14690 142672 14696
rect 143000 10674 143028 75140
rect 143092 33998 143120 75140
rect 143184 71913 143212 75140
rect 143276 72321 143304 75140
rect 143262 72312 143318 72321
rect 143262 72247 143318 72256
rect 143368 72185 143396 75140
rect 143354 72176 143410 72185
rect 143354 72111 143410 72120
rect 143460 72049 143488 75140
rect 143446 72040 143502 72049
rect 143446 71975 143502 71984
rect 143170 71904 143226 71913
rect 143170 71839 143226 71848
rect 143264 71800 143316 71806
rect 143264 71742 143316 71748
rect 143080 33992 143132 33998
rect 143080 33934 143132 33940
rect 143276 27606 143304 71742
rect 143264 27600 143316 27606
rect 143264 27542 143316 27548
rect 143552 24750 143580 75140
rect 143644 33930 143672 75140
rect 143736 74322 143764 75140
rect 143724 74316 143776 74322
rect 143724 74258 143776 74264
rect 143632 33924 143684 33930
rect 143632 33866 143684 33872
rect 143540 24744 143592 24750
rect 143540 24686 143592 24692
rect 142988 10668 143040 10674
rect 142988 10610 143040 10616
rect 142436 8016 142488 8022
rect 142436 7958 142488 7964
rect 139860 6724 139912 6730
rect 139860 6666 139912 6672
rect 143828 6662 143856 75140
rect 143920 16386 143948 75140
rect 143908 16380 143960 16386
rect 143908 16322 143960 16328
rect 144012 16318 144040 75140
rect 144000 16312 144052 16318
rect 144000 16254 144052 16260
rect 144104 7954 144132 75140
rect 144196 33862 144224 75140
rect 144184 33856 144236 33862
rect 144184 33798 144236 33804
rect 144288 16250 144316 75140
rect 144380 26042 144408 75140
rect 144368 26036 144420 26042
rect 144368 25978 144420 25984
rect 144276 16244 144328 16250
rect 144276 16186 144328 16192
rect 144472 10606 144500 75140
rect 144564 71913 144592 75140
rect 144656 72049 144684 75140
rect 144748 72185 144776 75140
rect 144734 72176 144790 72185
rect 144734 72111 144790 72120
rect 144642 72040 144698 72049
rect 144642 71975 144698 71984
rect 144840 71913 144868 75140
rect 144550 71904 144606 71913
rect 144550 71839 144606 71848
rect 144826 71904 144882 71913
rect 144826 71839 144882 71848
rect 144932 30258 144960 75140
rect 145024 33794 145052 75140
rect 145116 74254 145144 75140
rect 145104 74248 145156 74254
rect 145104 74190 145156 74196
rect 145104 73024 145156 73030
rect 145104 72966 145156 72972
rect 145116 72078 145144 72966
rect 145104 72072 145156 72078
rect 145104 72014 145156 72020
rect 145012 33788 145064 33794
rect 145012 33730 145064 33736
rect 144920 30252 144972 30258
rect 144920 30194 144972 30200
rect 145208 30190 145236 75140
rect 145300 35154 145328 75140
rect 145288 35148 145340 35154
rect 145288 35090 145340 35096
rect 145196 30184 145248 30190
rect 145196 30126 145248 30132
rect 144460 10600 144512 10606
rect 144460 10542 144512 10548
rect 145392 9518 145420 75140
rect 145484 72282 145512 75140
rect 145472 72276 145524 72282
rect 145472 72218 145524 72224
rect 145576 35902 145604 75140
rect 145564 35896 145616 35902
rect 145564 35838 145616 35844
rect 145380 9512 145432 9518
rect 145380 9454 145432 9460
rect 145668 9450 145696 75140
rect 145656 9444 145708 9450
rect 145656 9386 145708 9392
rect 145760 9382 145788 75140
rect 145852 71806 145880 75140
rect 145840 71800 145892 71806
rect 145840 71742 145892 71748
rect 145944 10538 145972 75140
rect 146036 72185 146064 75140
rect 146022 72176 146078 72185
rect 146022 72111 146078 72120
rect 146024 72072 146076 72078
rect 146024 72014 146076 72020
rect 146036 27402 146064 72014
rect 146128 71913 146156 75140
rect 146220 72049 146248 75140
rect 146206 72040 146262 72049
rect 146206 71975 146262 71984
rect 146114 71904 146170 71913
rect 146114 71839 146170 71848
rect 146024 27396 146076 27402
rect 146024 27338 146076 27344
rect 145932 10532 145984 10538
rect 145932 10474 145984 10480
rect 146312 10470 146340 75140
rect 146404 35766 146432 75140
rect 146496 74594 146524 75140
rect 146484 74588 146536 74594
rect 146484 74530 146536 74536
rect 146392 35760 146444 35766
rect 146392 35702 146444 35708
rect 146588 12034 146616 75140
rect 146680 35698 146708 75140
rect 146772 74186 146800 75140
rect 146760 74180 146812 74186
rect 146760 74122 146812 74128
rect 146760 72752 146812 72758
rect 146760 72694 146812 72700
rect 146772 71874 146800 72694
rect 146760 71868 146812 71874
rect 146760 71810 146812 71816
rect 146668 35692 146720 35698
rect 146668 35634 146720 35640
rect 146864 13326 146892 75140
rect 146956 35630 146984 75140
rect 146944 35624 146996 35630
rect 146944 35566 146996 35572
rect 147048 17610 147076 75140
rect 147036 17604 147088 17610
rect 147036 17546 147088 17552
rect 146852 13320 146904 13326
rect 146852 13262 146904 13268
rect 147140 13258 147168 75140
rect 147232 20330 147260 75140
rect 147324 71913 147352 75140
rect 147416 72049 147444 75140
rect 147508 72185 147536 75140
rect 147494 72176 147550 72185
rect 147494 72111 147550 72120
rect 147402 72040 147458 72049
rect 147402 71975 147458 71984
rect 147600 71913 147628 75140
rect 147310 71904 147366 71913
rect 147310 71839 147366 71848
rect 147586 71904 147642 71913
rect 147586 71839 147642 71848
rect 147312 71800 147364 71806
rect 147312 71742 147364 71748
rect 147324 35834 147352 71742
rect 147312 35828 147364 35834
rect 147312 35770 147364 35776
rect 147220 20324 147272 20330
rect 147220 20266 147272 20272
rect 147128 13252 147180 13258
rect 147128 13194 147180 13200
rect 146576 12028 146628 12034
rect 146576 11970 146628 11976
rect 146300 10464 146352 10470
rect 146300 10406 146352 10412
rect 145748 9376 145800 9382
rect 145748 9318 145800 9324
rect 144092 7948 144144 7954
rect 144092 7890 144144 7896
rect 147692 7886 147720 75140
rect 147784 35562 147812 75140
rect 147876 74662 147904 75140
rect 147864 74656 147916 74662
rect 147864 74598 147916 74604
rect 147864 73228 147916 73234
rect 147864 73170 147916 73176
rect 147876 72962 147904 73170
rect 147864 72956 147916 72962
rect 147864 72898 147916 72904
rect 147772 35556 147824 35562
rect 147772 35498 147824 35504
rect 147968 9314 147996 75140
rect 148060 22030 148088 75140
rect 148048 22024 148100 22030
rect 148048 21966 148100 21972
rect 147956 9308 148008 9314
rect 147956 9250 148008 9256
rect 148152 9246 148180 75140
rect 148244 11966 148272 75140
rect 148336 27062 148364 75140
rect 148324 27056 148376 27062
rect 148324 26998 148376 27004
rect 148232 11960 148284 11966
rect 148232 11902 148284 11908
rect 148428 11898 148456 75140
rect 148520 16182 148548 75140
rect 148612 35494 148640 75140
rect 148704 72729 148732 75140
rect 148690 72720 148746 72729
rect 148690 72655 148746 72664
rect 148796 72457 148824 75140
rect 148888 72593 148916 75140
rect 148980 72865 149008 75140
rect 148966 72856 149022 72865
rect 148966 72791 149022 72800
rect 148874 72584 148930 72593
rect 148874 72519 148930 72528
rect 148782 72448 148838 72457
rect 148782 72383 148838 72392
rect 148600 35488 148652 35494
rect 148600 35430 148652 35436
rect 148508 16176 148560 16182
rect 148508 16118 148560 16124
rect 149072 16114 149100 75140
rect 149164 72010 149192 75140
rect 149152 72004 149204 72010
rect 149152 71946 149204 71952
rect 149060 16108 149112 16114
rect 149060 16050 149112 16056
rect 148416 11892 148468 11898
rect 148416 11834 148468 11840
rect 149256 11830 149284 75140
rect 149348 25974 149376 75140
rect 149440 35358 149468 75140
rect 149428 35352 149480 35358
rect 149428 35294 149480 35300
rect 149336 25968 149388 25974
rect 149336 25910 149388 25916
rect 149532 18970 149560 75140
rect 149520 18964 149572 18970
rect 149520 18906 149572 18912
rect 149624 14686 149652 75140
rect 149716 71942 149744 75140
rect 149704 71936 149756 71942
rect 149704 71878 149756 71884
rect 149612 14680 149664 14686
rect 149612 14622 149664 14628
rect 149808 13190 149836 75140
rect 149796 13184 149848 13190
rect 149796 13126 149848 13132
rect 149244 11824 149296 11830
rect 149244 11766 149296 11772
rect 148140 9240 148192 9246
rect 148140 9182 148192 9188
rect 147680 7880 147732 7886
rect 147680 7822 147732 7828
rect 143816 6656 143868 6662
rect 143816 6598 143868 6604
rect 142436 5432 142488 5438
rect 142436 5374 142488 5380
rect 140042 3496 140098 3505
rect 140042 3431 140098 3440
rect 140056 480 140084 3431
rect 141240 2984 141292 2990
rect 141240 2926 141292 2932
rect 141252 480 141280 2926
rect 142448 480 142476 5374
rect 144736 5364 144788 5370
rect 144736 5306 144788 5312
rect 143540 4140 143592 4146
rect 143540 4082 143592 4088
rect 143552 480 143580 4082
rect 144748 480 144776 5306
rect 149900 5166 149928 75140
rect 149992 72729 150020 75140
rect 149978 72720 150034 72729
rect 149978 72655 150034 72664
rect 150084 72593 150112 75140
rect 150176 73001 150204 75140
rect 150162 72992 150218 73001
rect 150268 72962 150296 75140
rect 150162 72927 150218 72936
rect 150256 72956 150308 72962
rect 150256 72898 150308 72904
rect 150360 72865 150388 75140
rect 150346 72856 150402 72865
rect 150346 72791 150402 72800
rect 150070 72584 150126 72593
rect 149980 72548 150032 72554
rect 150070 72519 150126 72528
rect 149980 72490 150032 72496
rect 149992 70394 150020 72490
rect 150164 72208 150216 72214
rect 150164 72150 150216 72156
rect 149992 70366 150112 70394
rect 148324 5160 148376 5166
rect 148324 5102 148376 5108
rect 149888 5160 149940 5166
rect 149888 5102 149940 5108
rect 146944 4072 146996 4078
rect 146944 4014 146996 4020
rect 145932 4004 145984 4010
rect 145932 3946 145984 3952
rect 145944 480 145972 3946
rect 146956 3398 146984 4014
rect 147128 3596 147180 3602
rect 147128 3538 147180 3544
rect 146944 3392 146996 3398
rect 146944 3334 146996 3340
rect 147140 480 147168 3538
rect 148336 480 148364 5102
rect 149520 5092 149572 5098
rect 149520 5034 149572 5040
rect 149532 480 149560 5034
rect 150084 3330 150112 70366
rect 150176 28082 150204 72150
rect 150452 28422 150480 75140
rect 150440 28416 150492 28422
rect 150440 28358 150492 28364
rect 150164 28076 150216 28082
rect 150164 28018 150216 28024
rect 150544 25906 150572 75140
rect 150636 74118 150664 75140
rect 150624 74112 150676 74118
rect 150624 74054 150676 74060
rect 150624 72888 150676 72894
rect 150624 72830 150676 72836
rect 150636 28694 150664 72830
rect 150728 30122 150756 75140
rect 150820 72350 150848 75140
rect 150808 72344 150860 72350
rect 150808 72286 150860 72292
rect 150716 30116 150768 30122
rect 150716 30058 150768 30064
rect 150624 28688 150676 28694
rect 150624 28630 150676 28636
rect 150532 25900 150584 25906
rect 150532 25842 150584 25848
rect 150912 18902 150940 75140
rect 150900 18896 150952 18902
rect 150900 18838 150952 18844
rect 151004 13122 151032 75140
rect 150992 13116 151044 13122
rect 150992 13058 151044 13064
rect 151096 6594 151124 75140
rect 151188 18834 151216 75140
rect 151280 72622 151308 75140
rect 151268 72616 151320 72622
rect 151268 72558 151320 72564
rect 151372 72078 151400 75140
rect 151360 72072 151412 72078
rect 151360 72014 151412 72020
rect 151176 18828 151228 18834
rect 151176 18770 151228 18776
rect 151464 14618 151492 75140
rect 151556 72729 151584 75140
rect 151542 72720 151598 72729
rect 151542 72655 151598 72664
rect 151648 72457 151676 75140
rect 151740 72865 151768 75140
rect 151832 73030 151860 75140
rect 151820 73024 151872 73030
rect 151820 72966 151872 72972
rect 151726 72856 151782 72865
rect 151726 72791 151782 72800
rect 151820 72820 151872 72826
rect 151820 72762 151872 72768
rect 151634 72448 151690 72457
rect 151634 72383 151690 72392
rect 151832 72282 151860 72762
rect 151924 72758 151952 75140
rect 152016 74633 152044 75140
rect 152002 74624 152058 74633
rect 152002 74559 152058 74568
rect 152004 73024 152056 73030
rect 152004 72966 152056 72972
rect 151912 72752 151964 72758
rect 151912 72694 151964 72700
rect 152016 72554 152044 72966
rect 152004 72548 152056 72554
rect 152004 72490 152056 72496
rect 151820 72276 151872 72282
rect 151820 72218 151872 72224
rect 151636 71868 151688 71874
rect 151636 71810 151688 71816
rect 151648 64874 151676 71810
rect 151556 64846 151676 64874
rect 151556 28898 151584 64846
rect 151544 28892 151596 28898
rect 151544 28834 151596 28840
rect 151452 14612 151504 14618
rect 151452 14554 151504 14560
rect 152108 9178 152136 75140
rect 152200 72214 152228 75140
rect 152188 72208 152240 72214
rect 152188 72150 152240 72156
rect 152292 20194 152320 75140
rect 152280 20188 152332 20194
rect 152280 20130 152332 20136
rect 152096 9172 152148 9178
rect 152096 9114 152148 9120
rect 151084 6588 151136 6594
rect 151084 6530 151136 6536
rect 152384 6526 152412 75140
rect 152476 36650 152504 75140
rect 152464 36644 152516 36650
rect 152464 36586 152516 36592
rect 152568 20126 152596 75140
rect 152556 20120 152608 20126
rect 152556 20062 152608 20068
rect 152660 10402 152688 75140
rect 152752 73030 152780 75140
rect 152740 73024 152792 73030
rect 152740 72966 152792 72972
rect 152844 72457 152872 75140
rect 152936 72865 152964 75140
rect 152922 72856 152978 72865
rect 152922 72791 152978 72800
rect 153028 72729 153056 75140
rect 153014 72720 153070 72729
rect 152924 72684 152976 72690
rect 153014 72655 153070 72664
rect 152924 72626 152976 72632
rect 152936 72570 152964 72626
rect 153120 72593 153148 75140
rect 153106 72584 153162 72593
rect 152936 72542 153056 72570
rect 152830 72448 152886 72457
rect 153028 72434 153056 72542
rect 153106 72519 153162 72528
rect 152830 72383 152886 72392
rect 152924 72412 152976 72418
rect 153028 72406 153148 72434
rect 152924 72354 152976 72360
rect 152832 72344 152884 72350
rect 152832 72286 152884 72292
rect 152844 28354 152872 72286
rect 152936 28558 152964 72354
rect 153016 72276 153068 72282
rect 153016 72218 153068 72224
rect 152924 28552 152976 28558
rect 152924 28494 152976 28500
rect 153028 28490 153056 72218
rect 153120 40730 153148 72406
rect 153108 40724 153160 40730
rect 153108 40666 153160 40672
rect 153016 28484 153068 28490
rect 153016 28426 153068 28432
rect 152832 28348 152884 28354
rect 152832 28290 152884 28296
rect 153212 24682 153240 75140
rect 153304 71874 153332 75140
rect 153396 74050 153424 75140
rect 153384 74044 153436 74050
rect 153384 73986 153436 73992
rect 153384 73228 153436 73234
rect 153384 73170 153436 73176
rect 153396 72962 153424 73170
rect 153384 72956 153436 72962
rect 153384 72898 153436 72904
rect 153292 71868 153344 71874
rect 153292 71810 153344 71816
rect 153200 24676 153252 24682
rect 153200 24618 153252 24624
rect 152648 10396 152700 10402
rect 152648 10338 152700 10344
rect 153488 9110 153516 75140
rect 153476 9104 153528 9110
rect 153476 9046 153528 9052
rect 153580 9042 153608 75140
rect 153672 20058 153700 75140
rect 153764 25838 153792 75140
rect 153856 72214 153884 75140
rect 153844 72208 153896 72214
rect 153844 72150 153896 72156
rect 153752 25832 153804 25838
rect 153752 25774 153804 25780
rect 153660 20052 153712 20058
rect 153660 19994 153712 20000
rect 153948 16046 153976 75140
rect 153936 16040 153988 16046
rect 153936 15982 153988 15988
rect 153568 9036 153620 9042
rect 153568 8978 153620 8984
rect 154040 7818 154068 75140
rect 154132 72865 154160 75140
rect 154118 72856 154174 72865
rect 154118 72791 154174 72800
rect 154224 72729 154252 75140
rect 154316 73001 154344 75140
rect 154302 72992 154358 73001
rect 154302 72927 154358 72936
rect 154408 72826 154436 75140
rect 154396 72820 154448 72826
rect 154396 72762 154448 72768
rect 154210 72720 154266 72729
rect 154210 72655 154266 72664
rect 154120 72616 154172 72622
rect 154500 72593 154528 75140
rect 154120 72558 154172 72564
rect 154486 72584 154542 72593
rect 154132 64874 154160 72558
rect 154486 72519 154542 72528
rect 154304 72140 154356 72146
rect 154304 72082 154356 72088
rect 154132 64846 154252 64874
rect 154224 30054 154252 64846
rect 154316 30326 154344 72082
rect 154396 72004 154448 72010
rect 154396 71946 154448 71952
rect 154408 64874 154436 71946
rect 154408 64846 154528 64874
rect 154500 35426 154528 64846
rect 154488 35420 154540 35426
rect 154488 35362 154540 35368
rect 154304 30320 154356 30326
rect 154304 30262 154356 30268
rect 154212 30048 154264 30054
rect 154212 29990 154264 29996
rect 154592 26994 154620 75140
rect 154580 26988 154632 26994
rect 154580 26930 154632 26936
rect 154684 14550 154712 75140
rect 154776 74526 154804 75140
rect 154764 74520 154816 74526
rect 154764 74462 154816 74468
rect 154764 72888 154816 72894
rect 154764 72830 154816 72836
rect 154776 68882 154804 72830
rect 154764 68876 154816 68882
rect 154764 68818 154816 68824
rect 154868 17542 154896 75140
rect 154960 72282 154988 75140
rect 154948 72276 155000 72282
rect 154948 72218 155000 72224
rect 155052 21894 155080 75140
rect 155144 29918 155172 75140
rect 155132 29912 155184 29918
rect 155132 29854 155184 29860
rect 155040 21888 155092 21894
rect 155040 21830 155092 21836
rect 155236 21826 155264 75140
rect 155224 21820 155276 21826
rect 155224 21762 155276 21768
rect 154856 17536 154908 17542
rect 154856 17478 154908 17484
rect 155328 17474 155356 75140
rect 155316 17468 155368 17474
rect 155316 17410 155368 17416
rect 155420 17406 155448 75140
rect 155512 73710 155540 75140
rect 155500 73704 155552 73710
rect 155500 73646 155552 73652
rect 155500 72752 155552 72758
rect 155500 72694 155552 72700
rect 155512 36718 155540 72694
rect 155500 36712 155552 36718
rect 155500 36654 155552 36660
rect 155408 17400 155460 17406
rect 155408 17342 155460 17348
rect 155604 17338 155632 75140
rect 155696 72457 155724 75140
rect 155788 72865 155816 75140
rect 155774 72856 155830 72865
rect 155774 72791 155830 72800
rect 155880 72729 155908 75140
rect 155866 72720 155922 72729
rect 155866 72655 155922 72664
rect 155682 72448 155738 72457
rect 155682 72383 155738 72392
rect 155972 29782 156000 75140
rect 156064 72418 156092 75140
rect 156156 74934 156184 75140
rect 156144 74928 156196 74934
rect 156144 74870 156196 74876
rect 156144 74792 156196 74798
rect 156144 74734 156196 74740
rect 156156 73166 156184 74734
rect 156144 73160 156196 73166
rect 156144 73102 156196 73108
rect 156052 72412 156104 72418
rect 156052 72354 156104 72360
rect 155960 29776 156012 29782
rect 155960 29718 156012 29724
rect 156248 29714 156276 75140
rect 156236 29708 156288 29714
rect 156236 29650 156288 29656
rect 156340 21758 156368 75140
rect 156328 21752 156380 21758
rect 156328 21694 156380 21700
rect 156432 21690 156460 75140
rect 156420 21684 156472 21690
rect 156420 21626 156472 21632
rect 155592 17332 155644 17338
rect 155592 17274 155644 17280
rect 154672 14544 154724 14550
rect 154672 14486 154724 14492
rect 156524 10334 156552 75140
rect 156616 72894 156644 75140
rect 156604 72888 156656 72894
rect 156604 72830 156656 72836
rect 156604 72548 156656 72554
rect 156604 72490 156656 72496
rect 156616 69698 156644 72490
rect 156604 69692 156656 69698
rect 156604 69634 156656 69640
rect 156708 18766 156736 75140
rect 156800 29646 156828 75140
rect 156892 72729 156920 75140
rect 156984 72865 157012 75140
rect 156970 72856 157026 72865
rect 156970 72791 157026 72800
rect 156878 72720 156934 72729
rect 156878 72655 156934 72664
rect 157076 72593 157104 75140
rect 157062 72584 157118 72593
rect 157062 72519 157118 72528
rect 157062 72448 157118 72457
rect 157062 72383 157118 72392
rect 156880 71936 156932 71942
rect 156880 71878 156932 71884
rect 156788 29640 156840 29646
rect 156788 29582 156840 29588
rect 156892 21962 156920 71878
rect 156972 69692 157024 69698
rect 156972 69634 157024 69640
rect 156984 29986 157012 69634
rect 156972 29980 157024 29986
rect 156972 29922 157024 29928
rect 157076 29850 157104 72383
rect 157168 72185 157196 75140
rect 157260 72729 157288 75140
rect 157246 72720 157302 72729
rect 157246 72655 157302 72664
rect 157154 72176 157210 72185
rect 157154 72111 157210 72120
rect 157064 29844 157116 29850
rect 157064 29786 157116 29792
rect 157352 23458 157380 75140
rect 157444 72826 157472 75140
rect 157536 74798 157564 75140
rect 157524 74792 157576 74798
rect 157524 74734 157576 74740
rect 157524 74656 157576 74662
rect 157522 74624 157524 74633
rect 157576 74624 157578 74633
rect 157522 74559 157578 74568
rect 157432 72820 157484 72826
rect 157432 72762 157484 72768
rect 157628 31754 157656 75140
rect 157616 31748 157668 31754
rect 157616 31690 157668 31696
rect 157340 23452 157392 23458
rect 157340 23394 157392 23400
rect 156880 21956 156932 21962
rect 156880 21898 156932 21904
rect 156696 18760 156748 18766
rect 156696 18702 156748 18708
rect 157720 12306 157748 75140
rect 157812 74594 157840 75140
rect 157800 74588 157852 74594
rect 157800 74530 157852 74536
rect 157798 72176 157854 72185
rect 157798 72111 157854 72120
rect 157812 36582 157840 72111
rect 157800 36576 157852 36582
rect 157800 36518 157852 36524
rect 157904 14482 157932 75140
rect 157996 26926 158024 75140
rect 157984 26920 158036 26926
rect 157984 26862 158036 26868
rect 158088 19990 158116 75140
rect 158180 31686 158208 75140
rect 158272 72758 158300 75140
rect 158260 72752 158312 72758
rect 158364 72729 158392 75140
rect 158260 72694 158312 72700
rect 158350 72720 158406 72729
rect 158350 72655 158406 72664
rect 158456 72593 158484 75140
rect 158442 72584 158498 72593
rect 158442 72519 158498 72528
rect 158548 72457 158576 75140
rect 158640 72865 158668 75140
rect 158626 72856 158682 72865
rect 158626 72791 158682 72800
rect 158628 72752 158680 72758
rect 158628 72694 158680 72700
rect 158640 72622 158668 72694
rect 158628 72616 158680 72622
rect 158628 72558 158680 72564
rect 158534 72448 158590 72457
rect 158534 72383 158590 72392
rect 158444 72072 158496 72078
rect 158444 72014 158496 72020
rect 158352 68876 158404 68882
rect 158352 68818 158404 68824
rect 158364 35290 158392 68818
rect 158352 35284 158404 35290
rect 158352 35226 158404 35232
rect 158456 35222 158484 72014
rect 158444 35216 158496 35222
rect 158444 35158 158496 35164
rect 158168 31680 158220 31686
rect 158168 31622 158220 31628
rect 158732 31618 158760 75140
rect 158824 71913 158852 75140
rect 158916 72049 158944 75140
rect 158902 72040 158958 72049
rect 158902 71975 158958 71984
rect 158810 71904 158866 71913
rect 158810 71839 158866 71848
rect 158720 31612 158772 31618
rect 158720 31554 158772 31560
rect 159008 21622 159036 75140
rect 159100 31550 159128 75140
rect 159088 31544 159140 31550
rect 159088 31486 159140 31492
rect 158996 21616 159048 21622
rect 158996 21558 159048 21564
rect 158076 19984 158128 19990
rect 158076 19926 158128 19932
rect 157892 14476 157944 14482
rect 157892 14418 157944 14424
rect 157708 12300 157760 12306
rect 157708 12242 157760 12248
rect 156512 10328 156564 10334
rect 156512 10270 156564 10276
rect 154028 7812 154080 7818
rect 154028 7754 154080 7760
rect 152372 6520 152424 6526
rect 152372 6462 152424 6468
rect 153016 5024 153068 5030
rect 153016 4966 153068 4972
rect 155406 4992 155462 5001
rect 151820 4956 151872 4962
rect 151820 4898 151872 4904
rect 150624 3528 150676 3534
rect 150624 3470 150676 3476
rect 150072 3324 150124 3330
rect 150072 3266 150124 3272
rect 150636 480 150664 3470
rect 151832 480 151860 4898
rect 153028 480 153056 4966
rect 155406 4927 155462 4936
rect 154212 3460 154264 3466
rect 154212 3402 154264 3408
rect 154224 480 154252 3402
rect 155420 480 155448 4927
rect 158904 4888 158956 4894
rect 156602 4856 156658 4865
rect 158904 4830 158956 4836
rect 156602 4791 156658 4800
rect 156616 480 156644 4791
rect 157798 3360 157854 3369
rect 157798 3295 157854 3304
rect 157812 480 157840 3295
rect 158916 480 158944 4830
rect 159192 3602 159220 75140
rect 159284 21554 159312 75140
rect 159272 21548 159324 21554
rect 159272 21490 159324 21496
rect 159376 11762 159404 75140
rect 159364 11756 159416 11762
rect 159364 11698 159416 11704
rect 159180 3596 159232 3602
rect 159180 3538 159232 3544
rect 159468 3534 159496 75140
rect 159560 21486 159588 75140
rect 159652 72321 159680 75140
rect 159638 72312 159694 72321
rect 159638 72247 159694 72256
rect 159548 21480 159600 21486
rect 159548 21422 159600 21428
rect 159456 3528 159508 3534
rect 159456 3470 159508 3476
rect 159744 3466 159772 75140
rect 159836 21418 159864 75140
rect 159928 72865 159956 75140
rect 159914 72856 159970 72865
rect 159914 72791 159970 72800
rect 160020 72729 160048 75140
rect 160006 72720 160062 72729
rect 160006 72655 160062 72664
rect 160112 23390 160140 75140
rect 160204 31414 160232 75140
rect 160296 72185 160324 75140
rect 160282 72176 160338 72185
rect 160282 72111 160338 72120
rect 160192 31408 160244 31414
rect 160192 31350 160244 31356
rect 160100 23384 160152 23390
rect 160100 23326 160152 23332
rect 160388 23322 160416 75140
rect 160376 23316 160428 23322
rect 160376 23258 160428 23264
rect 159824 21412 159876 21418
rect 159824 21354 159876 21360
rect 160480 5098 160508 75140
rect 160468 5092 160520 5098
rect 160468 5034 160520 5040
rect 160572 5030 160600 75140
rect 160664 23254 160692 75140
rect 160756 31346 160784 75140
rect 160744 31340 160796 31346
rect 160744 31282 160796 31288
rect 160652 23248 160704 23254
rect 160652 23190 160704 23196
rect 160560 5024 160612 5030
rect 160560 4966 160612 4972
rect 160100 4072 160152 4078
rect 160100 4014 160152 4020
rect 159732 3460 159784 3466
rect 159732 3402 159784 3408
rect 160112 480 160140 4014
rect 160848 3913 160876 75140
rect 160940 23186 160968 75140
rect 161032 72729 161060 75140
rect 161018 72720 161074 72729
rect 161018 72655 161074 72664
rect 161124 72457 161152 75140
rect 161216 72865 161244 75140
rect 161308 73137 161336 75140
rect 161294 73128 161350 73137
rect 161294 73063 161350 73072
rect 161202 72856 161258 72865
rect 161202 72791 161258 72800
rect 161400 72593 161428 75140
rect 161386 72584 161442 72593
rect 161386 72519 161442 72528
rect 161110 72448 161166 72457
rect 161110 72383 161166 72392
rect 161018 72312 161074 72321
rect 161018 72247 161074 72256
rect 161032 31482 161060 72247
rect 161020 31476 161072 31482
rect 161020 31418 161072 31424
rect 160928 23180 160980 23186
rect 160928 23122 160980 23128
rect 161492 23118 161520 75140
rect 161480 23112 161532 23118
rect 161480 23054 161532 23060
rect 161584 6322 161612 75140
rect 161676 74361 161704 75140
rect 161662 74352 161718 74361
rect 161662 74287 161718 74296
rect 161664 73908 161716 73914
rect 161664 73850 161716 73856
rect 161676 73574 161704 73850
rect 161664 73568 161716 73574
rect 161664 73510 161716 73516
rect 161768 23050 161796 75140
rect 161860 31210 161888 75140
rect 161848 31204 161900 31210
rect 161848 31146 161900 31152
rect 161756 23044 161808 23050
rect 161756 22986 161808 22992
rect 161572 6316 161624 6322
rect 161572 6258 161624 6264
rect 161952 4962 161980 75140
rect 162044 22982 162072 75140
rect 162136 31074 162164 75140
rect 162124 31068 162176 31074
rect 162124 31010 162176 31016
rect 162032 22976 162084 22982
rect 162032 22918 162084 22924
rect 161940 4956 161992 4962
rect 161940 4898 161992 4904
rect 162228 4894 162256 75140
rect 162320 22914 162348 75140
rect 162412 74905 162440 75140
rect 162398 74896 162454 74905
rect 162398 74831 162454 74840
rect 162398 74352 162454 74361
rect 162398 74287 162454 74296
rect 162412 73273 162440 74287
rect 162398 73264 162454 73273
rect 162398 73199 162454 73208
rect 162398 73128 162454 73137
rect 162398 73063 162454 73072
rect 162412 64874 162440 73063
rect 162504 72729 162532 75140
rect 162596 73001 162624 75140
rect 162582 72992 162638 73001
rect 162582 72927 162638 72936
rect 162490 72720 162546 72729
rect 162490 72655 162546 72664
rect 162688 72593 162716 75140
rect 162780 72865 162808 75140
rect 162766 72856 162822 72865
rect 162766 72791 162822 72800
rect 162674 72584 162730 72593
rect 162674 72519 162730 72528
rect 162766 72448 162822 72457
rect 162766 72383 162822 72392
rect 162780 72078 162808 72383
rect 162768 72072 162820 72078
rect 162768 72014 162820 72020
rect 162412 64846 162624 64874
rect 162596 31278 162624 64846
rect 162584 31272 162636 31278
rect 162584 31214 162636 31220
rect 162872 24614 162900 75140
rect 162860 24608 162912 24614
rect 162860 24550 162912 24556
rect 162308 22908 162360 22914
rect 162308 22850 162360 22856
rect 162964 15910 162992 75140
rect 163056 73137 163084 75140
rect 163042 73128 163098 73137
rect 163042 73063 163098 73072
rect 163148 24546 163176 75140
rect 163136 24540 163188 24546
rect 163136 24482 163188 24488
rect 163240 18698 163268 75140
rect 163332 73001 163360 75140
rect 163318 72992 163374 73001
rect 163318 72927 163374 72936
rect 163424 24478 163452 75140
rect 163516 58682 163544 75140
rect 163504 58676 163556 58682
rect 163504 58618 163556 58624
rect 163412 24472 163464 24478
rect 163412 24414 163464 24420
rect 163228 18692 163280 18698
rect 163228 18634 163280 18640
rect 162952 15904 163004 15910
rect 162952 15846 163004 15852
rect 163608 6254 163636 75140
rect 163700 24410 163728 75140
rect 163688 24404 163740 24410
rect 163688 24346 163740 24352
rect 163792 19038 163820 75140
rect 163780 19032 163832 19038
rect 163780 18974 163832 18980
rect 163596 6248 163648 6254
rect 163596 6190 163648 6196
rect 163884 6186 163912 75140
rect 163976 72729 164004 75140
rect 164068 72865 164096 75140
rect 164054 72856 164110 72865
rect 164054 72791 164110 72800
rect 163962 72720 164018 72729
rect 163962 72655 164018 72664
rect 164160 72457 164188 75140
rect 164146 72448 164202 72457
rect 164146 72383 164202 72392
rect 164252 24342 164280 75140
rect 164344 32502 164372 75140
rect 164436 73846 164464 75140
rect 164424 73840 164476 73846
rect 164424 73782 164476 73788
rect 164332 32496 164384 32502
rect 164332 32438 164384 32444
rect 164240 24336 164292 24342
rect 164240 24278 164292 24284
rect 164528 24274 164556 75140
rect 164516 24268 164568 24274
rect 164516 24210 164568 24216
rect 164620 18630 164648 75140
rect 164608 18624 164660 18630
rect 164608 18566 164660 18572
rect 164712 7750 164740 75140
rect 164804 25770 164832 75140
rect 164792 25764 164844 25770
rect 164792 25706 164844 25712
rect 164896 17270 164924 75140
rect 164884 17264 164936 17270
rect 164884 17206 164936 17212
rect 164700 7744 164752 7750
rect 164700 7686 164752 7692
rect 164988 7682 165016 75140
rect 165080 71874 165108 75140
rect 165068 71868 165120 71874
rect 165068 71810 165120 71816
rect 165172 22846 165200 75140
rect 165264 72729 165292 75140
rect 165250 72720 165306 72729
rect 165250 72655 165306 72664
rect 165252 72480 165304 72486
rect 165356 72457 165384 75140
rect 165448 72593 165476 75140
rect 165540 72865 165568 75140
rect 165526 72856 165582 72865
rect 165526 72791 165582 72800
rect 165434 72584 165490 72593
rect 165434 72519 165490 72528
rect 165252 72422 165304 72428
rect 165342 72448 165398 72457
rect 165160 22840 165212 22846
rect 165160 22782 165212 22788
rect 164976 7676 165028 7682
rect 164976 7618 165028 7624
rect 163872 6180 163924 6186
rect 163872 6122 163924 6128
rect 162216 4888 162268 4894
rect 162216 4830 162268 4836
rect 163688 4820 163740 4826
rect 163688 4762 163740 4768
rect 161296 3936 161348 3942
rect 160834 3904 160890 3913
rect 161296 3878 161348 3884
rect 160834 3839 160890 3848
rect 161308 480 161336 3878
rect 162492 3868 162544 3874
rect 162492 3810 162544 3816
rect 162504 480 162532 3810
rect 163700 480 163728 4762
rect 164884 3800 164936 3806
rect 164884 3742 164936 3748
rect 164896 480 164924 3742
rect 165264 3262 165292 72422
rect 165342 72383 165398 72392
rect 165632 25634 165660 75140
rect 165620 25628 165672 25634
rect 165620 25570 165672 25576
rect 165724 24206 165752 75140
rect 165712 24200 165764 24206
rect 165712 24142 165764 24148
rect 165816 7614 165844 75140
rect 165908 24138 165936 75140
rect 166000 28286 166028 75140
rect 165988 28280 166040 28286
rect 165988 28222 166040 28228
rect 165896 24132 165948 24138
rect 165896 24074 165948 24080
rect 166092 8974 166120 75140
rect 166184 25566 166212 75140
rect 166276 32434 166304 75140
rect 166368 72593 166396 75140
rect 166460 72729 166488 75140
rect 166446 72720 166502 72729
rect 166446 72655 166502 72664
rect 166354 72584 166410 72593
rect 166354 72519 166410 72528
rect 166552 72457 166580 75140
rect 166644 72758 166672 75140
rect 166632 72752 166684 72758
rect 166632 72694 166684 72700
rect 166736 72554 166764 75140
rect 166828 72729 166856 75140
rect 166814 72720 166870 72729
rect 166814 72655 166870 72664
rect 166814 72584 166870 72593
rect 166724 72548 166776 72554
rect 166814 72519 166870 72528
rect 166724 72490 166776 72496
rect 166538 72448 166594 72457
rect 166538 72383 166594 72392
rect 166724 72072 166776 72078
rect 166828 72049 166856 72519
rect 166920 72486 166948 75140
rect 167012 73930 167040 75140
rect 167104 74526 167132 75140
rect 167092 74520 167144 74526
rect 167196 74497 167224 75140
rect 167092 74462 167144 74468
rect 167182 74488 167238 74497
rect 167182 74423 167238 74432
rect 167288 74225 167316 75140
rect 167274 74216 167330 74225
rect 167274 74151 167330 74160
rect 167012 73902 167316 73930
rect 167184 73500 167236 73506
rect 167184 73442 167236 73448
rect 166908 72480 166960 72486
rect 166908 72422 166960 72428
rect 166724 72014 166776 72020
rect 166814 72040 166870 72049
rect 166632 71868 166684 71874
rect 166632 71810 166684 71816
rect 166264 32428 166316 32434
rect 166264 32370 166316 32376
rect 166644 25702 166672 71810
rect 166736 31142 166764 72014
rect 166814 71975 166870 71984
rect 166906 31784 166962 31793
rect 166906 31719 166962 31728
rect 166724 31136 166776 31142
rect 166724 31078 166776 31084
rect 166632 25696 166684 25702
rect 166632 25638 166684 25644
rect 166172 25560 166224 25566
rect 166172 25502 166224 25508
rect 166080 8968 166132 8974
rect 166080 8910 166132 8916
rect 165804 7608 165856 7614
rect 165804 7550 165856 7556
rect 166920 4826 166948 31719
rect 167196 6390 167224 73442
rect 167288 72010 167316 73902
rect 167380 73681 167408 75140
rect 167472 74905 167500 75140
rect 167458 74896 167514 74905
rect 167564 74866 167592 75140
rect 167458 74831 167514 74840
rect 167552 74860 167604 74866
rect 167552 74802 167604 74808
rect 167656 74769 167684 75140
rect 167748 74905 167776 75140
rect 167734 74896 167790 74905
rect 167734 74831 167790 74840
rect 167736 74792 167788 74798
rect 167642 74760 167698 74769
rect 167736 74734 167788 74740
rect 167642 74695 167698 74704
rect 167552 74588 167604 74594
rect 167552 74530 167604 74536
rect 167748 74534 167776 74734
rect 167366 73672 167422 73681
rect 167366 73607 167422 73616
rect 167368 72140 167420 72146
rect 167368 72082 167420 72088
rect 167276 72004 167328 72010
rect 167276 71946 167328 71952
rect 167276 69624 167328 69630
rect 167276 69566 167328 69572
rect 167184 6384 167236 6390
rect 167184 6326 167236 6332
rect 167184 5296 167236 5302
rect 167184 5238 167236 5244
rect 166908 4820 166960 4826
rect 166908 4762 166960 4768
rect 166080 3732 166132 3738
rect 166080 3674 166132 3680
rect 165252 3256 165304 3262
rect 165252 3198 165304 3204
rect 166092 480 166120 3674
rect 167196 480 167224 5238
rect 167288 3874 167316 69566
rect 167380 4010 167408 72082
rect 167564 69698 167592 74530
rect 167656 74506 167776 74534
rect 167656 72944 167684 74506
rect 167840 73098 167868 75140
rect 167932 73166 167960 75140
rect 167920 73160 167972 73166
rect 168024 73137 168052 75140
rect 168116 74633 168144 75140
rect 168102 74624 168158 74633
rect 168208 74594 168236 75140
rect 168102 74559 168158 74568
rect 168196 74588 168248 74594
rect 168196 74530 168248 74536
rect 168194 74488 168250 74497
rect 168194 74423 168250 74432
rect 168208 73817 168236 74423
rect 168300 73914 168328 75140
rect 168392 73982 168420 75140
rect 168380 73976 168432 73982
rect 168380 73918 168432 73924
rect 168288 73908 168340 73914
rect 168288 73850 168340 73856
rect 168194 73808 168250 73817
rect 168194 73743 168250 73752
rect 168196 73704 168248 73710
rect 168196 73646 168248 73652
rect 167920 73102 167972 73108
rect 168010 73128 168066 73137
rect 167828 73092 167880 73098
rect 168010 73063 168066 73072
rect 167828 73034 167880 73040
rect 168012 73024 168064 73030
rect 168012 72966 168064 72972
rect 167920 72956 167972 72962
rect 167656 72916 167868 72944
rect 167644 72344 167696 72350
rect 167644 72286 167696 72292
rect 167552 69692 167604 69698
rect 167552 69634 167604 69640
rect 167656 69578 167684 72286
rect 167736 72208 167788 72214
rect 167736 72150 167788 72156
rect 167472 69550 167684 69578
rect 167368 4004 167420 4010
rect 167368 3946 167420 3952
rect 167276 3868 167328 3874
rect 167276 3810 167328 3816
rect 167472 3398 167500 69550
rect 167552 69488 167604 69494
rect 167748 69442 167776 72150
rect 167552 69430 167604 69436
rect 167564 4146 167592 69430
rect 167656 69414 167776 69442
rect 167552 4140 167604 4146
rect 167552 4082 167604 4088
rect 167656 3942 167684 69414
rect 167840 67634 167868 72916
rect 167920 72898 167972 72904
rect 167932 69494 167960 72898
rect 167920 69488 167972 69494
rect 167920 69430 167972 69436
rect 167748 67606 167868 67634
rect 167644 3936 167696 3942
rect 167644 3878 167696 3884
rect 167748 3738 167776 67606
rect 168024 64874 168052 72966
rect 168024 64846 168144 64874
rect 168116 4078 168144 64846
rect 168104 4072 168156 4078
rect 168104 4014 168156 4020
rect 168208 3806 168236 73646
rect 168288 73160 168340 73166
rect 168288 73102 168340 73108
rect 168300 72962 168328 73102
rect 168484 73030 168512 75140
rect 168576 74866 168604 75140
rect 168564 74860 168616 74866
rect 168564 74802 168616 74808
rect 168472 73024 168524 73030
rect 168472 72966 168524 72972
rect 168288 72956 168340 72962
rect 168288 72898 168340 72904
rect 168668 71670 168696 75140
rect 168656 71664 168708 71670
rect 168656 71606 168708 71612
rect 168760 71602 168788 75140
rect 168748 71596 168800 71602
rect 168748 71538 168800 71544
rect 168852 71466 168880 75140
rect 168944 71534 168972 75140
rect 169036 73953 169064 75140
rect 169128 74361 169156 75140
rect 169114 74352 169170 74361
rect 169114 74287 169170 74296
rect 169220 74089 169248 75140
rect 169312 74769 169340 75140
rect 169298 74760 169354 74769
rect 169298 74695 169354 74704
rect 169206 74080 169262 74089
rect 169206 74015 169262 74024
rect 169022 73944 169078 73953
rect 169022 73879 169078 73888
rect 169404 73545 169432 75140
rect 169496 74905 169524 75140
rect 169482 74896 169538 74905
rect 169482 74831 169538 74840
rect 169390 73536 169446 73545
rect 169390 73471 169446 73480
rect 169588 73438 169616 75140
rect 169680 74905 169708 75140
rect 169666 74896 169722 74905
rect 169666 74831 169722 74840
rect 169772 74458 169800 75140
rect 169760 74452 169812 74458
rect 169760 74394 169812 74400
rect 169864 74390 169892 75140
rect 169852 74384 169904 74390
rect 169852 74326 169904 74332
rect 169956 73778 169984 75140
rect 169944 73772 169996 73778
rect 169944 73714 169996 73720
rect 170048 73574 170076 75140
rect 170140 73642 170168 75140
rect 170128 73636 170180 73642
rect 170128 73578 170180 73584
rect 170036 73568 170088 73574
rect 170036 73510 170088 73516
rect 169576 73432 169628 73438
rect 169576 73374 169628 73380
rect 169024 72276 169076 72282
rect 169024 72218 169076 72224
rect 168932 71528 168984 71534
rect 168932 71470 168984 71476
rect 168840 71460 168892 71466
rect 168840 71402 168892 71408
rect 169036 6458 169064 72218
rect 170232 45558 170260 75140
rect 170220 45552 170272 45558
rect 170220 45494 170272 45500
rect 170324 22710 170352 75140
rect 170416 74905 170444 75618
rect 171324 75472 171376 75478
rect 171416 75472 171468 75478
rect 171324 75414 171376 75420
rect 171414 75440 171416 75449
rect 171468 75440 171470 75449
rect 171140 75404 171192 75410
rect 171140 75346 171192 75352
rect 170496 75268 170548 75274
rect 170496 75210 170548 75216
rect 170402 74896 170458 74905
rect 170402 74831 170458 74840
rect 170508 73710 170536 75210
rect 171152 75206 171180 75346
rect 171140 75200 171192 75206
rect 171140 75142 171192 75148
rect 171336 75138 171364 75414
rect 171414 75375 171470 75384
rect 171690 75304 171746 75313
rect 171690 75239 171746 75248
rect 171324 75132 171376 75138
rect 171324 75074 171376 75080
rect 171704 74633 171732 75239
rect 171690 74624 171746 74633
rect 171690 74559 171746 74568
rect 170496 73704 170548 73710
rect 170496 73646 170548 73652
rect 171784 72412 171836 72418
rect 171784 72354 171836 72360
rect 170312 22704 170364 22710
rect 170312 22646 170364 22652
rect 171796 15978 171824 72354
rect 175568 33114 175596 132359
rect 175660 126993 175688 132466
rect 175646 126984 175702 126993
rect 175646 126919 175702 126928
rect 175936 124166 175964 136478
rect 176568 134768 176620 134774
rect 176568 134710 176620 134716
rect 176580 132494 176608 134710
rect 176580 132466 176792 132494
rect 175924 124160 175976 124166
rect 175924 124102 175976 124108
rect 176764 107545 176792 132466
rect 177316 115938 177344 140286
rect 177868 121281 177896 231066
rect 188344 205692 188396 205698
rect 188344 205634 188396 205640
rect 185584 165640 185636 165646
rect 185584 165582 185636 165588
rect 178776 136400 178828 136406
rect 178776 136342 178828 136348
rect 178040 136332 178092 136338
rect 178040 136274 178092 136280
rect 177854 121272 177910 121281
rect 177854 121207 177910 121216
rect 178052 118289 178080 136274
rect 178408 136264 178460 136270
rect 178408 136206 178460 136212
rect 178316 134700 178368 134706
rect 178316 134642 178368 134648
rect 178132 134632 178184 134638
rect 178132 134574 178184 134580
rect 178038 118280 178094 118289
rect 178038 118215 178094 118224
rect 177304 115932 177356 115938
rect 177304 115874 177356 115880
rect 178040 115932 178092 115938
rect 178040 115874 178092 115880
rect 178052 110401 178080 115874
rect 178144 113121 178172 134574
rect 178224 124160 178276 124166
rect 178224 124102 178276 124108
rect 178130 113112 178186 113121
rect 178130 113047 178186 113056
rect 178038 110392 178094 110401
rect 178038 110327 178094 110336
rect 178236 109041 178264 124102
rect 178328 115297 178356 134642
rect 178420 119785 178448 136206
rect 178684 136196 178736 136202
rect 178684 136138 178736 136144
rect 178500 136060 178552 136066
rect 178500 136002 178552 136008
rect 178512 124137 178540 136002
rect 178590 131200 178646 131209
rect 178590 131135 178646 131144
rect 178498 124128 178554 124137
rect 178498 124063 178554 124072
rect 178406 119776 178462 119785
rect 178406 119711 178462 119720
rect 178314 115288 178370 115297
rect 178314 115223 178370 115232
rect 178222 109032 178278 109041
rect 178222 108967 178278 108976
rect 176750 107536 176806 107545
rect 176750 107471 176806 107480
rect 178040 106276 178092 106282
rect 178040 106218 178092 106224
rect 178052 106049 178080 106218
rect 178038 106040 178094 106049
rect 178038 105975 178094 105984
rect 178040 104848 178092 104854
rect 178040 104790 178092 104796
rect 178052 104553 178080 104790
rect 178038 104544 178094 104553
rect 178038 104479 178094 104488
rect 178040 103488 178092 103494
rect 178040 103430 178092 103436
rect 178052 103057 178080 103430
rect 178038 103048 178094 103057
rect 178038 102983 178094 102992
rect 178040 102128 178092 102134
rect 178040 102070 178092 102076
rect 178052 101697 178080 102070
rect 178038 101688 178094 101697
rect 178038 101623 178094 101632
rect 178040 100700 178092 100706
rect 178040 100642 178092 100648
rect 178052 100201 178080 100642
rect 178038 100192 178094 100201
rect 178038 100127 178094 100136
rect 175924 99408 175976 99414
rect 175924 99350 175976 99356
rect 175936 75585 175964 99350
rect 178040 99340 178092 99346
rect 178040 99282 178092 99288
rect 178052 98841 178080 99282
rect 178038 98832 178094 98841
rect 178038 98767 178094 98776
rect 178040 97980 178092 97986
rect 178040 97922 178092 97928
rect 178052 97345 178080 97922
rect 178038 97336 178094 97345
rect 178038 97271 178094 97280
rect 178040 95192 178092 95198
rect 178038 95160 178040 95169
rect 178092 95160 178094 95169
rect 178038 95095 178094 95104
rect 178040 93832 178092 93838
rect 178038 93800 178040 93809
rect 178092 93800 178094 93809
rect 178038 93735 178094 93744
rect 178040 92472 178092 92478
rect 178040 92414 178092 92420
rect 178052 92313 178080 92414
rect 178038 92304 178094 92313
rect 178038 92239 178094 92248
rect 178040 91044 178092 91050
rect 178040 90986 178092 90992
rect 178052 90953 178080 90986
rect 178038 90944 178094 90953
rect 178038 90879 178094 90888
rect 178040 89684 178092 89690
rect 178040 89626 178092 89632
rect 178052 89457 178080 89626
rect 178038 89448 178094 89457
rect 178038 89383 178094 89392
rect 178040 88324 178092 88330
rect 178040 88266 178092 88272
rect 178052 88097 178080 88266
rect 178038 88088 178094 88097
rect 178038 88023 178094 88032
rect 178040 86964 178092 86970
rect 178040 86906 178092 86912
rect 178052 86601 178080 86906
rect 178038 86592 178094 86601
rect 178038 86527 178094 86536
rect 178040 85536 178092 85542
rect 178040 85478 178092 85484
rect 178052 85105 178080 85478
rect 178038 85096 178094 85105
rect 178038 85031 178094 85040
rect 178040 84176 178092 84182
rect 178040 84118 178092 84124
rect 178052 83745 178080 84118
rect 178038 83736 178094 83745
rect 178038 83671 178094 83680
rect 178040 82816 178092 82822
rect 178040 82758 178092 82764
rect 178052 82249 178080 82758
rect 178038 82240 178094 82249
rect 178038 82175 178094 82184
rect 178038 76664 178094 76673
rect 178038 76599 178094 76608
rect 178052 75954 178080 76599
rect 178040 75948 178092 75954
rect 178040 75890 178092 75896
rect 175922 75576 175978 75585
rect 175922 75511 175978 75520
rect 176568 75472 176620 75478
rect 176568 75414 176620 75420
rect 176384 75064 176436 75070
rect 176384 75006 176436 75012
rect 176396 74866 176424 75006
rect 176384 74860 176436 74866
rect 176384 74802 176436 74808
rect 176580 74798 176608 75414
rect 176568 74792 176620 74798
rect 176568 74734 176620 74740
rect 178604 72078 178632 131135
rect 178696 116793 178724 136138
rect 178788 122505 178816 136342
rect 178868 136128 178920 136134
rect 178868 136070 178920 136076
rect 178880 125497 178908 136070
rect 184204 125656 184256 125662
rect 184204 125598 184256 125604
rect 178866 125488 178922 125497
rect 178866 125423 178922 125432
rect 178774 122496 178830 122505
rect 178774 122431 178830 122440
rect 178682 116784 178738 116793
rect 178682 116719 178738 116728
rect 178684 85604 178736 85610
rect 178684 85546 178736 85552
rect 178696 80889 178724 85546
rect 184216 82822 184244 125598
rect 185596 84182 185624 165582
rect 188356 85542 188384 205634
rect 207032 198014 207060 230588
rect 236012 230574 236578 230602
rect 207020 198008 207072 198014
rect 207020 197950 207072 197956
rect 236012 196654 236040 230574
rect 266556 228478 266584 230588
rect 266544 228472 266596 228478
rect 266544 228414 266596 228420
rect 236644 228404 236696 228410
rect 236644 228346 236696 228352
rect 236656 196722 236684 228346
rect 296732 199442 296760 230588
rect 327092 228478 327120 230588
rect 356072 230574 356546 230602
rect 297364 228472 297416 228478
rect 297364 228414 297416 228420
rect 327080 228472 327132 228478
rect 327080 228414 327132 228420
rect 296720 199436 296772 199442
rect 296720 199378 296772 199384
rect 236644 196716 236696 196722
rect 236644 196658 236696 196664
rect 236000 196648 236052 196654
rect 236000 196590 236052 196596
rect 297376 195906 297404 228414
rect 356072 195974 356100 230574
rect 386524 228410 386552 230588
rect 387800 230444 387852 230450
rect 387800 230386 387852 230392
rect 387812 229094 387840 230386
rect 387720 229066 387840 229094
rect 386512 228404 386564 228410
rect 386512 228346 386564 228352
rect 387720 223718 387748 229066
rect 387800 224936 387852 224942
rect 387800 224878 387852 224884
rect 384948 223712 385000 223718
rect 384948 223654 385000 223660
rect 387708 223712 387760 223718
rect 387708 223654 387760 223660
rect 384960 219502 384988 223654
rect 387064 223576 387116 223582
rect 387064 223518 387116 223524
rect 385040 220516 385092 220522
rect 385040 220458 385092 220464
rect 381360 219496 381412 219502
rect 381360 219438 381412 219444
rect 384948 219496 385000 219502
rect 384948 219438 385000 219444
rect 380900 213920 380952 213926
rect 380900 213862 380952 213868
rect 378784 213648 378836 213654
rect 378784 213590 378836 213596
rect 378140 211676 378192 211682
rect 378140 211618 378192 211624
rect 378152 207074 378180 211618
rect 378060 207046 378180 207074
rect 378060 204678 378088 207046
rect 375748 204672 375800 204678
rect 375748 204614 375800 204620
rect 378048 204672 378100 204678
rect 378048 204614 378100 204620
rect 375760 203590 375788 204614
rect 366364 203584 366416 203590
rect 366364 203526 366416 203532
rect 375748 203584 375800 203590
rect 375748 203526 375800 203532
rect 366376 197402 366404 203526
rect 378796 203046 378824 213590
rect 380912 211682 380940 213862
rect 381372 213654 381400 219438
rect 384304 218136 384356 218142
rect 384304 218078 384356 218084
rect 381360 213648 381412 213654
rect 381360 213590 381412 213596
rect 380900 211676 380952 211682
rect 380900 211618 380952 211624
rect 382924 206304 382976 206310
rect 382924 206246 382976 206252
rect 377128 203040 377180 203046
rect 377128 202982 377180 202988
rect 378784 203040 378836 203046
rect 378784 202982 378836 202988
rect 377140 200802 377168 202982
rect 375380 200796 375432 200802
rect 375380 200738 375432 200744
rect 377128 200796 377180 200802
rect 377128 200738 377180 200744
rect 375392 200114 375420 200738
rect 375300 200086 375420 200114
rect 364984 197396 365036 197402
rect 364984 197338 365036 197344
rect 366364 197396 366416 197402
rect 366364 197338 366416 197344
rect 356060 195968 356112 195974
rect 356060 195910 356112 195916
rect 297364 195900 297416 195906
rect 297364 195842 297416 195848
rect 217324 193860 217376 193866
rect 217324 193802 217376 193808
rect 188344 85536 188396 85542
rect 188344 85478 188396 85484
rect 185584 84176 185636 84182
rect 185584 84118 185636 84124
rect 184204 82816 184256 82822
rect 184204 82758 184256 82764
rect 178682 80880 178738 80889
rect 178682 80815 178738 80824
rect 178682 78704 178738 78713
rect 178682 78639 178738 78648
rect 178592 72072 178644 72078
rect 178592 72014 178644 72020
rect 178696 46918 178724 78639
rect 195980 75336 196032 75342
rect 195980 75278 196032 75284
rect 178684 46912 178736 46918
rect 178684 46854 178736 46860
rect 175556 33108 175608 33114
rect 175556 33050 175608 33056
rect 176660 32972 176712 32978
rect 176660 32914 176712 32920
rect 173898 32736 173954 32745
rect 173898 32671 173954 32680
rect 172518 25664 172574 25673
rect 172518 25599 172574 25608
rect 172532 16574 172560 25599
rect 172532 16546 172744 16574
rect 171784 15972 171836 15978
rect 171784 15914 171836 15920
rect 169116 12300 169168 12306
rect 169116 12242 169168 12248
rect 169024 6452 169076 6458
rect 169024 6394 169076 6400
rect 168196 3800 168248 3806
rect 168196 3742 168248 3748
rect 167736 3732 167788 3738
rect 167736 3674 167788 3680
rect 169128 3670 169156 12242
rect 170312 10872 170364 10878
rect 170312 10814 170364 10820
rect 169666 8120 169722 8129
rect 169666 8055 169722 8064
rect 168380 3664 168432 3670
rect 168380 3606 168432 3612
rect 169116 3664 169168 3670
rect 169116 3606 169168 3612
rect 167460 3392 167512 3398
rect 167460 3334 167512 3340
rect 168392 480 168420 3606
rect 169680 3330 169708 8055
rect 169576 3324 169628 3330
rect 169576 3266 169628 3272
rect 169668 3324 169720 3330
rect 169668 3266 169720 3272
rect 169588 480 169616 3266
rect 130538 326 131068 354
rect 130538 -960 130650 326
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170324 354 170352 10814
rect 171968 8900 172020 8906
rect 171968 8842 172020 8848
rect 171980 480 172008 8842
rect 170742 354 170854 480
rect 170324 326 170854 354
rect 170742 -960 170854 326
rect 171938 -960 172050 480
rect 172716 354 172744 16546
rect 173134 354 173246 480
rect 172716 326 173246 354
rect 173912 354 173940 32671
rect 176672 11694 176700 32914
rect 180800 32904 180852 32910
rect 180800 32846 180852 32852
rect 179420 25492 179472 25498
rect 179420 25434 179472 25440
rect 176752 25424 176804 25430
rect 176752 25366 176804 25372
rect 176660 11688 176712 11694
rect 176660 11630 176712 11636
rect 176764 6914 176792 25366
rect 179432 16574 179460 25434
rect 180812 16574 180840 32846
rect 184940 32836 184992 32842
rect 184940 32778 184992 32784
rect 183560 26240 183612 26246
rect 183560 26182 183612 26188
rect 183572 16574 183600 26182
rect 179432 16546 180288 16574
rect 180812 16546 181024 16574
rect 183572 16546 183784 16574
rect 177856 11688 177908 11694
rect 177856 11630 177908 11636
rect 176672 6886 176792 6914
rect 175464 3324 175516 3330
rect 175464 3266 175516 3272
rect 175476 480 175504 3266
rect 176672 480 176700 6886
rect 177868 480 177896 11630
rect 179052 9648 179104 9654
rect 179052 9590 179104 9596
rect 179064 480 179092 9590
rect 180260 480 180288 16546
rect 174238 354 174350 480
rect 173912 326 174350 354
rect 173134 -960 173246 326
rect 174238 -960 174350 326
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 180996 354 181024 16546
rect 182548 3256 182600 3262
rect 182548 3198 182600 3204
rect 182560 480 182588 3198
rect 183756 480 183784 16546
rect 184952 480 184980 32778
rect 194600 32768 194652 32774
rect 194600 32710 194652 32716
rect 187698 32600 187754 32609
rect 187698 32535 187754 32544
rect 186320 27532 186372 27538
rect 186320 27474 186372 27480
rect 186332 16574 186360 27474
rect 187712 16574 187740 32535
rect 191838 32464 191894 32473
rect 191838 32399 191894 32408
rect 190458 27160 190514 27169
rect 190458 27095 190514 27104
rect 186332 16546 186912 16574
rect 187712 16546 188568 16574
rect 186136 9580 186188 9586
rect 186136 9522 186188 9528
rect 186148 480 186176 9522
rect 181414 354 181526 480
rect 180996 326 181526 354
rect 181414 -960 181526 326
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 186884 354 186912 16546
rect 188540 480 188568 16546
rect 189724 4140 189776 4146
rect 189724 4082 189776 4088
rect 189736 480 189764 4082
rect 187302 354 187414 480
rect 186884 326 187414 354
rect 187302 -960 187414 326
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190472 354 190500 27095
rect 191852 16574 191880 32399
rect 193220 27600 193272 27606
rect 193220 27542 193272 27548
rect 191852 16546 192064 16574
rect 192036 480 192064 16546
rect 193232 3330 193260 27542
rect 194612 16574 194640 32710
rect 195992 16574 196020 75278
rect 207020 73228 207072 73234
rect 207020 73170 207072 73176
rect 198740 32700 198792 32706
rect 198740 32642 198792 32648
rect 197360 27464 197412 27470
rect 197360 27406 197412 27412
rect 197372 16574 197400 27406
rect 194612 16546 195192 16574
rect 195992 16546 196848 16574
rect 197372 16546 197952 16574
rect 193310 4720 193366 4729
rect 193310 4655 193366 4664
rect 193220 3324 193272 3330
rect 193220 3266 193272 3272
rect 193324 2394 193352 4655
rect 194416 3324 194468 3330
rect 194416 3266 194468 3272
rect 193232 2366 193352 2394
rect 193232 480 193260 2366
rect 194428 480 194456 3266
rect 190798 354 190910 480
rect 190472 326 190910 354
rect 190798 -960 190910 326
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195164 354 195192 16546
rect 196820 480 196848 16546
rect 197924 480 197952 16546
rect 195582 354 195694 480
rect 195164 326 195694 354
rect 195582 -960 195694 326
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 198752 354 198780 32642
rect 205640 32632 205692 32638
rect 205640 32574 205692 32580
rect 201500 27328 201552 27334
rect 201500 27270 201552 27276
rect 200304 10804 200356 10810
rect 200304 10746 200356 10752
rect 200316 480 200344 10746
rect 201512 480 201540 27270
rect 204260 27260 204312 27266
rect 204260 27202 204312 27208
rect 204272 16574 204300 27202
rect 205652 16574 205680 32574
rect 204272 16546 205128 16574
rect 205652 16546 206232 16574
rect 203432 10736 203484 10742
rect 203432 10678 203484 10684
rect 202696 5228 202748 5234
rect 202696 5170 202748 5176
rect 202708 480 202736 5170
rect 199078 354 199190 480
rect 198752 326 199190 354
rect 199078 -960 199190 326
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203444 354 203472 10678
rect 205100 480 205128 16546
rect 206204 480 206232 16546
rect 203862 354 203974 480
rect 203444 326 203974 354
rect 203862 -960 203974 326
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207032 354 207060 73170
rect 217336 72962 217364 193802
rect 358544 170400 358596 170406
rect 358544 170342 358596 170348
rect 358556 167074 358584 170342
rect 364996 169114 365024 197338
rect 375300 194410 375328 200086
rect 382936 197402 382964 206246
rect 379520 197396 379572 197402
rect 379520 197338 379572 197344
rect 382924 197396 382976 197402
rect 382924 197338 382976 197344
rect 379532 195226 379560 197338
rect 376024 195220 376076 195226
rect 376024 195162 376076 195168
rect 379520 195220 379572 195226
rect 379520 195162 379572 195168
rect 371240 194404 371292 194410
rect 371240 194346 371292 194352
rect 375288 194404 375340 194410
rect 375288 194346 375340 194352
rect 371252 191894 371280 194346
rect 371240 191888 371292 191894
rect 371240 191830 371292 191836
rect 365076 191820 365128 191826
rect 365076 191762 365128 191768
rect 362960 169108 363012 169114
rect 362960 169050 363012 169056
rect 364984 169108 365036 169114
rect 364984 169050 365036 169056
rect 355324 167068 355376 167074
rect 355324 167010 355376 167016
rect 358544 167068 358596 167074
rect 358544 167010 358596 167016
rect 355336 157350 355364 167010
rect 362972 162926 363000 169050
rect 365088 165170 365116 191762
rect 376036 169046 376064 195162
rect 384316 182850 384344 218078
rect 385052 213994 385080 220458
rect 387076 218142 387104 223518
rect 387812 222306 387840 224878
rect 390388 223582 390416 231095
rect 394620 229158 394648 232047
rect 394712 230518 394740 232086
rect 394700 230512 394752 230518
rect 394700 230454 394752 230460
rect 391940 229152 391992 229158
rect 391940 229094 391992 229100
rect 394608 229152 394660 229158
rect 394608 229094 394660 229100
rect 391952 226386 391980 229094
rect 391860 226358 391980 226386
rect 391860 225010 391888 226358
rect 391848 225004 391900 225010
rect 391848 224946 391900 224952
rect 390376 223576 390428 223582
rect 390376 223518 390428 223524
rect 387720 222278 387840 222306
rect 387720 220522 387748 222278
rect 387708 220516 387760 220522
rect 387708 220458 387760 220464
rect 387064 218136 387116 218142
rect 387064 218078 387116 218084
rect 385040 213988 385092 213994
rect 385040 213930 385092 213936
rect 393320 209976 393372 209982
rect 393320 209918 393372 209924
rect 393332 206310 393360 209918
rect 393320 206304 393372 206310
rect 393320 206246 393372 206252
rect 376116 182844 376168 182850
rect 376116 182786 376168 182792
rect 384304 182844 384356 182850
rect 384304 182786 384356 182792
rect 376128 170406 376156 182786
rect 376116 170400 376168 170406
rect 376116 170342 376168 170348
rect 366364 169040 366416 169046
rect 366364 168982 366416 168988
rect 376024 169040 376076 169046
rect 376024 168982 376076 168988
rect 363604 165164 363656 165170
rect 363604 165106 363656 165112
rect 365076 165164 365128 165170
rect 365076 165106 365128 165112
rect 362960 162920 363012 162926
rect 362960 162862 363012 162868
rect 358452 162852 358504 162858
rect 358452 162794 358504 162800
rect 358464 157418 358492 162794
rect 356060 157412 356112 157418
rect 356060 157354 356112 157360
rect 358452 157412 358504 157418
rect 358452 157354 358504 157360
rect 352564 157344 352616 157350
rect 352564 157286 352616 157292
rect 355324 157344 355376 157350
rect 355324 157286 355376 157292
rect 349804 153196 349856 153202
rect 349804 153138 349856 153144
rect 349816 151094 349844 153138
rect 343640 151088 343692 151094
rect 343640 151030 343692 151036
rect 349804 151088 349856 151094
rect 349804 151030 349856 151036
rect 343652 147694 343680 151030
rect 341524 147688 341576 147694
rect 341524 147630 341576 147636
rect 343640 147688 343692 147694
rect 343640 147630 343692 147636
rect 341536 117298 341564 147630
rect 351184 146940 351236 146946
rect 351184 146882 351236 146888
rect 351196 139466 351224 146882
rect 347044 139460 347096 139466
rect 347044 139402 347096 139408
rect 351184 139460 351236 139466
rect 351184 139402 351236 139408
rect 342260 137624 342312 137630
rect 342260 137566 342312 137572
rect 342272 134570 342300 137566
rect 342260 134564 342312 134570
rect 342260 134506 342312 134512
rect 347056 131170 347084 139402
rect 352576 137630 352604 157286
rect 356072 153270 356100 157354
rect 356060 153264 356112 153270
rect 356060 153206 356112 153212
rect 363616 146946 363644 165106
rect 366376 148850 366404 168982
rect 363696 148844 363748 148850
rect 363696 148786 363748 148792
rect 366364 148844 366416 148850
rect 366364 148786 366416 148792
rect 363604 146940 363656 146946
rect 363604 146882 363656 146888
rect 352564 137624 352616 137630
rect 352564 137566 352616 137572
rect 363708 136338 363736 148786
rect 360844 136332 360896 136338
rect 360844 136274 360896 136280
rect 363696 136332 363748 136338
rect 363696 136274 363748 136280
rect 345664 131164 345716 131170
rect 345664 131106 345716 131112
rect 347044 131164 347096 131170
rect 347044 131106 347096 131112
rect 345676 124234 345704 131106
rect 344284 124228 344336 124234
rect 344284 124170 344336 124176
rect 345664 124228 345716 124234
rect 345664 124170 345716 124176
rect 338764 117292 338816 117298
rect 338764 117234 338816 117240
rect 341524 117292 341576 117298
rect 341524 117234 341576 117240
rect 338776 106826 338804 117234
rect 337016 106820 337068 106826
rect 337016 106762 337068 106768
rect 338764 106820 338816 106826
rect 338764 106762 338816 106768
rect 337028 104854 337056 106762
rect 344296 106282 344324 124170
rect 360856 124166 360884 136274
rect 358084 124160 358136 124166
rect 358084 124102 358136 124108
rect 360844 124160 360896 124166
rect 360844 124102 360896 124108
rect 358096 111110 358124 124102
rect 348424 111104 348476 111110
rect 348424 111046 348476 111052
rect 358084 111104 358136 111110
rect 358084 111046 358136 111052
rect 344284 106276 344336 106282
rect 344284 106218 344336 106224
rect 337016 104848 337068 104854
rect 337016 104790 337068 104796
rect 348436 95946 348464 111046
rect 341524 95940 341576 95946
rect 341524 95882 341576 95888
rect 348424 95940 348476 95946
rect 348424 95882 348476 95888
rect 341536 82142 341564 95882
rect 332600 82136 332652 82142
rect 332600 82078 332652 82084
rect 341524 82136 341576 82142
rect 341524 82078 341576 82084
rect 332612 79354 332640 82078
rect 324320 79348 324372 79354
rect 324320 79290 324372 79296
rect 332600 79348 332652 79354
rect 332600 79290 332652 79296
rect 249800 75200 249852 75206
rect 249800 75142 249852 75148
rect 217324 72956 217376 72962
rect 217324 72898 217376 72904
rect 231124 72888 231176 72894
rect 231124 72830 231176 72836
rect 226340 40724 226392 40730
rect 226340 40666 226392 40672
rect 212540 34468 212592 34474
rect 212540 34410 212592 34416
rect 209778 34096 209834 34105
rect 209778 34031 209834 34040
rect 208400 27396 208452 27402
rect 208400 27338 208452 27344
rect 208412 16574 208440 27338
rect 208412 16546 208624 16574
rect 208596 480 208624 16546
rect 209792 480 209820 34031
rect 211160 28144 211212 28150
rect 211160 28086 211212 28092
rect 211172 16574 211200 28086
rect 212552 16574 212580 34410
rect 216680 34400 216732 34406
rect 216680 34342 216732 34348
rect 215300 28212 215352 28218
rect 215300 28154 215352 28160
rect 211172 16546 211752 16574
rect 212552 16546 213408 16574
rect 210974 12200 211030 12209
rect 210974 12135 211030 12144
rect 210988 480 211016 12135
rect 207358 354 207470 480
rect 207032 326 207470 354
rect 207358 -960 207470 326
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 211724 354 211752 16546
rect 213380 480 213408 16546
rect 214472 12232 214524 12238
rect 214472 12174 214524 12180
rect 214484 480 214512 12174
rect 212142 354 212254 480
rect 211724 326 212254 354
rect 212142 -960 212254 326
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215312 354 215340 28154
rect 216692 16574 216720 34342
rect 219440 34332 219492 34338
rect 219440 34274 219492 34280
rect 218060 27192 218112 27198
rect 218060 27134 218112 27140
rect 216692 16546 216904 16574
rect 216876 480 216904 16546
rect 218072 11694 218100 27134
rect 219452 16574 219480 34274
rect 222200 28076 222252 28082
rect 222200 28018 222252 28024
rect 222212 16574 222240 28018
rect 223578 20224 223634 20233
rect 223578 20159 223634 20168
rect 219452 16546 220032 16574
rect 222212 16546 222792 16574
rect 218152 12164 218204 12170
rect 218152 12106 218204 12112
rect 218060 11688 218112 11694
rect 218060 11630 218112 11636
rect 218164 6914 218192 12106
rect 219256 11688 219308 11694
rect 219256 11630 219308 11636
rect 218072 6886 218192 6914
rect 218072 480 218100 6886
rect 219268 480 219296 11630
rect 215638 354 215750 480
rect 215312 326 215750 354
rect 215638 -960 215750 326
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220004 354 220032 16546
rect 221096 12096 221148 12102
rect 221096 12038 221148 12044
rect 220422 354 220534 480
rect 220004 326 220534 354
rect 221108 354 221136 12038
rect 222764 480 222792 16546
rect 221526 354 221638 480
rect 221108 326 221638 354
rect 220422 -960 220534 326
rect 221526 -960 221638 326
rect 222722 -960 222834 480
rect 223592 354 223620 20159
rect 225142 12880 225198 12889
rect 225142 12815 225198 12824
rect 225156 480 225184 12815
rect 226352 3330 226380 40666
rect 229100 28960 229152 28966
rect 229100 28902 229152 28908
rect 229112 16574 229140 28902
rect 231136 20262 231164 72830
rect 239220 72820 239272 72826
rect 239220 72762 239272 72768
rect 239232 68338 239260 72762
rect 239220 68332 239272 68338
rect 239220 68274 239272 68280
rect 234620 34264 234672 34270
rect 234620 34206 234672 34212
rect 233240 27124 233292 27130
rect 233240 27066 233292 27072
rect 230480 20256 230532 20262
rect 230480 20198 230532 20204
rect 231124 20256 231176 20262
rect 231124 20198 231176 20204
rect 230492 16574 230520 20198
rect 233252 16574 233280 27066
rect 229112 16546 229416 16574
rect 230492 16546 231072 16574
rect 233252 16546 233464 16574
rect 226430 6896 226486 6905
rect 226430 6831 226486 6840
rect 226340 3324 226392 3330
rect 226340 3266 226392 3272
rect 226444 3210 226472 6831
rect 228730 6760 228786 6769
rect 228730 6695 228786 6704
rect 227536 3324 227588 3330
rect 227536 3266 227588 3272
rect 226352 3182 226472 3210
rect 226352 480 226380 3182
rect 227548 480 227576 3266
rect 228744 480 228772 6695
rect 223918 354 224030 480
rect 223592 326 224030 354
rect 223918 -960 224030 326
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229388 354 229416 16546
rect 231044 480 231072 16546
rect 231860 13456 231912 13462
rect 231860 13398 231912 13404
rect 229806 354 229918 480
rect 229388 326 229918 354
rect 229806 -960 229918 326
rect 231002 -960 231114 480
rect 231872 354 231900 13398
rect 233436 480 233464 16546
rect 234632 480 234660 34206
rect 248420 34196 248472 34202
rect 248420 34138 248472 34144
rect 241518 33960 241574 33969
rect 241518 33895 241574 33904
rect 240140 28824 240192 28830
rect 240140 28766 240192 28772
rect 236000 26172 236052 26178
rect 236000 26114 236052 26120
rect 236012 16574 236040 26114
rect 237380 20460 237432 20466
rect 237380 20402 237432 20408
rect 237392 16574 237420 20402
rect 236012 16546 236592 16574
rect 237392 16546 237696 16574
rect 235816 6724 235868 6730
rect 235816 6666 235868 6672
rect 235828 480 235856 6666
rect 232198 354 232310 480
rect 231872 326 232310 354
rect 232198 -960 232310 326
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236564 354 236592 16546
rect 236982 354 237094 480
rect 236564 326 237094 354
rect 237668 354 237696 16546
rect 239312 13388 239364 13394
rect 239312 13330 239364 13336
rect 239324 480 239352 13330
rect 238086 354 238198 480
rect 237668 326 238198 354
rect 236982 -960 237094 326
rect 238086 -960 238198 326
rect 239282 -960 239394 480
rect 240152 354 240180 28766
rect 241532 16574 241560 33895
rect 242900 28892 242952 28898
rect 242900 28834 242952 28840
rect 241532 16546 241744 16574
rect 241716 480 241744 16546
rect 242912 11694 242940 28834
rect 247040 28756 247092 28762
rect 247040 28698 247092 28704
rect 244278 20088 244334 20097
rect 244278 20023 244334 20032
rect 244292 16574 244320 20023
rect 247052 16574 247080 28698
rect 244292 16546 245240 16574
rect 247052 16546 247632 16574
rect 242990 13696 243046 13705
rect 242990 13631 243046 13640
rect 242900 11688 242952 11694
rect 242900 11630 242952 11636
rect 243004 6914 243032 13631
rect 244096 11688 244148 11694
rect 244096 11630 244148 11636
rect 242912 6886 243032 6914
rect 242912 480 242940 6886
rect 244108 480 244136 11630
rect 245212 480 245240 16546
rect 246394 6624 246450 6633
rect 246394 6559 246450 6568
rect 246408 480 246436 6559
rect 247604 480 247632 16546
rect 240478 354 240590 480
rect 240152 326 240590 354
rect 240478 -960 240590 326
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248432 354 248460 34138
rect 249812 16574 249840 75142
rect 259460 75132 259512 75138
rect 259460 75074 259512 75080
rect 259368 72752 259420 72758
rect 259368 72694 259420 72700
rect 259380 71058 259408 72694
rect 259368 71052 259420 71058
rect 259368 70994 259420 71000
rect 255320 34128 255372 34134
rect 255320 34070 255372 34076
rect 251180 28620 251232 28626
rect 251180 28562 251232 28568
rect 249812 16546 250024 16574
rect 249996 480 250024 16546
rect 251192 480 251220 28562
rect 253940 24812 253992 24818
rect 253940 24754 253992 24760
rect 251272 19100 251324 19106
rect 251272 19042 251324 19048
rect 251284 16574 251312 19042
rect 253952 16574 253980 24754
rect 255332 16574 255360 34070
rect 258080 28688 258132 28694
rect 258080 28630 258132 28636
rect 258092 16574 258120 28630
rect 251284 16546 252416 16574
rect 253952 16546 254256 16574
rect 255332 16546 255912 16574
rect 258092 16546 258304 16574
rect 252388 480 252416 16546
rect 253480 14952 253532 14958
rect 253480 14894 253532 14900
rect 253492 480 253520 14894
rect 248758 354 248870 480
rect 248432 326 248870 354
rect 248758 -960 248870 326
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254228 354 254256 16546
rect 255884 480 255912 16546
rect 256700 14884 256752 14890
rect 256700 14826 256752 14832
rect 254646 354 254758 480
rect 254228 326 254758 354
rect 254646 -960 254758 326
rect 255842 -960 255954 480
rect 256712 354 256740 14826
rect 258276 480 258304 16546
rect 259472 11694 259500 75074
rect 324332 75070 324360 79290
rect 324320 75064 324372 75070
rect 324320 75006 324372 75012
rect 320180 74996 320232 75002
rect 320180 74938 320232 74944
rect 284300 74316 284352 74322
rect 284300 74258 284352 74264
rect 269120 34060 269172 34066
rect 269120 34002 269172 34008
rect 262218 33824 262274 33833
rect 262218 33759 262274 33768
rect 260840 26104 260892 26110
rect 260840 26046 260892 26052
rect 259552 20392 259604 20398
rect 259552 20334 259604 20340
rect 259460 11688 259512 11694
rect 259460 11630 259512 11636
rect 259564 6914 259592 20334
rect 260852 16574 260880 26046
rect 262232 16574 262260 33759
rect 266360 32564 266412 32570
rect 266360 32506 266412 32512
rect 264980 28552 265032 28558
rect 264980 28494 265032 28500
rect 260852 16546 261800 16574
rect 262232 16546 262536 16574
rect 260656 11688 260708 11694
rect 260656 11630 260708 11636
rect 259472 6886 259592 6914
rect 259472 480 259500 6886
rect 260668 480 260696 11630
rect 261772 480 261800 16546
rect 257038 354 257150 480
rect 256712 326 257150 354
rect 257038 -960 257150 326
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262508 354 262536 16546
rect 264150 15192 264206 15201
rect 264150 15127 264206 15136
rect 264164 480 264192 15127
rect 262926 354 263038 480
rect 262508 326 263038 354
rect 262926 -960 263038 326
rect 264122 -960 264234 480
rect 264992 354 265020 28494
rect 266372 16574 266400 32506
rect 269132 16574 269160 34002
rect 276020 33992 276072 33998
rect 276020 33934 276072 33940
rect 271880 28484 271932 28490
rect 271880 28426 271932 28432
rect 271892 16574 271920 28426
rect 273260 17672 273312 17678
rect 273260 17614 273312 17620
rect 266372 16546 266584 16574
rect 269132 16546 270080 16574
rect 271892 16546 272472 16574
rect 266556 480 266584 16546
rect 267740 14816 267792 14822
rect 267740 14758 267792 14764
rect 267752 480 267780 14758
rect 268844 8016 268896 8022
rect 268844 7958 268896 7964
rect 268856 480 268884 7958
rect 270052 480 270080 16546
rect 270776 14748 270828 14754
rect 270776 14690 270828 14696
rect 265318 354 265430 480
rect 264992 326 265430 354
rect 265318 -960 265430 326
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 270788 354 270816 14690
rect 272444 480 272472 16546
rect 271206 354 271318 480
rect 270788 326 271318 354
rect 271206 -960 271318 326
rect 272402 -960 272514 480
rect 273272 354 273300 17614
rect 274824 16448 274876 16454
rect 274824 16390 274876 16396
rect 274836 480 274864 16390
rect 276032 4146 276060 33934
rect 278778 27024 278834 27033
rect 278778 26959 278834 26968
rect 278792 16574 278820 26959
rect 282920 24744 282972 24750
rect 282920 24686 282972 24692
rect 282932 16574 282960 24686
rect 278792 16546 279096 16574
rect 282932 16546 283144 16574
rect 276112 10668 276164 10674
rect 276112 10610 276164 10616
rect 276020 4140 276072 4146
rect 276020 4082 276072 4088
rect 276124 3482 276152 10610
rect 278318 7984 278374 7993
rect 278318 7919 278374 7928
rect 276756 4140 276808 4146
rect 276756 4082 276808 4088
rect 276032 3454 276152 3482
rect 276032 480 276060 3454
rect 273598 354 273710 480
rect 273272 326 273710 354
rect 273598 -960 273710 326
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 276768 354 276796 4082
rect 278332 480 278360 7919
rect 277094 354 277206 480
rect 276768 326 277206 354
rect 277094 -960 277206 326
rect 278290 -960 278402 480
rect 279068 354 279096 16546
rect 280710 13560 280766 13569
rect 280710 13495 280766 13504
rect 280724 480 280752 13495
rect 281906 7848 281962 7857
rect 281906 7783 281962 7792
rect 281920 480 281948 7783
rect 283116 480 283144 16546
rect 284312 4146 284340 74258
rect 302240 74248 302292 74254
rect 302240 74190 302292 74196
rect 298098 35320 298154 35329
rect 298098 35255 298154 35264
rect 284392 33924 284444 33930
rect 284392 33866 284444 33872
rect 284300 4140 284352 4146
rect 284300 4082 284352 4088
rect 284404 3482 284432 33866
rect 291200 33856 291252 33862
rect 291200 33798 291252 33804
rect 291212 16574 291240 33798
rect 292580 26036 292632 26042
rect 292580 25978 292632 25984
rect 291212 16546 291424 16574
rect 287336 16380 287388 16386
rect 287336 16322 287388 16328
rect 286600 6656 286652 6662
rect 286600 6598 286652 6604
rect 285036 4140 285088 4146
rect 285036 4082 285088 4088
rect 284312 3454 284432 3482
rect 284312 480 284340 3454
rect 279486 354 279598 480
rect 279068 326 279598 354
rect 279486 -960 279598 326
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285048 354 285076 4082
rect 286612 480 286640 6598
rect 285374 354 285486 480
rect 285048 326 285486 354
rect 285374 -960 285486 326
rect 286570 -960 286682 480
rect 287348 354 287376 16322
rect 288992 16312 289044 16318
rect 288992 16254 289044 16260
rect 289004 480 289032 16254
rect 290188 7948 290240 7954
rect 290188 7890 290240 7896
rect 290200 480 290228 7890
rect 291396 480 291424 16546
rect 292592 4146 292620 25978
rect 295614 16280 295670 16289
rect 292672 16244 292724 16250
rect 295614 16215 295670 16224
rect 292672 16186 292724 16192
rect 292580 4140 292632 4146
rect 292580 4082 292632 4088
rect 292684 3482 292712 16186
rect 294880 10600 294932 10606
rect 294880 10542 294932 10548
rect 293316 4140 293368 4146
rect 293316 4082 293368 4088
rect 292592 3454 292712 3482
rect 292592 480 292620 3454
rect 287766 354 287878 480
rect 287348 326 287878 354
rect 287766 -960 287878 326
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293328 354 293356 4082
rect 294892 480 294920 10542
rect 293654 354 293766 480
rect 293328 326 293766 354
rect 293654 -960 293766 326
rect 294850 -960 294962 480
rect 295628 354 295656 16215
rect 297270 15056 297326 15065
rect 297270 14991 297326 15000
rect 297284 480 297312 14991
rect 296046 354 296158 480
rect 295628 326 296158 354
rect 296046 -960 296158 326
rect 297242 -960 297354 480
rect 298112 354 298140 35255
rect 300860 33788 300912 33794
rect 300860 33730 300912 33736
rect 299480 30252 299532 30258
rect 299480 30194 299532 30200
rect 299492 3330 299520 30194
rect 300872 16574 300900 33730
rect 302252 16574 302280 74190
rect 307760 35896 307812 35902
rect 307760 35838 307812 35844
rect 305000 35148 305052 35154
rect 305000 35090 305052 35096
rect 303620 30184 303672 30190
rect 303620 30126 303672 30132
rect 303632 16574 303660 30126
rect 305012 16574 305040 35090
rect 300872 16546 301544 16574
rect 302252 16546 303200 16574
rect 303632 16546 303936 16574
rect 305012 16546 305592 16574
rect 299662 9208 299718 9217
rect 299662 9143 299718 9152
rect 299480 3324 299532 3330
rect 299480 3266 299532 3272
rect 299676 480 299704 9143
rect 300768 3324 300820 3330
rect 300768 3266 300820 3272
rect 300780 480 300808 3266
rect 298438 354 298550 480
rect 298112 326 298550 354
rect 298438 -960 298550 326
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301516 354 301544 16546
rect 303172 480 303200 16546
rect 301934 354 302046 480
rect 301516 326 302046 354
rect 301934 -960 302046 326
rect 303130 -960 303242 480
rect 303908 354 303936 16546
rect 305564 480 305592 16546
rect 306748 9512 306800 9518
rect 306748 9454 306800 9460
rect 306760 480 306788 9454
rect 307772 3330 307800 35838
rect 311900 35828 311952 35834
rect 311900 35770 311952 35776
rect 307852 30320 307904 30326
rect 307852 30262 307904 30268
rect 307864 16574 307892 30262
rect 311912 16574 311940 35770
rect 318800 35760 318852 35766
rect 318800 35702 318852 35708
rect 314658 29608 314714 29617
rect 314658 29543 314714 29552
rect 312544 19032 312596 19038
rect 312544 18974 312596 18980
rect 307864 16546 307984 16574
rect 311912 16546 312216 16574
rect 307760 3324 307812 3330
rect 307760 3266 307812 3272
rect 307956 480 307984 16546
rect 310244 9444 310296 9450
rect 310244 9386 310296 9392
rect 309048 3324 309100 3330
rect 309048 3266 309100 3272
rect 309060 480 309088 3266
rect 310256 480 310284 9386
rect 311440 9376 311492 9382
rect 311440 9318 311492 9324
rect 311452 480 311480 9318
rect 304326 354 304438 480
rect 303908 326 304438 354
rect 304326 -960 304438 326
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312188 354 312216 16546
rect 312556 4146 312584 18974
rect 313832 10532 313884 10538
rect 313832 10474 313884 10480
rect 312544 4140 312596 4146
rect 312544 4082 312596 4088
rect 313844 480 313872 10474
rect 312606 354 312718 480
rect 312188 326 312718 354
rect 312606 -960 312718 326
rect 313802 -960 313914 480
rect 314672 354 314700 29543
rect 316038 17640 316094 17649
rect 316038 17575 316094 17584
rect 316052 3330 316080 17575
rect 318812 16574 318840 35702
rect 320192 16574 320220 74938
rect 338120 74928 338172 74934
rect 396736 74905 396764 378150
rect 396908 364404 396960 364410
rect 396908 364346 396960 364352
rect 396816 324352 396868 324358
rect 396816 324294 396868 324300
rect 338120 74870 338172 74876
rect 396722 74896 396778 74905
rect 324320 74180 324372 74186
rect 324320 74122 324372 74128
rect 322940 35692 322992 35698
rect 322940 35634 322992 35640
rect 318812 16546 319760 16574
rect 320192 16546 320496 16574
rect 316222 14920 316278 14929
rect 316222 14855 316278 14864
rect 316040 3324 316092 3330
rect 316040 3266 316092 3272
rect 316236 480 316264 14855
rect 318064 10464 318116 10470
rect 318064 10406 318116 10412
rect 317328 3324 317380 3330
rect 317328 3266 317380 3272
rect 317340 480 317368 3266
rect 314998 354 315110 480
rect 314672 326 315110 354
rect 314998 -960 315110 326
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 354 318104 10406
rect 319732 480 319760 16546
rect 318494 354 318606 480
rect 318076 326 318606 354
rect 318494 -960 318606 326
rect 319690 -960 319802 480
rect 320468 354 320496 16546
rect 322112 12028 322164 12034
rect 322112 11970 322164 11976
rect 322124 480 322152 11970
rect 320886 354 320998 480
rect 320468 326 320998 354
rect 320886 -960 320998 326
rect 322082 -960 322194 480
rect 322952 354 322980 35634
rect 324332 3210 324360 74122
rect 326344 58676 326396 58682
rect 326344 58618 326396 58624
rect 325700 35624 325752 35630
rect 325700 35566 325752 35572
rect 324412 13320 324464 13326
rect 324412 13262 324464 13268
rect 324424 3330 324452 13262
rect 325712 6914 325740 35566
rect 326356 16574 326384 58618
rect 336740 35556 336792 35562
rect 336740 35498 336792 35504
rect 332598 35184 332654 35193
rect 332598 35119 332654 35128
rect 329840 20324 329892 20330
rect 329840 20266 329892 20272
rect 327080 17604 327132 17610
rect 327080 17546 327132 17552
rect 327092 16574 327120 17546
rect 329852 16574 329880 20266
rect 326356 16546 326476 16574
rect 327092 16546 328040 16574
rect 329852 16546 330432 16574
rect 325712 6886 326384 6914
rect 324412 3324 324464 3330
rect 324412 3266 324464 3272
rect 325608 3324 325660 3330
rect 325608 3266 325660 3272
rect 324332 3182 324452 3210
rect 324424 480 324452 3182
rect 325620 480 325648 3266
rect 323278 354 323390 480
rect 322952 326 323390 354
rect 323278 -960 323390 326
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326356 354 326384 6886
rect 326448 3262 326476 16546
rect 326436 3256 326488 3262
rect 326436 3198 326488 3204
rect 328012 480 328040 16546
rect 328736 13252 328788 13258
rect 328736 13194 328788 13200
rect 326774 354 326886 480
rect 326356 326 326886 354
rect 326774 -960 326886 326
rect 327970 -960 328082 480
rect 328748 354 328776 13194
rect 330404 480 330432 16546
rect 331218 10432 331274 10441
rect 331218 10367 331274 10376
rect 329166 354 329278 480
rect 328748 326 329278 354
rect 329166 -960 329278 326
rect 330362 -960 330474 480
rect 331232 354 331260 10367
rect 332612 3330 332640 35119
rect 336752 16574 336780 35498
rect 338132 16574 338160 74870
rect 396828 74866 396856 324294
rect 396920 137562 396948 364346
rect 397092 311908 397144 311914
rect 397092 311850 397144 311856
rect 397000 271924 397052 271930
rect 397000 271866 397052 271872
rect 396908 137556 396960 137562
rect 396908 137498 396960 137504
rect 396722 74831 396778 74840
rect 396816 74860 396868 74866
rect 396816 74802 396868 74808
rect 397012 74798 397040 271866
rect 397104 137494 397132 311850
rect 397184 258120 397236 258126
rect 397184 258062 397236 258068
rect 397092 137488 397144 137494
rect 397092 137430 397144 137436
rect 397196 137426 397224 258062
rect 397184 137420 397236 137426
rect 397184 137362 397236 137368
rect 397000 74792 397052 74798
rect 397000 74734 397052 74740
rect 390560 74724 390612 74730
rect 390560 74666 390612 74672
rect 374000 74112 374052 74118
rect 374000 74054 374052 74060
rect 347780 35488 347832 35494
rect 347780 35430 347832 35436
rect 343640 27056 343692 27062
rect 343640 26998 343692 27004
rect 340880 22024 340932 22030
rect 340880 21966 340932 21972
rect 340892 16574 340920 21966
rect 343652 16574 343680 26998
rect 347792 16574 347820 35430
rect 354680 35420 354732 35426
rect 354680 35362 354732 35368
rect 350538 21584 350594 21593
rect 350538 21519 350594 21528
rect 350552 16574 350580 21519
rect 354692 16574 354720 35362
rect 357440 35352 357492 35358
rect 357440 35294 357492 35300
rect 336752 16546 337056 16574
rect 338132 16546 338712 16574
rect 340892 16546 341012 16574
rect 343652 16546 344600 16574
rect 347792 16546 348096 16574
rect 350552 16546 351224 16574
rect 354692 16546 355272 16574
rect 332690 14784 332746 14793
rect 332690 14719 332746 14728
rect 332600 3324 332652 3330
rect 332600 3266 332652 3272
rect 332704 480 332732 14719
rect 334622 10296 334678 10305
rect 334622 10231 334678 10240
rect 333888 3324 333940 3330
rect 333888 3266 333940 3272
rect 333900 480 333928 3266
rect 331558 354 331670 480
rect 331232 326 331670 354
rect 331558 -960 331670 326
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 354 334664 10231
rect 336280 7880 336332 7886
rect 336280 7822 336332 7828
rect 336292 480 336320 7822
rect 335054 354 335166 480
rect 334636 326 335166 354
rect 335054 -960 335166 326
rect 336250 -960 336362 480
rect 337028 354 337056 16546
rect 338684 480 338712 16546
rect 339868 9308 339920 9314
rect 339868 9250 339920 9256
rect 339880 480 339908 9250
rect 340984 480 341012 16546
rect 342904 11960 342956 11966
rect 342904 11902 342956 11908
rect 342168 9240 342220 9246
rect 342168 9182 342220 9188
rect 342180 480 342208 9182
rect 337446 354 337558 480
rect 337028 326 337558 354
rect 337446 -960 337558 326
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342916 354 342944 11902
rect 344572 480 344600 16546
rect 346952 16176 347004 16182
rect 346952 16118 347004 16124
rect 345296 11892 345348 11898
rect 345296 11834 345348 11840
rect 343334 354 343446 480
rect 342916 326 343446 354
rect 343334 -960 343446 326
rect 344530 -960 344642 480
rect 345308 354 345336 11834
rect 346964 480 346992 16118
rect 348068 480 348096 16546
rect 349158 16144 349214 16153
rect 349158 16079 349214 16088
rect 349172 3262 349200 16079
rect 349250 12064 349306 12073
rect 349250 11999 349306 12008
rect 349160 3256 349212 3262
rect 349160 3198 349212 3204
rect 349264 480 349292 11999
rect 350448 3256 350500 3262
rect 350448 3198 350500 3204
rect 350460 480 350488 3198
rect 345726 354 345838 480
rect 345308 326 345838 354
rect 345726 -960 345838 326
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351196 354 351224 16546
rect 353576 16108 353628 16114
rect 353576 16050 353628 16056
rect 352838 11928 352894 11937
rect 352838 11863 352894 11872
rect 352852 480 352880 11863
rect 351614 354 351726 480
rect 351196 326 351726 354
rect 351614 -960 351726 326
rect 352810 -960 352922 480
rect 353588 354 353616 16050
rect 355244 480 355272 16546
rect 356336 11824 356388 11830
rect 356336 11766 356388 11772
rect 356348 480 356376 11766
rect 357452 3262 357480 35294
rect 368480 35284 368532 35290
rect 368480 35226 368532 35232
rect 367098 26888 367154 26897
rect 367098 26823 367154 26832
rect 357532 25968 357584 25974
rect 357532 25910 357584 25916
rect 357440 3256 357492 3262
rect 357440 3198 357492 3204
rect 357544 480 357572 25910
rect 361580 21956 361632 21962
rect 361580 21898 361632 21904
rect 358820 18964 358872 18970
rect 358820 18906 358872 18912
rect 358832 16574 358860 18906
rect 361592 16574 361620 21898
rect 367112 16574 367140 26823
rect 368492 16574 368520 35226
rect 371240 28416 371292 28422
rect 371240 28358 371292 28364
rect 358832 16546 359504 16574
rect 361592 16546 361896 16574
rect 367112 16546 367784 16574
rect 368492 16546 369440 16574
rect 358728 3256 358780 3262
rect 358728 3198 358780 3204
rect 358740 480 358768 3198
rect 354006 354 354118 480
rect 353588 326 354118 354
rect 354006 -960 354118 326
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359476 354 359504 16546
rect 361120 14680 361172 14686
rect 361120 14622 361172 14628
rect 361132 480 361160 14622
rect 359894 354 360006 480
rect 359476 326 360006 354
rect 359894 -960 360006 326
rect 361090 -960 361202 480
rect 361868 354 361896 16546
rect 365718 13424 365774 13433
rect 365718 13359 365774 13368
rect 363512 13184 363564 13190
rect 363512 13126 363564 13132
rect 363524 480 363552 13126
rect 364616 5160 364668 5166
rect 364616 5102 364668 5108
rect 364628 480 364656 5102
rect 365732 3262 365760 13359
rect 365810 11792 365866 11801
rect 365810 11727 365866 11736
rect 365720 3256 365772 3262
rect 365720 3198 365772 3204
rect 365824 480 365852 11727
rect 367008 3256 367060 3262
rect 367008 3198 367060 3204
rect 367020 480 367048 3198
rect 362286 354 362398 480
rect 361868 326 362398 354
rect 362286 -960 362398 326
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 367756 354 367784 16546
rect 369412 480 369440 16546
rect 370134 13288 370190 13297
rect 370134 13223 370190 13232
rect 368174 354 368286 480
rect 367756 326 368286 354
rect 368174 -960 368286 326
rect 369370 -960 369482 480
rect 370148 354 370176 13223
rect 370566 354 370678 480
rect 370148 326 370678 354
rect 371252 354 371280 28358
rect 372620 25900 372672 25906
rect 372620 25842 372672 25848
rect 372632 16574 372660 25842
rect 372632 16546 372936 16574
rect 372908 480 372936 16546
rect 374012 3074 374040 74054
rect 382280 35216 382332 35222
rect 382280 35158 382332 35164
rect 374092 30116 374144 30122
rect 374092 30058 374144 30064
rect 374104 3262 374132 30058
rect 375380 28348 375432 28354
rect 375380 28290 375432 28296
rect 375392 16574 375420 28290
rect 376760 18896 376812 18902
rect 376760 18838 376812 18844
rect 376772 16574 376800 18838
rect 380900 18828 380952 18834
rect 380900 18770 380952 18776
rect 380912 16574 380940 18770
rect 375392 16546 376064 16574
rect 376772 16546 377720 16574
rect 380912 16546 381216 16574
rect 374092 3256 374144 3262
rect 374092 3198 374144 3204
rect 375288 3256 375340 3262
rect 375288 3198 375340 3204
rect 374012 3046 374132 3074
rect 374104 480 374132 3046
rect 375300 480 375328 3198
rect 371670 354 371782 480
rect 371252 326 371782 354
rect 370566 -960 370678 326
rect 371670 -960 371782 326
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376036 354 376064 16546
rect 377692 480 377720 16546
rect 378416 13116 378468 13122
rect 378416 13058 378468 13064
rect 376454 354 376566 480
rect 376036 326 376566 354
rect 376454 -960 376566 326
rect 377650 -960 377762 480
rect 378428 354 378456 13058
rect 379980 6588 380032 6594
rect 379980 6530 380032 6536
rect 379992 480 380020 6530
rect 381188 480 381216 16546
rect 382292 3262 382320 35158
rect 382372 30048 382424 30054
rect 382372 29990 382424 29996
rect 382280 3256 382332 3262
rect 382280 3198 382332 3204
rect 382384 480 382412 29990
rect 389180 29980 389232 29986
rect 389180 29922 389232 29928
rect 386418 24440 386474 24449
rect 386418 24375 386474 24384
rect 386432 16574 386460 24375
rect 389192 16574 389220 29922
rect 386432 16546 386736 16574
rect 389192 16546 389496 16574
rect 384304 14612 384356 14618
rect 384304 14554 384356 14560
rect 383568 3256 383620 3262
rect 383568 3198 383620 3204
rect 383580 480 383608 3198
rect 378846 354 378958 480
rect 378428 326 378958 354
rect 378846 -960 378958 326
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384316 354 384344 14554
rect 385958 6488 386014 6497
rect 385958 6423 386014 6432
rect 385972 480 386000 6423
rect 384734 354 384846 480
rect 384316 326 384846 354
rect 384734 -960 384846 326
rect 385930 -960 386042 480
rect 386708 354 386736 16546
rect 387798 14648 387854 14657
rect 387798 14583 387854 14592
rect 387126 354 387238 480
rect 386708 326 387238 354
rect 387812 354 387840 14583
rect 389468 480 389496 16546
rect 390572 3262 390600 74666
rect 397472 73030 397500 703520
rect 410524 700392 410576 700398
rect 410524 700334 410576 700340
rect 409144 700324 409196 700330
rect 409144 700266 409196 700272
rect 407764 670744 407816 670750
rect 407764 670686 407816 670692
rect 406384 616888 406436 616894
rect 406384 616830 406436 616836
rect 405004 563100 405056 563106
rect 405004 563042 405056 563048
rect 397552 534132 397604 534138
rect 397552 534074 397604 534080
rect 397564 209982 397592 534074
rect 403624 510672 403676 510678
rect 403624 510614 403676 510620
rect 400864 456816 400916 456822
rect 400864 456758 400916 456764
rect 399576 444440 399628 444446
rect 399576 444382 399628 444388
rect 398104 418192 398156 418198
rect 398104 418134 398156 418140
rect 397552 209976 397604 209982
rect 397552 209918 397604 209924
rect 398116 137358 398144 418134
rect 399484 404388 399536 404394
rect 399484 404330 399536 404336
rect 398104 137352 398156 137358
rect 398104 137294 398156 137300
rect 399496 91050 399524 404330
rect 399588 187678 399616 444382
rect 399576 187672 399628 187678
rect 399576 187614 399628 187620
rect 400876 92478 400904 456758
rect 403636 93838 403664 510614
rect 405016 95198 405044 563042
rect 406396 97986 406424 616830
rect 407776 99346 407804 670686
rect 409156 100706 409184 700266
rect 410536 102134 410564 700334
rect 412652 135998 412680 703582
rect 413480 703474 413508 703582
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 413664 703474 413692 703520
rect 413480 703446 413692 703474
rect 429856 700466 429884 703520
rect 413284 700460 413336 700466
rect 413284 700402 413336 700408
rect 429844 700460 429896 700466
rect 429844 700402 429896 700408
rect 412640 135992 412692 135998
rect 412640 135934 412692 135940
rect 413296 103494 413324 700402
rect 418804 351960 418856 351966
rect 418804 351902 418856 351908
rect 417424 298172 417476 298178
rect 417424 298114 417476 298120
rect 414664 244316 414716 244322
rect 414664 244258 414716 244264
rect 413284 103488 413336 103494
rect 413284 103430 413336 103436
rect 410524 102128 410576 102134
rect 410524 102070 410576 102076
rect 409144 100700 409196 100706
rect 409144 100642 409196 100648
rect 407764 99340 407816 99346
rect 407764 99282 407816 99288
rect 406384 97980 406436 97986
rect 406384 97922 406436 97928
rect 405004 95192 405056 95198
rect 405004 95134 405056 95140
rect 403624 93832 403676 93838
rect 403624 93774 403676 93780
rect 400864 92472 400916 92478
rect 400864 92414 400916 92420
rect 399484 91044 399536 91050
rect 399484 90986 399536 90992
rect 414676 86970 414704 244258
rect 417436 88330 417464 298114
rect 418816 89690 418844 351902
rect 418804 89684 418856 89690
rect 418804 89626 418856 89632
rect 417424 88324 417476 88330
rect 417424 88266 417476 88272
rect 414664 86964 414716 86970
rect 414664 86906 414716 86912
rect 408500 74044 408552 74050
rect 408500 73986 408552 73992
rect 397460 73024 397512 73030
rect 397460 72966 397512 72972
rect 405002 72720 405058 72729
rect 405002 72655 405058 72664
rect 390652 36712 390704 36718
rect 390652 36654 390704 36660
rect 390560 3256 390612 3262
rect 390560 3198 390612 3204
rect 390664 480 390692 36654
rect 397460 36644 397512 36650
rect 397460 36586 397512 36592
rect 394700 20188 394752 20194
rect 394700 20130 394752 20136
rect 394712 16574 394740 20130
rect 397472 16574 397500 36586
rect 398840 20120 398892 20126
rect 398840 20062 398892 20068
rect 394712 16546 395384 16574
rect 397472 16546 397776 16574
rect 393044 9172 393096 9178
rect 393044 9114 393096 9120
rect 391848 3256 391900 3262
rect 391848 3198 391900 3204
rect 391860 480 391888 3198
rect 393056 480 393084 9114
rect 394240 3392 394292 3398
rect 394240 3334 394292 3340
rect 394252 480 394280 3334
rect 395356 480 395384 16546
rect 396540 6520 396592 6526
rect 396540 6462 396592 6468
rect 396552 480 396580 6462
rect 397748 480 397776 16546
rect 398852 3210 398880 20062
rect 402518 14512 402574 14521
rect 402518 14447 402574 14456
rect 398932 10396 398984 10402
rect 398932 10338 398984 10344
rect 398944 3398 398972 10338
rect 401324 4072 401376 4078
rect 401324 4014 401376 4020
rect 398932 3392 398984 3398
rect 398932 3334 398984 3340
rect 400128 3392 400180 3398
rect 400128 3334 400180 3340
rect 398852 3182 398972 3210
rect 398944 480 398972 3182
rect 400140 480 400168 3334
rect 401336 480 401364 4014
rect 402532 480 402560 14447
rect 403622 11656 403678 11665
rect 403622 11591 403678 11600
rect 403636 480 403664 11591
rect 404818 5536 404874 5545
rect 404818 5471 404874 5480
rect 404832 480 404860 5471
rect 405016 5166 405044 72655
rect 407212 24676 407264 24682
rect 407212 24618 407264 24624
rect 406014 16008 406070 16017
rect 406014 15943 406070 15952
rect 405004 5160 405056 5166
rect 405004 5102 405056 5108
rect 406028 480 406056 15943
rect 407224 480 407252 24618
rect 408512 16574 408540 73986
rect 462332 73982 462360 703520
rect 478524 702434 478552 703520
rect 477512 702406 478552 702434
rect 477512 142866 477540 702406
rect 494808 700398 494836 703520
rect 494796 700392 494848 700398
rect 494796 700334 494848 700340
rect 477500 142860 477552 142866
rect 477500 142802 477552 142808
rect 465172 74656 465224 74662
rect 465172 74598 465224 74604
rect 462320 73976 462372 73982
rect 462320 73918 462372 73924
rect 422300 72684 422352 72690
rect 422300 72626 422352 72632
rect 414020 25832 414072 25838
rect 414020 25774 414072 25780
rect 412640 20052 412692 20058
rect 412640 19994 412692 20000
rect 408512 16546 409184 16574
rect 408408 4004 408460 4010
rect 408408 3946 408460 3952
rect 408420 480 408448 3946
rect 388230 354 388342 480
rect 387812 326 388342 354
rect 387126 -960 387238 326
rect 388230 -960 388342 326
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409156 354 409184 16546
rect 410800 9104 410852 9110
rect 410800 9046 410852 9052
rect 410812 480 410840 9046
rect 411904 9036 411956 9042
rect 411904 8978 411956 8984
rect 411916 480 411944 8978
rect 409574 354 409686 480
rect 409156 326 409686 354
rect 409574 -960 409686 326
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 412652 354 412680 19994
rect 414032 16574 414060 25774
rect 420918 17504 420974 17513
rect 420918 17439 420974 17448
rect 414032 16546 414336 16574
rect 414308 480 414336 16546
rect 415492 16040 415544 16046
rect 415492 15982 415544 15988
rect 415400 3936 415452 3942
rect 415400 3878 415452 3884
rect 415412 1986 415440 3878
rect 415504 3398 415532 15982
rect 420182 15872 420238 15881
rect 420182 15807 420238 15816
rect 418526 13152 418582 13161
rect 418526 13087 418582 13096
rect 417884 7812 417936 7818
rect 417884 7754 417936 7760
rect 415492 3392 415544 3398
rect 415492 3334 415544 3340
rect 416688 3392 416740 3398
rect 416688 3334 416740 3340
rect 415412 1958 415532 1986
rect 415504 480 415532 1958
rect 416700 480 416728 3334
rect 417896 480 417924 7754
rect 413070 354 413182 480
rect 412652 326 413182 354
rect 413070 -960 413182 326
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418540 354 418568 13087
rect 420196 480 420224 15807
rect 418958 354 419070 480
rect 418540 326 419070 354
rect 418958 -960 419070 326
rect 420154 -960 420266 480
rect 420932 354 420960 17439
rect 422312 16574 422340 72626
rect 460940 68332 460992 68338
rect 460940 68274 460992 68280
rect 456800 36576 456852 36582
rect 456800 36518 456852 36524
rect 445022 31240 445078 31249
rect 445022 31175 445078 31184
rect 431960 29912 432012 29918
rect 431960 29854 432012 29860
rect 423680 26988 423732 26994
rect 423680 26930 423732 26936
rect 422312 16546 422616 16574
rect 422588 480 422616 16546
rect 423692 3398 423720 26930
rect 430580 21888 430632 21894
rect 430580 21830 430632 21836
rect 427820 17536 427872 17542
rect 427820 17478 427872 17484
rect 423770 17368 423826 17377
rect 423770 17303 423826 17312
rect 423680 3392 423732 3398
rect 423680 3334 423732 3340
rect 423784 480 423812 17303
rect 427832 16574 427860 17478
rect 430592 16574 430620 21830
rect 427832 16546 428504 16574
rect 430592 16546 430896 16574
rect 425704 14544 425756 14550
rect 425704 14486 425756 14492
rect 424968 3392 425020 3398
rect 424968 3334 425020 3340
rect 424980 480 425008 3334
rect 421350 354 421462 480
rect 420932 326 421462 354
rect 421350 -960 421462 326
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 425716 354 425744 14486
rect 427268 3868 427320 3874
rect 427268 3810 427320 3816
rect 427280 480 427308 3810
rect 428476 480 428504 16546
rect 429660 6452 429712 6458
rect 429660 6394 429712 6400
rect 429672 480 429700 6394
rect 430868 480 430896 16546
rect 431972 1714 432000 29854
rect 438860 29844 438912 29850
rect 438860 29786 438912 29792
rect 432052 21820 432104 21826
rect 432052 21762 432104 21768
rect 432064 1834 432092 21762
rect 433340 17468 433392 17474
rect 433340 17410 433392 17416
rect 433352 16574 433380 17410
rect 434720 17400 434772 17406
rect 434720 17342 434772 17348
rect 434732 16574 434760 17342
rect 437480 17332 437532 17338
rect 437480 17274 437532 17280
rect 433352 16546 434024 16574
rect 434732 16546 435128 16574
rect 432052 1828 432104 1834
rect 432052 1770 432104 1776
rect 433248 1828 433300 1834
rect 433248 1770 433300 1776
rect 431972 1686 432092 1714
rect 432064 480 432092 1686
rect 433260 480 433288 1770
rect 426134 354 426246 480
rect 425716 326 426246 354
rect 426134 -960 426246 326
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 433996 354 434024 16546
rect 434414 354 434526 480
rect 433996 326 434526 354
rect 435100 354 435128 16546
rect 436744 6384 436796 6390
rect 436744 6326 436796 6332
rect 436756 480 436784 6326
rect 435518 354 435630 480
rect 435100 326 435630 354
rect 434414 -960 434526 326
rect 435518 -960 435630 326
rect 436714 -960 436826 480
rect 437492 354 437520 17274
rect 438872 16574 438900 29786
rect 441620 29776 441672 29782
rect 441620 29718 441672 29724
rect 440238 21448 440294 21457
rect 440238 21383 440294 21392
rect 438872 16546 439176 16574
rect 439148 480 439176 16546
rect 440252 3210 440280 21383
rect 440330 17232 440386 17241
rect 440330 17167 440386 17176
rect 440344 3398 440372 17167
rect 441632 16574 441660 29718
rect 445036 16574 445064 31175
rect 445760 29708 445812 29714
rect 445760 29650 445812 29656
rect 441632 16546 442672 16574
rect 445036 16546 445156 16574
rect 440332 3392 440384 3398
rect 440332 3334 440384 3340
rect 441528 3392 441580 3398
rect 441528 3334 441580 3340
rect 440252 3182 440372 3210
rect 440344 480 440372 3182
rect 441540 480 441568 3334
rect 442644 480 442672 16546
rect 443368 15972 443420 15978
rect 443368 15914 443420 15920
rect 437910 354 438022 480
rect 437492 326 438022 354
rect 437910 -960 438022 326
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443380 354 443408 15914
rect 445128 3806 445156 16546
rect 445024 3800 445076 3806
rect 445024 3742 445076 3748
rect 445116 3800 445168 3806
rect 445116 3742 445168 3748
rect 445036 480 445064 3742
rect 443798 354 443910 480
rect 443380 326 443910 354
rect 443798 -960 443910 326
rect 444994 -960 445106 480
rect 445772 354 445800 29650
rect 452660 29640 452712 29646
rect 452660 29582 452712 29588
rect 447140 21752 447192 21758
rect 447140 21694 447192 21700
rect 447152 16574 447180 21694
rect 448520 21684 448572 21690
rect 448520 21626 448572 21632
rect 447152 16546 447456 16574
rect 447428 480 447456 16546
rect 448532 3210 448560 21626
rect 449900 20256 449952 20262
rect 449900 20198 449952 20204
rect 449912 16574 449940 20198
rect 451280 18760 451332 18766
rect 451280 18702 451332 18708
rect 451292 16574 451320 18702
rect 452672 16574 452700 29582
rect 454038 22808 454094 22817
rect 454038 22743 454094 22752
rect 449912 16546 450952 16574
rect 451292 16546 451688 16574
rect 452672 16546 453344 16574
rect 448612 10328 448664 10334
rect 448612 10270 448664 10276
rect 448624 3398 448652 10270
rect 448612 3392 448664 3398
rect 448612 3334 448664 3340
rect 449808 3392 449860 3398
rect 449808 3334 449860 3340
rect 448532 3182 448652 3210
rect 448624 480 448652 3182
rect 449820 480 449848 3334
rect 450924 480 450952 16546
rect 446190 354 446302 480
rect 445772 326 446302 354
rect 446190 -960 446302 326
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 451660 354 451688 16546
rect 453316 480 453344 16546
rect 452078 354 452190 480
rect 451660 326 452190 354
rect 452078 -960 452190 326
rect 453274 -960 453386 480
rect 454052 354 454080 22743
rect 455418 18864 455474 18873
rect 455418 18799 455474 18808
rect 455432 16574 455460 18799
rect 455432 16546 455736 16574
rect 455708 480 455736 16546
rect 456812 3398 456840 36518
rect 456890 25528 456946 25537
rect 456890 25463 456946 25472
rect 456800 3392 456852 3398
rect 456800 3334 456852 3340
rect 456904 480 456932 25463
rect 459560 23452 459612 23458
rect 459560 23394 459612 23400
rect 458178 18728 458234 18737
rect 458178 18663 458234 18672
rect 458192 16574 458220 18663
rect 459572 16574 459600 23394
rect 460952 16574 460980 68274
rect 463700 31748 463752 31754
rect 463700 31690 463752 31696
rect 463712 16574 463740 31690
rect 465184 16574 465212 74598
rect 527192 73914 527220 703520
rect 543476 702434 543504 703520
rect 542372 702406 543504 702434
rect 542372 137290 542400 702406
rect 559668 700330 559696 703520
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 580446 683904 580502 683913
rect 580446 683839 580502 683848
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580262 644056 580318 644065
rect 580262 643991 580318 644000
rect 579986 617536 580042 617545
rect 579986 617471 580042 617480
rect 580000 616894 580028 617471
rect 579988 616888 580040 616894
rect 579988 616830 580040 616836
rect 580170 564360 580226 564369
rect 580170 564295 580226 564304
rect 580184 563106 580212 564295
rect 580172 563100 580224 563106
rect 580172 563042 580224 563048
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 579802 511320 579858 511329
rect 579802 511255 579858 511264
rect 579816 510678 579844 511255
rect 579804 510672 579856 510678
rect 579804 510614 579856 510620
rect 579986 458144 580042 458153
rect 579986 458079 580042 458088
rect 580000 456822 580028 458079
rect 579988 456816 580040 456822
rect 579988 456758 580040 456764
rect 580078 444816 580134 444825
rect 580078 444751 580134 444760
rect 580092 444446 580120 444751
rect 580080 444440 580132 444446
rect 580080 444382 580132 444388
rect 580078 418296 580134 418305
rect 580078 418231 580134 418240
rect 580092 418198 580120 418231
rect 580080 418192 580132 418198
rect 580080 418134 580132 418140
rect 580078 404968 580134 404977
rect 580078 404903 580134 404912
rect 580092 404394 580120 404903
rect 580080 404388 580132 404394
rect 580080 404330 580132 404336
rect 580078 378448 580134 378457
rect 580078 378383 580134 378392
rect 580092 378214 580120 378383
rect 580080 378208 580132 378214
rect 580080 378150 580132 378156
rect 579802 365120 579858 365129
rect 579802 365055 579858 365064
rect 579816 364410 579844 365055
rect 579804 364404 579856 364410
rect 579804 364346 579856 364352
rect 580080 351960 580132 351966
rect 580078 351928 580080 351937
rect 580132 351928 580134 351937
rect 580078 351863 580134 351872
rect 580078 325272 580134 325281
rect 580078 325207 580134 325216
rect 580092 324358 580120 325207
rect 580080 324352 580132 324358
rect 580080 324294 580132 324300
rect 580078 312080 580134 312089
rect 580078 312015 580134 312024
rect 580092 311914 580120 312015
rect 580080 311908 580132 311914
rect 580080 311850 580132 311856
rect 580078 298752 580134 298761
rect 580078 298687 580134 298696
rect 580092 298178 580120 298687
rect 580080 298172 580132 298178
rect 580080 298114 580132 298120
rect 579802 272232 579858 272241
rect 579802 272167 579858 272176
rect 579816 271930 579844 272167
rect 579804 271924 579856 271930
rect 579804 271866 579856 271872
rect 579986 258904 580042 258913
rect 579986 258839 580042 258848
rect 580000 258126 580028 258839
rect 579988 258120 580040 258126
rect 579988 258062 580040 258068
rect 579986 245576 580042 245585
rect 579986 245511 580042 245520
rect 580000 244322 580028 245511
rect 579988 244316 580040 244322
rect 579988 244258 580040 244264
rect 580078 232384 580134 232393
rect 580078 232319 580134 232328
rect 579802 219056 579858 219065
rect 579802 218991 579858 219000
rect 579816 218074 579844 218991
rect 579804 218068 579856 218074
rect 579804 218010 579856 218016
rect 579986 205728 580042 205737
rect 579986 205663 579988 205672
rect 580040 205663 580042 205672
rect 579988 205634 580040 205640
rect 579894 192536 579950 192545
rect 579894 192471 579950 192480
rect 579802 165880 579858 165889
rect 579802 165815 579858 165824
rect 579816 165646 579844 165815
rect 579804 165640 579856 165646
rect 579804 165582 579856 165588
rect 579618 139360 579674 139369
rect 579618 139295 579674 139304
rect 579632 138038 579660 139295
rect 579620 138032 579672 138038
rect 579620 137974 579672 137980
rect 542360 137284 542412 137290
rect 542360 137226 542412 137232
rect 579710 126032 579766 126041
rect 579710 125967 579766 125976
rect 579724 125662 579752 125967
rect 579712 125656 579764 125662
rect 579712 125598 579764 125604
rect 562324 75948 562376 75954
rect 562324 75890 562376 75896
rect 527180 73908 527232 73914
rect 527180 73850 527232 73856
rect 550640 73840 550692 73846
rect 550640 73782 550692 73788
rect 471980 72616 472032 72622
rect 471980 72558 472032 72564
rect 480258 72584 480314 72593
rect 470600 31680 470652 31686
rect 470600 31622 470652 31628
rect 467840 26920 467892 26926
rect 467840 26862 467892 26868
rect 467852 16574 467880 26862
rect 469220 19984 469272 19990
rect 469220 19926 469272 19932
rect 469232 16574 469260 19926
rect 458192 16546 459232 16574
rect 459572 16546 459968 16574
rect 460952 16546 461624 16574
rect 463712 16546 464016 16574
rect 465184 16546 465856 16574
rect 467852 16546 468248 16574
rect 469232 16546 469904 16574
rect 458088 3392 458140 3398
rect 458088 3334 458140 3340
rect 458100 480 458128 3334
rect 459204 480 459232 16546
rect 454470 354 454582 480
rect 454052 326 454582 354
rect 454470 -960 454582 326
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459940 354 459968 16546
rect 461596 480 461624 16546
rect 462780 3732 462832 3738
rect 462780 3674 462832 3680
rect 462792 480 462820 3674
rect 463988 480 464016 16546
rect 465172 3664 465224 3670
rect 465172 3606 465224 3612
rect 465184 480 465212 3606
rect 460358 354 460470 480
rect 459940 326 460470 354
rect 460358 -960 460470 326
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 465828 354 465856 16546
rect 467472 14476 467524 14482
rect 467472 14418 467524 14424
rect 467484 480 467512 14418
rect 466246 354 466358 480
rect 465828 326 466358 354
rect 466246 -960 466358 326
rect 467442 -960 467554 480
rect 468220 354 468248 16546
rect 469876 480 469904 16546
rect 468638 354 468750 480
rect 468220 326 468750 354
rect 468638 -960 468750 326
rect 469834 -960 469946 480
rect 470612 354 470640 31622
rect 471992 16574 472020 72558
rect 480258 72519 480314 72528
rect 520924 72548 520976 72554
rect 474738 65512 474794 65521
rect 474738 65447 474794 65456
rect 473358 31104 473414 31113
rect 473358 31039 473414 31048
rect 471992 16546 472296 16574
rect 472268 480 472296 16546
rect 473372 3398 473400 31039
rect 473450 19952 473506 19961
rect 473450 19887 473506 19896
rect 473360 3392 473412 3398
rect 473360 3334 473412 3340
rect 473464 480 473492 19887
rect 474752 16574 474780 65447
rect 477500 31612 477552 31618
rect 477500 31554 477552 31560
rect 476118 21312 476174 21321
rect 476118 21247 476174 21256
rect 476132 16574 476160 21247
rect 477512 16574 477540 31554
rect 480272 16574 480300 72519
rect 520924 72490 520976 72496
rect 498198 72448 498254 72457
rect 498198 72383 498254 72392
rect 481640 31544 481692 31550
rect 481640 31486 481692 31492
rect 474752 16546 475792 16574
rect 476132 16546 476528 16574
rect 477512 16546 478184 16574
rect 480272 16546 480576 16574
rect 474188 3392 474240 3398
rect 474188 3334 474240 3340
rect 471030 354 471142 480
rect 470612 326 471142 354
rect 471030 -960 471142 326
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474200 354 474228 3334
rect 475764 480 475792 16546
rect 474526 354 474638 480
rect 474200 326 474638 354
rect 474526 -960 474638 326
rect 475722 -960 475834 480
rect 476500 354 476528 16546
rect 478052 3528 478104 3534
rect 478052 3470 478104 3476
rect 478064 3398 478092 3470
rect 478052 3392 478104 3398
rect 478052 3334 478104 3340
rect 478156 480 478184 16546
rect 479340 5160 479392 5166
rect 479340 5102 479392 5108
rect 479352 480 479380 5102
rect 480548 480 480576 16546
rect 481652 7546 481680 31486
rect 490012 31476 490064 31482
rect 490012 31418 490064 31424
rect 481732 21616 481784 21622
rect 481732 21558 481784 21564
rect 481640 7540 481692 7546
rect 481640 7482 481692 7488
rect 481744 480 481772 21558
rect 484400 21548 484452 21554
rect 484400 21490 484452 21496
rect 484412 16574 484440 21490
rect 488540 21480 488592 21486
rect 488540 21422 488592 21428
rect 488552 16574 488580 21422
rect 484412 16546 484808 16574
rect 488552 16546 488856 16574
rect 482468 7540 482520 7546
rect 482468 7482 482520 7488
rect 476918 354 477030 480
rect 476500 326 477030 354
rect 476918 -960 477030 326
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482480 354 482508 7482
rect 484032 3596 484084 3602
rect 484032 3538 484084 3544
rect 484044 480 484072 3538
rect 482806 354 482918 480
rect 482480 326 482918 354
rect 482806 -960 482918 326
rect 484002 -960 484114 480
rect 484780 354 484808 16546
rect 486424 11756 486476 11762
rect 486424 11698 486476 11704
rect 486436 480 486464 11698
rect 487620 3392 487672 3398
rect 487620 3334 487672 3340
rect 487632 480 487660 3334
rect 488828 480 488856 16546
rect 490024 6914 490052 31418
rect 496820 31408 496872 31414
rect 496820 31350 496872 31356
rect 492678 30968 492734 30977
rect 492678 30903 492734 30912
rect 491300 21412 491352 21418
rect 491300 21354 491352 21360
rect 491312 16574 491340 21354
rect 492692 16574 492720 30903
rect 495440 23384 495492 23390
rect 495440 23326 495492 23332
rect 491312 16546 492352 16574
rect 492692 16546 493088 16574
rect 489932 6886 490052 6914
rect 489932 480 489960 6886
rect 491116 3460 491168 3466
rect 491116 3402 491168 3408
rect 491128 480 491156 3402
rect 492324 480 492352 16546
rect 485198 354 485310 480
rect 484780 326 485310 354
rect 485198 -960 485310 326
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493060 354 493088 16546
rect 494702 4040 494758 4049
rect 494702 3975 494758 3984
rect 494716 480 494744 3975
rect 493478 354 493590 480
rect 493060 326 493590 354
rect 493478 -960 493590 326
rect 494674 -960 494786 480
rect 495452 354 495480 23326
rect 496832 16574 496860 31350
rect 496832 16546 497136 16574
rect 497108 480 497136 16546
rect 498212 480 498240 72383
rect 503720 31340 503772 31346
rect 503720 31282 503772 31288
rect 498292 23316 498344 23322
rect 498292 23258 498344 23264
rect 498304 16574 498332 23258
rect 502340 23248 502392 23254
rect 502340 23190 502392 23196
rect 502352 16574 502380 23190
rect 498304 16546 498976 16574
rect 502352 16546 503024 16574
rect 495870 354 495982 480
rect 495452 326 495982 354
rect 495870 -960 495982 326
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 498948 354 498976 16546
rect 500592 5092 500644 5098
rect 500592 5034 500644 5040
rect 500604 480 500632 5034
rect 501788 5024 501840 5030
rect 501788 4966 501840 4972
rect 501800 480 501828 4966
rect 502996 480 503024 16546
rect 499366 354 499478 480
rect 498948 326 499478 354
rect 499366 -960 499478 326
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 503732 354 503760 31282
rect 510620 31272 510672 31278
rect 510620 31214 510672 31220
rect 506480 23180 506532 23186
rect 506480 23122 506532 23128
rect 505374 3904 505430 3913
rect 505374 3839 505430 3848
rect 505388 480 505416 3839
rect 506492 480 506520 23122
rect 509238 22672 509294 22681
rect 509238 22607 509294 22616
rect 509252 16574 509280 22607
rect 510632 16574 510660 31214
rect 517520 31204 517572 31210
rect 517520 31146 517572 31152
rect 513380 23112 513432 23118
rect 513380 23054 513432 23060
rect 509252 16546 509648 16574
rect 510632 16546 511304 16574
rect 507214 13016 507270 13025
rect 507214 12951 507270 12960
rect 504150 354 504262 480
rect 503732 326 504262 354
rect 504150 -960 504262 326
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507228 354 507256 12951
rect 508870 5400 508926 5409
rect 508870 5335 508926 5344
rect 508884 480 508912 5335
rect 507646 354 507758 480
rect 507228 326 507758 354
rect 507646 -960 507758 326
rect 508842 -960 508954 480
rect 509620 354 509648 16546
rect 511276 480 511304 16546
rect 512458 5264 512514 5273
rect 512458 5199 512514 5208
rect 512472 480 512500 5199
rect 510038 354 510150 480
rect 509620 326 510150 354
rect 510038 -960 510150 326
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513392 354 513420 23054
rect 516140 23044 516192 23050
rect 516140 22986 516192 22992
rect 516152 16574 516180 22986
rect 517532 16574 517560 31146
rect 520280 22976 520332 22982
rect 520280 22918 520332 22924
rect 516152 16546 517192 16574
rect 517532 16546 517928 16574
rect 514760 6316 514812 6322
rect 514760 6258 514812 6264
rect 514772 480 514800 6258
rect 515954 3768 516010 3777
rect 515954 3703 516010 3712
rect 515968 480 515996 3703
rect 517164 480 517192 16546
rect 513534 354 513646 480
rect 513392 326 513646 354
rect 513534 -960 513646 326
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 517900 354 517928 16546
rect 519544 4956 519596 4962
rect 519544 4898 519596 4904
rect 519556 480 519584 4898
rect 518318 354 518430 480
rect 517900 326 518430 354
rect 518318 -960 518430 326
rect 519514 -960 519626 480
rect 520292 354 520320 22918
rect 520936 3466 520964 72490
rect 549260 32496 549312 32502
rect 549260 32438 549312 32444
rect 524420 31136 524472 31142
rect 524420 31078 524472 31084
rect 521660 31068 521712 31074
rect 521660 31010 521712 31016
rect 520924 3460 520976 3466
rect 520924 3402 520976 3408
rect 520710 354 520822 480
rect 520292 326 520822 354
rect 521672 354 521700 31010
rect 523040 22908 523092 22914
rect 523040 22850 523092 22856
rect 523052 16574 523080 22850
rect 524432 16574 524460 31078
rect 531320 24608 531372 24614
rect 531320 24550 531372 24556
rect 527178 24304 527234 24313
rect 527178 24239 527234 24248
rect 527192 16574 527220 24239
rect 528558 18592 528614 18601
rect 528558 18527 528614 18536
rect 523052 16546 523816 16574
rect 524432 16546 525472 16574
rect 527192 16546 527864 16574
rect 523040 4888 523092 4894
rect 523040 4830 523092 4836
rect 523052 480 523080 4830
rect 521814 354 521926 480
rect 521672 326 521926 354
rect 520710 -960 520822 326
rect 521814 -960 521926 326
rect 523010 -960 523122 480
rect 523788 354 523816 16546
rect 525444 480 525472 16546
rect 526626 6352 526682 6361
rect 526626 6287 526682 6296
rect 526640 480 526668 6287
rect 527836 480 527864 16546
rect 524206 354 524318 480
rect 523788 326 524318 354
rect 524206 -960 524318 326
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528572 354 528600 18527
rect 530122 6216 530178 6225
rect 530122 6151 530178 6160
rect 530136 480 530164 6151
rect 531332 480 531360 24550
rect 534080 24540 534132 24546
rect 534080 24482 534132 24488
rect 534092 16574 534120 24482
rect 538220 24472 538272 24478
rect 538220 24414 538272 24420
rect 535460 18692 535512 18698
rect 535460 18634 535512 18640
rect 535472 16574 535500 18634
rect 534092 16546 534488 16574
rect 535472 16546 536144 16574
rect 532056 15904 532108 15910
rect 532056 15846 532108 15852
rect 528990 354 529102 480
rect 528572 326 529102 354
rect 528990 -960 529102 326
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532068 354 532096 15846
rect 533710 3632 533766 3641
rect 533710 3567 533766 3576
rect 533724 480 533752 3567
rect 532486 354 532598 480
rect 532068 326 532598 354
rect 532486 -960 532598 326
rect 533682 -960 533794 480
rect 534460 354 534488 16546
rect 536116 480 536144 16546
rect 537206 3496 537262 3505
rect 537206 3431 537262 3440
rect 537220 480 537248 3431
rect 534878 354 534990 480
rect 534460 326 534990 354
rect 534878 -960 534990 326
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538232 354 538260 24414
rect 540980 24404 541032 24410
rect 540980 24346 541032 24352
rect 540992 16574 541020 24346
rect 547880 24336 547932 24342
rect 547880 24278 547932 24284
rect 545118 24168 545174 24177
rect 545118 24103 545174 24112
rect 545132 16574 545160 24103
rect 547892 16574 547920 24278
rect 549272 16574 549300 32438
rect 550652 16574 550680 73782
rect 556160 25764 556212 25770
rect 556160 25706 556212 25712
rect 552020 24268 552072 24274
rect 552020 24210 552072 24216
rect 552032 16574 552060 24210
rect 553400 18624 553452 18630
rect 553400 18566 553452 18572
rect 553412 16574 553440 18566
rect 540992 16546 542032 16574
rect 545132 16546 545528 16574
rect 547892 16546 548656 16574
rect 549272 16546 550312 16574
rect 550652 16546 551048 16574
rect 552032 16546 552704 16574
rect 553412 16546 553808 16574
rect 540796 6248 540848 6254
rect 540796 6190 540848 6196
rect 539600 3324 539652 3330
rect 539600 3266 539652 3272
rect 539612 480 539640 3266
rect 540808 480 540836 6190
rect 542004 480 542032 16546
rect 544384 6180 544436 6186
rect 544384 6122 544436 6128
rect 543188 4140 543240 4146
rect 543188 4082 543240 4088
rect 543200 480 543228 4082
rect 544396 480 544424 6122
rect 545500 480 545528 16546
rect 547878 5128 547934 5137
rect 547878 5063 547934 5072
rect 546684 3800 546736 3806
rect 546684 3742 546736 3748
rect 546696 480 546724 3742
rect 547892 480 547920 5063
rect 538374 354 538486 480
rect 538232 326 538486 354
rect 538374 -960 538486 326
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 548628 354 548656 16546
rect 550284 480 550312 16546
rect 549046 354 549158 480
rect 548628 326 549158 354
rect 549046 -960 549158 326
rect 550242 -960 550354 480
rect 551020 354 551048 16546
rect 552676 480 552704 16546
rect 553780 480 553808 16546
rect 554964 7744 555016 7750
rect 554964 7686 555016 7692
rect 554976 480 555004 7686
rect 556172 480 556200 25706
rect 558920 25696 558972 25702
rect 558920 25638 558972 25644
rect 556252 17264 556304 17270
rect 556252 17206 556304 17212
rect 556264 16574 556292 17206
rect 558932 16574 558960 25638
rect 560300 22840 560352 22846
rect 560300 22782 560352 22788
rect 560312 16574 560340 22782
rect 556264 16546 556936 16574
rect 558932 16546 559328 16574
rect 560312 16546 560432 16574
rect 551438 354 551550 480
rect 551020 326 551550 354
rect 551438 -960 551550 326
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 556908 354 556936 16546
rect 558552 7676 558604 7682
rect 558552 7618 558604 7624
rect 558564 480 558592 7618
rect 557326 354 557438 480
rect 556908 326 557438 354
rect 557326 -960 557438 326
rect 558522 -960 558634 480
rect 559300 354 559328 16546
rect 559718 354 559830 480
rect 559300 326 559830 354
rect 560404 354 560432 16546
rect 562046 7712 562102 7721
rect 562046 7647 562102 7656
rect 562060 480 562088 7647
rect 562336 6866 562364 75890
rect 579618 75304 579674 75313
rect 579618 75239 579674 75248
rect 579632 74594 579660 75239
rect 579620 74588 579672 74594
rect 579620 74530 579672 74536
rect 579908 74225 579936 192471
rect 579986 179208 580042 179217
rect 579986 179143 580042 179152
rect 580000 178090 580028 179143
rect 579988 178084 580040 178090
rect 579988 178026 580040 178032
rect 579894 74216 579950 74225
rect 579894 74151 579950 74160
rect 580092 73681 580120 232319
rect 580184 193866 580212 537775
rect 580172 193860 580224 193866
rect 580172 193802 580224 193808
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 580184 99414 580212 99447
rect 580172 99408 580224 99414
rect 580172 99350 580224 99356
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 580184 85610 580212 86119
rect 580172 85604 580224 85610
rect 580172 85546 580224 85552
rect 580276 74769 580304 643991
rect 580354 591016 580410 591025
rect 580354 590951 580410 590960
rect 580262 74760 580318 74769
rect 580262 74695 580318 74704
rect 580078 73672 580134 73681
rect 580078 73607 580134 73616
rect 580368 73137 580396 590951
rect 580460 174350 580488 683839
rect 580538 630864 580594 630873
rect 580538 630799 580594 630808
rect 580448 174344 580500 174350
rect 580448 174286 580500 174292
rect 580446 152688 580502 152697
rect 580446 152623 580502 152632
rect 580460 73817 580488 152623
rect 580552 149734 580580 630799
rect 580630 577688 580686 577697
rect 580630 577623 580686 577632
rect 580540 149728 580592 149734
rect 580540 149670 580592 149676
rect 580644 144226 580672 577623
rect 580814 524512 580870 524521
rect 580814 524447 580870 524456
rect 580722 484664 580778 484673
rect 580722 484599 580778 484608
rect 580632 144220 580684 144226
rect 580632 144162 580684 144168
rect 580538 112840 580594 112849
rect 580538 112775 580594 112784
rect 580552 74526 580580 112775
rect 580540 74520 580592 74526
rect 580540 74462 580592 74468
rect 580446 73808 580502 73817
rect 580446 73743 580502 73752
rect 580354 73128 580410 73137
rect 580736 73098 580764 484599
rect 580828 135930 580856 524447
rect 580906 431624 580962 431633
rect 580906 431559 580962 431568
rect 580816 135924 580868 135930
rect 580816 135866 580868 135872
rect 580920 74633 580948 431559
rect 580906 74624 580962 74633
rect 580906 74559 580962 74568
rect 580354 73063 580410 73072
rect 580724 73092 580776 73098
rect 580724 73034 580776 73040
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 580184 72010 580212 72927
rect 580264 72480 580316 72486
rect 580264 72422 580316 72428
rect 580172 72004 580224 72010
rect 580172 71946 580224 71952
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 580276 33153 580304 72422
rect 581092 71052 581144 71058
rect 581092 70994 581144 71000
rect 580262 33144 580318 33153
rect 580262 33079 580318 33088
rect 574100 32428 574152 32434
rect 574100 32370 574152 32376
rect 571340 28280 571392 28286
rect 571340 28222 571392 28228
rect 565820 25628 565872 25634
rect 565820 25570 565872 25576
rect 565832 16574 565860 25570
rect 567200 24200 567252 24206
rect 567200 24142 567252 24148
rect 567212 16574 567240 24142
rect 569960 24132 570012 24138
rect 569960 24074 570012 24080
rect 569972 16574 570000 24074
rect 565832 16546 566872 16574
rect 567212 16546 567608 16574
rect 569972 16546 570368 16574
rect 564438 7576 564494 7585
rect 564438 7511 564494 7520
rect 562324 6860 562376 6866
rect 562324 6802 562376 6808
rect 563242 4992 563298 5001
rect 563242 4927 563298 4936
rect 563256 480 563284 4927
rect 564452 480 564480 7511
rect 565634 4856 565690 4865
rect 565634 4791 565690 4800
rect 565648 480 565676 4791
rect 566844 480 566872 16546
rect 560822 354 560934 480
rect 560404 326 560934 354
rect 559718 -960 559830 326
rect 560822 -960 560934 326
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567580 354 567608 16546
rect 569132 7608 569184 7614
rect 569132 7550 569184 7556
rect 569144 480 569172 7550
rect 570340 480 570368 16546
rect 567998 354 568110 480
rect 567580 326 568110 354
rect 567998 -960 568110 326
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571352 354 571380 28222
rect 572720 25560 572772 25566
rect 572720 25502 572772 25508
rect 572732 16574 572760 25502
rect 574112 16574 574140 32370
rect 580172 22772 580224 22778
rect 580172 22714 580224 22720
rect 580184 19825 580212 22714
rect 580170 19816 580226 19825
rect 580170 19751 580226 19760
rect 572732 16546 573496 16574
rect 574112 16546 575152 16574
rect 572720 8968 572772 8974
rect 572720 8910 572772 8916
rect 572732 480 572760 8910
rect 571494 354 571606 480
rect 571352 326 571606 354
rect 571494 -960 571606 326
rect 572690 -960 572802 480
rect 573468 354 573496 16546
rect 575124 480 575152 16546
rect 576306 9072 576362 9081
rect 576306 9007 576362 9016
rect 576320 480 576348 9007
rect 578606 8936 578662 8945
rect 578606 8871 578662 8880
rect 577412 4820 577464 4826
rect 577412 4762 577464 4768
rect 577424 480 577452 4762
rect 578620 480 578648 8871
rect 581104 6914 581132 70994
rect 581012 6886 581132 6914
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 581012 480 581040 6886
rect 582196 3460 582248 3466
rect 582196 3402 582248 3408
rect 582208 480 582236 3402
rect 583390 3360 583446 3369
rect 583390 3295 583446 3304
rect 583404 480 583432 3295
rect 573886 354 573998 480
rect 573468 326 573998 354
rect 573886 -960 573998 326
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3330 566888 3386 566944
rect 2778 553852 2834 553888
rect 2778 553832 2780 553852
rect 2780 553832 2832 553852
rect 2832 553832 2834 553852
rect 3330 514820 3386 514856
rect 3330 514800 3332 514820
rect 3332 514800 3384 514820
rect 3384 514800 3386 514820
rect 2778 501744 2834 501800
rect 2778 462596 2834 462632
rect 2778 462576 2780 462596
rect 2780 462576 2832 462596
rect 2832 462576 2834 462596
rect 2778 449520 2834 449576
rect 3330 410488 3386 410544
rect 2778 397468 2780 397488
rect 2780 397468 2832 397488
rect 2832 397468 2834 397488
rect 2778 397432 2834 397468
rect 3330 358400 3386 358456
rect 2778 345344 2834 345400
rect 3330 319232 3386 319288
rect 3238 306176 3294 306232
rect 3238 293120 3294 293176
rect 3238 267144 3294 267200
rect 3146 254088 3202 254144
rect 3054 241032 3110 241088
rect 3146 214920 3202 214976
rect 3146 201864 3202 201920
rect 3146 188808 3202 188864
rect 3146 162868 3148 162888
rect 3148 162868 3200 162888
rect 3200 162868 3202 162888
rect 3146 162832 3202 162868
rect 3146 149776 3202 149832
rect 3514 671200 3570 671256
rect 3606 632032 3662 632088
rect 3514 619112 3570 619168
rect 3514 606056 3570 606112
rect 3422 136720 3478 136776
rect 3330 84632 3386 84688
rect 2870 32408 2926 32464
rect 3698 579944 3754 580000
rect 3790 527856 3846 527912
rect 3882 475632 3938 475688
rect 4066 423544 4122 423600
rect 3974 371320 4030 371376
rect 3514 74296 3570 74352
rect 3514 71576 3570 71632
rect 3790 110608 3846 110664
rect 3698 97552 3754 97608
rect 4802 74976 4858 75032
rect 4986 75112 5042 75168
rect 4894 73888 4950 73944
rect 395526 240080 395582 240136
rect 395342 239944 395398 240000
rect 394606 232056 394662 232112
rect 6918 74024 6974 74080
rect 114006 137264 114062 137320
rect 113730 131164 113786 131200
rect 113730 131144 113732 131164
rect 113732 131144 113784 131164
rect 113784 131144 113786 131164
rect 113730 128968 113786 129024
rect 113638 127472 113694 127528
rect 113730 126792 113786 126848
rect 113546 125296 113602 125352
rect 113730 123800 113786 123856
rect 113362 122748 113364 122768
rect 113364 122748 113416 122768
rect 113416 122748 113418 122768
rect 113362 122712 113418 122748
rect 113730 121216 113786 121272
rect 113730 119720 113786 119776
rect 113638 118224 113694 118280
rect 113730 116728 113786 116784
rect 113730 115232 113786 115288
rect 113730 113092 113732 113112
rect 113732 113092 113784 113112
rect 113784 113092 113786 113112
rect 113730 113056 113786 113092
rect 113730 111732 113732 111752
rect 113732 111732 113784 111752
rect 113784 111732 113786 111752
rect 113730 111696 113786 111732
rect 113730 110372 113732 110392
rect 113732 110372 113784 110392
rect 113784 110372 113786 110392
rect 113730 110336 113786 110372
rect 113730 108840 113786 108896
rect 113546 107344 113602 107400
rect 113730 106120 113786 106176
rect 113362 104796 113364 104816
rect 113364 104796 113416 104816
rect 113416 104796 113418 104816
rect 113362 104760 113418 104796
rect 113822 101768 113878 101824
rect 113914 98776 113970 98832
rect 114006 91024 114062 91080
rect 114098 89664 114154 89720
rect 114190 88168 114246 88224
rect 114282 86808 114338 86864
rect 114374 85312 114430 85368
rect 115110 133184 115166 133240
rect 114466 80824 114522 80880
rect 114374 76608 114430 76664
rect 22742 72528 22798 72584
rect 3606 58520 3662 58576
rect 3514 45500 3516 45520
rect 3516 45500 3568 45520
rect 3568 45500 3570 45520
rect 3514 45464 3570 45500
rect 3422 19352 3478 19408
rect 3514 6432 3570 6488
rect 1674 3440 1730 3496
rect 570 3304 626 3360
rect 18234 6160 18290 6216
rect 17038 3576 17094 3632
rect 34794 8880 34850 8936
rect 38382 9016 38438 9072
rect 37186 4800 37242 4856
rect 53746 9152 53802 9208
rect 52550 6296 52606 6352
rect 56046 6432 56102 6488
rect 54942 3712 54998 3768
rect 71502 10240 71558 10296
rect 70306 7520 70362 7576
rect 114466 75384 114522 75440
rect 115294 103128 115350 103184
rect 115662 96668 115718 96724
rect 115570 95104 115626 95160
rect 115478 93744 115534 93800
rect 115386 92384 115442 92440
rect 390374 231104 390430 231160
rect 138110 195880 138166 195936
rect 140410 195880 140466 195936
rect 141422 195916 141424 195936
rect 141424 195916 141476 195936
rect 141476 195916 141478 195936
rect 141422 195880 141478 195916
rect 158902 195872 158958 195928
rect 160834 195880 160890 195936
rect 157154 195608 157210 195664
rect 139398 195472 139454 195528
rect 140870 191800 140926 191856
rect 140778 191664 140834 191720
rect 140778 184184 140834 184240
rect 115938 100272 115994 100328
rect 115846 83204 115902 83260
rect 115754 81708 115810 81764
rect 116490 78376 116546 78432
rect 116490 75520 116546 75576
rect 140962 190848 141018 190904
rect 140962 184320 141018 184376
rect 140870 184048 140926 184104
rect 144366 190984 144422 191040
rect 145838 189760 145894 189816
rect 144826 189216 144882 189272
rect 157338 188944 157394 189000
rect 144918 182008 144974 182064
rect 141238 181056 141294 181112
rect 144642 180920 144698 180976
rect 142666 179016 142722 179072
rect 144090 178880 144146 178936
rect 141698 178744 141754 178800
rect 141790 178608 141846 178664
rect 157798 178064 157854 178120
rect 158534 178064 158590 178120
rect 139674 137944 139730 138000
rect 147494 174528 147550 174584
rect 161570 137672 161626 137728
rect 167826 137536 167882 137592
rect 169390 137400 169446 137456
rect 175370 129920 175426 129976
rect 175370 128288 175426 128344
rect 175554 132368 175610 132424
rect 175462 111832 175518 111888
rect 89166 10376 89222 10432
rect 87970 7656 88026 7712
rect 91558 7792 91614 7848
rect 90362 4936 90418 4992
rect 105726 9288 105782 9344
rect 109314 9424 109370 9480
rect 108118 6568 108174 6624
rect 121642 71984 121698 72040
rect 121550 71848 121606 71904
rect 121918 72528 121974 72584
rect 122838 71984 122894 72040
rect 122930 71848 122986 71904
rect 124218 72120 124274 72176
rect 124402 71984 124458 72040
rect 124494 71848 124550 71904
rect 125690 72256 125746 72312
rect 125782 72120 125838 72176
rect 125598 71984 125654 72040
rect 125874 71848 125930 71904
rect 127070 71984 127126 72040
rect 126978 71848 127034 71904
rect 128542 73072 128598 73128
rect 128450 72120 128506 72176
rect 128358 71984 128414 72040
rect 128634 71848 128690 71904
rect 129738 72120 129794 72176
rect 130014 71984 130070 72040
rect 129922 71848 129978 71904
rect 123482 3576 123538 3632
rect 124678 3440 124734 3496
rect 131210 71984 131266 72040
rect 131118 71848 131174 71904
rect 132222 71984 132278 72040
rect 132406 71848 132462 71904
rect 133602 72120 133658 72176
rect 133694 71984 133750 72040
rect 133786 71848 133842 71904
rect 135074 72120 135130 72176
rect 134982 71984 135038 72040
rect 135166 71848 135222 71904
rect 136454 72120 136510 72176
rect 136362 71984 136418 72040
rect 136178 71848 136234 71904
rect 136546 71848 136602 71904
rect 137834 71984 137890 72040
rect 137926 71848 137982 71904
rect 137650 3576 137706 3632
rect 139030 71984 139086 72040
rect 139306 72120 139362 72176
rect 138938 71848 138994 71904
rect 139122 71848 139178 71904
rect 140318 72120 140374 72176
rect 140594 71984 140650 72040
rect 140410 71848 140466 71904
rect 140686 71848 140742 71904
rect 141974 71984 142030 72040
rect 142066 71848 142122 71904
rect 143262 72256 143318 72312
rect 143354 72120 143410 72176
rect 143446 71984 143502 72040
rect 143170 71848 143226 71904
rect 144734 72120 144790 72176
rect 144642 71984 144698 72040
rect 144550 71848 144606 71904
rect 144826 71848 144882 71904
rect 146022 72120 146078 72176
rect 146206 71984 146262 72040
rect 146114 71848 146170 71904
rect 147494 72120 147550 72176
rect 147402 71984 147458 72040
rect 147310 71848 147366 71904
rect 147586 71848 147642 71904
rect 148690 72664 148746 72720
rect 148966 72800 149022 72856
rect 148874 72528 148930 72584
rect 148782 72392 148838 72448
rect 140042 3440 140098 3496
rect 149978 72664 150034 72720
rect 150162 72936 150218 72992
rect 150346 72800 150402 72856
rect 150070 72528 150126 72584
rect 151542 72664 151598 72720
rect 151726 72800 151782 72856
rect 151634 72392 151690 72448
rect 152002 74568 152058 74624
rect 152922 72800 152978 72856
rect 153014 72664 153070 72720
rect 152830 72392 152886 72448
rect 153106 72528 153162 72584
rect 154118 72800 154174 72856
rect 154302 72936 154358 72992
rect 154210 72664 154266 72720
rect 154486 72528 154542 72584
rect 155774 72800 155830 72856
rect 155866 72664 155922 72720
rect 155682 72392 155738 72448
rect 156970 72800 157026 72856
rect 156878 72664 156934 72720
rect 157062 72528 157118 72584
rect 157062 72392 157118 72448
rect 157246 72664 157302 72720
rect 157154 72120 157210 72176
rect 157522 74604 157524 74624
rect 157524 74604 157576 74624
rect 157576 74604 157578 74624
rect 157522 74568 157578 74604
rect 157798 72120 157854 72176
rect 158350 72664 158406 72720
rect 158442 72528 158498 72584
rect 158626 72800 158682 72856
rect 158534 72392 158590 72448
rect 158902 71984 158958 72040
rect 158810 71848 158866 71904
rect 155406 4936 155462 4992
rect 156602 4800 156658 4856
rect 157798 3304 157854 3360
rect 159638 72256 159694 72312
rect 159914 72800 159970 72856
rect 160006 72664 160062 72720
rect 160282 72120 160338 72176
rect 161018 72664 161074 72720
rect 161294 73072 161350 73128
rect 161202 72800 161258 72856
rect 161386 72528 161442 72584
rect 161110 72392 161166 72448
rect 161018 72256 161074 72312
rect 161662 74296 161718 74352
rect 162398 74840 162454 74896
rect 162398 74296 162454 74352
rect 162398 73208 162454 73264
rect 162398 73072 162454 73128
rect 162582 72936 162638 72992
rect 162490 72664 162546 72720
rect 162766 72800 162822 72856
rect 162674 72528 162730 72584
rect 162766 72392 162822 72448
rect 163042 73072 163098 73128
rect 163318 72936 163374 72992
rect 164054 72800 164110 72856
rect 163962 72664 164018 72720
rect 164146 72392 164202 72448
rect 165250 72664 165306 72720
rect 165526 72800 165582 72856
rect 165434 72528 165490 72584
rect 160834 3848 160890 3904
rect 165342 72392 165398 72448
rect 166446 72664 166502 72720
rect 166354 72528 166410 72584
rect 166814 72664 166870 72720
rect 166814 72528 166870 72584
rect 166538 72392 166594 72448
rect 167182 74432 167238 74488
rect 167274 74160 167330 74216
rect 166814 71984 166870 72040
rect 166906 31728 166962 31784
rect 167458 74840 167514 74896
rect 167734 74840 167790 74896
rect 167642 74704 167698 74760
rect 167366 73616 167422 73672
rect 168102 74568 168158 74624
rect 168194 74432 168250 74488
rect 168194 73752 168250 73808
rect 168010 73072 168066 73128
rect 169114 74296 169170 74352
rect 169298 74704 169354 74760
rect 169206 74024 169262 74080
rect 169022 73888 169078 73944
rect 169482 74840 169538 74896
rect 169390 73480 169446 73536
rect 169666 74840 169722 74896
rect 171414 75420 171416 75440
rect 171416 75420 171468 75440
rect 171468 75420 171470 75440
rect 170402 74840 170458 74896
rect 171414 75384 171470 75420
rect 171690 75248 171746 75304
rect 171690 74568 171746 74624
rect 175646 126928 175702 126984
rect 177854 121216 177910 121272
rect 178038 118224 178094 118280
rect 178130 113056 178186 113112
rect 178038 110336 178094 110392
rect 178590 131144 178646 131200
rect 178498 124072 178554 124128
rect 178406 119720 178462 119776
rect 178314 115232 178370 115288
rect 178222 108976 178278 109032
rect 176750 107480 176806 107536
rect 178038 105984 178094 106040
rect 178038 104488 178094 104544
rect 178038 102992 178094 103048
rect 178038 101632 178094 101688
rect 178038 100136 178094 100192
rect 178038 98776 178094 98832
rect 178038 97280 178094 97336
rect 178038 95140 178040 95160
rect 178040 95140 178092 95160
rect 178092 95140 178094 95160
rect 178038 95104 178094 95140
rect 178038 93780 178040 93800
rect 178040 93780 178092 93800
rect 178092 93780 178094 93800
rect 178038 93744 178094 93780
rect 178038 92248 178094 92304
rect 178038 90888 178094 90944
rect 178038 89392 178094 89448
rect 178038 88032 178094 88088
rect 178038 86536 178094 86592
rect 178038 85040 178094 85096
rect 178038 83680 178094 83736
rect 178038 82184 178094 82240
rect 178038 76608 178094 76664
rect 175922 75520 175978 75576
rect 178866 125432 178922 125488
rect 178774 122440 178830 122496
rect 178682 116728 178738 116784
rect 178682 80824 178738 80880
rect 178682 78648 178738 78704
rect 173898 32680 173954 32736
rect 172518 25608 172574 25664
rect 169666 8064 169722 8120
rect 187698 32544 187754 32600
rect 191838 32408 191894 32464
rect 190458 27104 190514 27160
rect 193310 4664 193366 4720
rect 209778 34040 209834 34096
rect 210974 12144 211030 12200
rect 223578 20168 223634 20224
rect 225142 12824 225198 12880
rect 226430 6840 226486 6896
rect 228730 6704 228786 6760
rect 241518 33904 241574 33960
rect 244278 20032 244334 20088
rect 242990 13640 243046 13696
rect 246394 6568 246450 6624
rect 262218 33768 262274 33824
rect 264150 15136 264206 15192
rect 278778 26968 278834 27024
rect 278318 7928 278374 7984
rect 280710 13504 280766 13560
rect 281906 7792 281962 7848
rect 298098 35264 298154 35320
rect 295614 16224 295670 16280
rect 297270 15000 297326 15056
rect 299662 9152 299718 9208
rect 314658 29552 314714 29608
rect 316038 17584 316094 17640
rect 316222 14864 316278 14920
rect 332598 35128 332654 35184
rect 331218 10376 331274 10432
rect 396722 74840 396778 74896
rect 350538 21528 350594 21584
rect 332690 14728 332746 14784
rect 334622 10240 334678 10296
rect 349158 16088 349214 16144
rect 349250 12008 349306 12064
rect 352838 11872 352894 11928
rect 367098 26832 367154 26888
rect 365718 13368 365774 13424
rect 365810 11736 365866 11792
rect 370134 13232 370190 13288
rect 386418 24384 386474 24440
rect 385958 6432 386014 6488
rect 387798 14592 387854 14648
rect 405002 72664 405058 72720
rect 402518 14456 402574 14512
rect 403622 11600 403678 11656
rect 404818 5480 404874 5536
rect 406014 15952 406070 16008
rect 420918 17448 420974 17504
rect 420182 15816 420238 15872
rect 418526 13096 418582 13152
rect 445022 31184 445078 31240
rect 423770 17312 423826 17368
rect 440238 21392 440294 21448
rect 440330 17176 440386 17232
rect 454038 22752 454094 22808
rect 455418 18808 455474 18864
rect 456890 25472 456946 25528
rect 458178 18672 458234 18728
rect 580446 683848 580502 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580262 644000 580318 644056
rect 579986 617480 580042 617536
rect 580170 564304 580226 564360
rect 580170 537784 580226 537840
rect 579802 511264 579858 511320
rect 579986 458088 580042 458144
rect 580078 444760 580134 444816
rect 580078 418240 580134 418296
rect 580078 404912 580134 404968
rect 580078 378392 580134 378448
rect 579802 365064 579858 365120
rect 580078 351908 580080 351928
rect 580080 351908 580132 351928
rect 580132 351908 580134 351928
rect 580078 351872 580134 351908
rect 580078 325216 580134 325272
rect 580078 312024 580134 312080
rect 580078 298696 580134 298752
rect 579802 272176 579858 272232
rect 579986 258848 580042 258904
rect 579986 245520 580042 245576
rect 580078 232328 580134 232384
rect 579802 219000 579858 219056
rect 579986 205692 580042 205728
rect 579986 205672 579988 205692
rect 579988 205672 580040 205692
rect 580040 205672 580042 205692
rect 579894 192480 579950 192536
rect 579802 165824 579858 165880
rect 579618 139304 579674 139360
rect 579710 125976 579766 126032
rect 480258 72528 480314 72584
rect 474738 65456 474794 65512
rect 473358 31048 473414 31104
rect 473450 19896 473506 19952
rect 476118 21256 476174 21312
rect 498198 72392 498254 72448
rect 492678 30912 492734 30968
rect 494702 3984 494758 4040
rect 505374 3848 505430 3904
rect 509238 22616 509294 22672
rect 507214 12960 507270 13016
rect 508870 5344 508926 5400
rect 512458 5208 512514 5264
rect 515954 3712 516010 3768
rect 527178 24248 527234 24304
rect 528558 18536 528614 18592
rect 526626 6296 526682 6352
rect 530122 6160 530178 6216
rect 533710 3576 533766 3632
rect 537206 3440 537262 3496
rect 545118 24112 545174 24168
rect 547878 5072 547934 5128
rect 562046 7656 562102 7712
rect 579618 75248 579674 75304
rect 579986 179152 580042 179208
rect 579894 74160 579950 74216
rect 580170 99456 580226 99512
rect 580170 86128 580226 86184
rect 580354 590960 580410 591016
rect 580262 74704 580318 74760
rect 580078 73616 580134 73672
rect 580538 630808 580594 630864
rect 580446 152632 580502 152688
rect 580630 577632 580686 577688
rect 580814 524456 580870 524512
rect 580722 484608 580778 484664
rect 580538 112784 580594 112840
rect 580446 73752 580502 73808
rect 580354 73072 580410 73128
rect 580906 431568 580962 431624
rect 580906 74568 580962 74624
rect 580170 72936 580226 72992
rect 580170 59608 580226 59664
rect 580170 46280 580226 46336
rect 580262 33088 580318 33144
rect 564438 7520 564494 7576
rect 563242 4936 563298 4992
rect 565634 4800 565690 4856
rect 580170 19760 580226 19816
rect 576306 9016 576362 9072
rect 578606 8880 578662 8936
rect 580170 6568 580226 6624
rect 583390 3304 583446 3360
<< metal3 >>
rect -960 697220 480 697460
rect 580758 697172 580764 697236
rect 580828 697234 580834 697236
rect 583520 697234 584960 697324
rect 580828 697174 584960 697234
rect 580828 697172 580834 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580441 683906 580507 683909
rect 583520 683906 584960 683996
rect 580441 683904 584960 683906
rect 580441 683848 580446 683904
rect 580502 683848 584960 683904
rect 580441 683846 584960 683848
rect 580441 683843 580507 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3366 658202 3372 658204
rect -960 658142 3372 658202
rect -960 658052 480 658142
rect 3366 658140 3372 658142
rect 3436 658140 3442 658204
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580257 644058 580323 644061
rect 583520 644058 584960 644148
rect 580257 644056 584960 644058
rect 580257 644000 580262 644056
rect 580318 644000 584960 644056
rect 580257 643998 584960 644000
rect 580257 643995 580323 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3601 632090 3667 632093
rect -960 632088 3667 632090
rect -960 632032 3606 632088
rect 3662 632032 3667 632088
rect -960 632030 3667 632032
rect -960 631940 480 632030
rect 3601 632027 3667 632030
rect 580533 630866 580599 630869
rect 583520 630866 584960 630956
rect 580533 630864 584960 630866
rect 580533 630808 580538 630864
rect 580594 630808 584960 630864
rect 580533 630806 584960 630808
rect 580533 630803 580599 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3509 619170 3575 619173
rect -960 619168 3575 619170
rect -960 619112 3514 619168
rect 3570 619112 3575 619168
rect -960 619110 3575 619112
rect -960 619020 480 619110
rect 3509 619107 3575 619110
rect 579981 617538 580047 617541
rect 583520 617538 584960 617628
rect 579981 617536 584960 617538
rect 579981 617480 579986 617536
rect 580042 617480 584960 617536
rect 579981 617478 584960 617480
rect 579981 617475 580047 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3509 606114 3575 606117
rect -960 606112 3575 606114
rect -960 606056 3514 606112
rect 3570 606056 3575 606112
rect -960 606054 3575 606056
rect -960 605964 480 606054
rect 3509 606051 3575 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 580349 591018 580415 591021
rect 583520 591018 584960 591108
rect 580349 591016 584960 591018
rect 580349 590960 580354 591016
rect 580410 590960 584960 591016
rect 580349 590958 584960 590960
rect 580349 590955 580415 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3693 580002 3759 580005
rect -960 580000 3759 580002
rect -960 579944 3698 580000
rect 3754 579944 3759 580000
rect -960 579942 3759 579944
rect -960 579852 480 579942
rect 3693 579939 3759 579942
rect 580625 577690 580691 577693
rect 583520 577690 584960 577780
rect 580625 577688 584960 577690
rect 580625 577632 580630 577688
rect 580686 577632 584960 577688
rect 580625 577630 584960 577632
rect 580625 577627 580691 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3325 566946 3391 566949
rect -960 566944 3391 566946
rect -960 566888 3330 566944
rect 3386 566888 3391 566944
rect -960 566886 3391 566888
rect -960 566796 480 566886
rect 3325 566883 3391 566886
rect 580165 564362 580231 564365
rect 583520 564362 584960 564452
rect 580165 564360 584960 564362
rect 580165 564304 580170 564360
rect 580226 564304 584960 564360
rect 580165 564302 584960 564304
rect 580165 564299 580231 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 2773 553890 2839 553893
rect -960 553888 2839 553890
rect -960 553832 2778 553888
rect 2834 553832 2839 553888
rect -960 553830 2839 553832
rect -960 553740 480 553830
rect 2773 553827 2839 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 3785 527914 3851 527917
rect -960 527912 3851 527914
rect -960 527856 3790 527912
rect 3846 527856 3851 527912
rect -960 527854 3851 527856
rect -960 527764 480 527854
rect 3785 527851 3851 527854
rect 580809 524514 580875 524517
rect 583520 524514 584960 524604
rect 580809 524512 584960 524514
rect 580809 524456 580814 524512
rect 580870 524456 584960 524512
rect 580809 524454 584960 524456
rect 580809 524451 580875 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3325 514858 3391 514861
rect -960 514856 3391 514858
rect -960 514800 3330 514856
rect 3386 514800 3391 514856
rect -960 514798 3391 514800
rect -960 514708 480 514798
rect 3325 514795 3391 514798
rect 579797 511322 579863 511325
rect 583520 511322 584960 511412
rect 579797 511320 584960 511322
rect 579797 511264 579802 511320
rect 579858 511264 584960 511320
rect 579797 511262 584960 511264
rect 579797 511259 579863 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 2773 501802 2839 501805
rect -960 501800 2839 501802
rect -960 501744 2778 501800
rect 2834 501744 2839 501800
rect -960 501742 2839 501744
rect -960 501652 480 501742
rect 2773 501739 2839 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580717 484666 580783 484669
rect 583520 484666 584960 484756
rect 580717 484664 584960 484666
rect 580717 484608 580722 484664
rect 580778 484608 584960 484664
rect 580717 484606 584960 484608
rect 580717 484603 580783 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3877 475690 3943 475693
rect -960 475688 3943 475690
rect -960 475632 3882 475688
rect 3938 475632 3943 475688
rect -960 475630 3943 475632
rect -960 475540 480 475630
rect 3877 475627 3943 475630
rect 583520 471474 584960 471564
rect 583342 471414 584960 471474
rect 583342 471338 583402 471414
rect 583520 471338 584960 471414
rect 583342 471324 584960 471338
rect 583342 471278 583586 471324
rect 396574 470596 396580 470660
rect 396644 470658 396650 470660
rect 583526 470658 583586 471278
rect 396644 470598 583586 470658
rect 396644 470596 396650 470598
rect -960 462634 480 462724
rect 2773 462634 2839 462637
rect -960 462632 2839 462634
rect -960 462576 2778 462632
rect 2834 462576 2839 462632
rect -960 462574 2839 462576
rect -960 462484 480 462574
rect 2773 462571 2839 462574
rect 579981 458146 580047 458149
rect 583520 458146 584960 458236
rect 579981 458144 584960 458146
rect 579981 458088 579986 458144
rect 580042 458088 584960 458144
rect 579981 458086 584960 458088
rect 579981 458083 580047 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 2773 449578 2839 449581
rect -960 449576 2839 449578
rect -960 449520 2778 449576
rect 2834 449520 2839 449576
rect -960 449518 2839 449520
rect -960 449428 480 449518
rect 2773 449515 2839 449518
rect 580073 444818 580139 444821
rect 583520 444818 584960 444908
rect 580073 444816 584960 444818
rect 580073 444760 580078 444816
rect 580134 444760 584960 444816
rect 580073 444758 584960 444760
rect 580073 444755 580139 444758
rect 583520 444668 584960 444758
rect -960 436508 480 436748
rect 580901 431626 580967 431629
rect 583520 431626 584960 431716
rect 580901 431624 584960 431626
rect 580901 431568 580906 431624
rect 580962 431568 584960 431624
rect 580901 431566 584960 431568
rect 580901 431563 580967 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 4061 423602 4127 423605
rect -960 423600 4127 423602
rect -960 423544 4066 423600
rect 4122 423544 4127 423600
rect -960 423542 4127 423544
rect -960 423452 480 423542
rect 4061 423539 4127 423542
rect 580073 418298 580139 418301
rect 583520 418298 584960 418388
rect 580073 418296 584960 418298
rect 580073 418240 580078 418296
rect 580134 418240 584960 418296
rect 580073 418238 584960 418240
rect 580073 418235 580139 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3325 410546 3391 410549
rect -960 410544 3391 410546
rect -960 410488 3330 410544
rect 3386 410488 3391 410544
rect -960 410486 3391 410488
rect -960 410396 480 410486
rect 3325 410483 3391 410486
rect 580073 404970 580139 404973
rect 583520 404970 584960 405060
rect 580073 404968 584960 404970
rect 580073 404912 580078 404968
rect 580134 404912 584960 404968
rect 580073 404910 584960 404912
rect 580073 404907 580139 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 2773 397490 2839 397493
rect -960 397488 2839 397490
rect -960 397432 2778 397488
rect 2834 397432 2839 397488
rect -960 397430 2839 397432
rect -960 397340 480 397430
rect 2773 397427 2839 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580073 378450 580139 378453
rect 583520 378450 584960 378540
rect 580073 378448 584960 378450
rect 580073 378392 580078 378448
rect 580134 378392 584960 378448
rect 580073 378390 584960 378392
rect 580073 378387 580139 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 3969 371378 4035 371381
rect -960 371376 4035 371378
rect -960 371320 3974 371376
rect 4030 371320 4035 371376
rect -960 371318 4035 371320
rect -960 371228 480 371318
rect 3969 371315 4035 371318
rect 579797 365122 579863 365125
rect 583520 365122 584960 365212
rect 579797 365120 584960 365122
rect 579797 365064 579802 365120
rect 579858 365064 584960 365120
rect 579797 365062 584960 365064
rect 579797 365059 579863 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 3325 358458 3391 358461
rect -960 358456 3391 358458
rect -960 358400 3330 358456
rect 3386 358400 3391 358456
rect -960 358398 3391 358400
rect -960 358308 480 358398
rect 3325 358395 3391 358398
rect 580073 351930 580139 351933
rect 583520 351930 584960 352020
rect 580073 351928 584960 351930
rect 580073 351872 580078 351928
rect 580134 351872 584960 351928
rect 580073 351870 584960 351872
rect 580073 351867 580139 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 2773 345402 2839 345405
rect -960 345400 2839 345402
rect -960 345344 2778 345400
rect 2834 345344 2839 345400
rect -960 345342 2839 345344
rect -960 345252 480 345342
rect 2773 345339 2839 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 580073 325274 580139 325277
rect 583520 325274 584960 325364
rect 580073 325272 584960 325274
rect 580073 325216 580078 325272
rect 580134 325216 584960 325272
rect 580073 325214 584960 325216
rect 580073 325211 580139 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3325 319290 3391 319293
rect -960 319288 3391 319290
rect -960 319232 3330 319288
rect 3386 319232 3391 319288
rect -960 319230 3391 319232
rect -960 319140 480 319230
rect 3325 319227 3391 319230
rect 580073 312082 580139 312085
rect 583520 312082 584960 312172
rect 580073 312080 584960 312082
rect 580073 312024 580078 312080
rect 580134 312024 584960 312080
rect 580073 312022 584960 312024
rect 580073 312019 580139 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3233 306234 3299 306237
rect -960 306232 3299 306234
rect -960 306176 3238 306232
rect 3294 306176 3299 306232
rect -960 306174 3299 306176
rect -960 306084 480 306174
rect 3233 306171 3299 306174
rect 580073 298754 580139 298757
rect 583520 298754 584960 298844
rect 580073 298752 584960 298754
rect 580073 298696 580078 298752
rect 580134 298696 584960 298752
rect 580073 298694 584960 298696
rect 580073 298691 580139 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 3233 293178 3299 293181
rect -960 293176 3299 293178
rect -960 293120 3238 293176
rect 3294 293120 3299 293176
rect -960 293118 3299 293120
rect -960 293028 480 293118
rect 3233 293115 3299 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 579797 272234 579863 272237
rect 583520 272234 584960 272324
rect 579797 272232 584960 272234
rect 579797 272176 579802 272232
rect 579858 272176 584960 272232
rect 579797 272174 584960 272176
rect 579797 272171 579863 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 3233 267202 3299 267205
rect -960 267200 3299 267202
rect -960 267144 3238 267200
rect 3294 267144 3299 267200
rect -960 267142 3299 267144
rect -960 267052 480 267142
rect 3233 267139 3299 267142
rect 579981 258906 580047 258909
rect 583520 258906 584960 258996
rect 579981 258904 584960 258906
rect 579981 258848 579986 258904
rect 580042 258848 584960 258904
rect 579981 258846 584960 258848
rect 579981 258843 580047 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 3141 254146 3207 254149
rect -960 254144 3207 254146
rect -960 254088 3146 254144
rect 3202 254088 3207 254144
rect -960 254086 3207 254088
rect -960 253996 480 254086
rect 3141 254083 3207 254086
rect 579981 245578 580047 245581
rect 583520 245578 584960 245668
rect 579981 245576 584960 245578
rect 579981 245520 579986 245576
rect 580042 245520 584960 245576
rect 579981 245518 584960 245520
rect 579981 245515 580047 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 3049 241090 3115 241093
rect -960 241088 3115 241090
rect -960 241032 3054 241088
rect 3110 241032 3115 241088
rect -960 241030 3115 241032
rect -960 240940 480 241030
rect 3049 241027 3115 241030
rect 395521 240138 395587 240141
rect 396758 240138 396764 240140
rect 395521 240136 396764 240138
rect 395521 240080 395526 240136
rect 395582 240080 396764 240136
rect 395521 240078 396764 240080
rect 395521 240075 395587 240078
rect 396758 240076 396764 240078
rect 396828 240076 396834 240140
rect 395337 240002 395403 240005
rect 396942 240002 396948 240004
rect 395337 240000 396948 240002
rect 395337 239944 395342 240000
rect 395398 239944 396948 240000
rect 395337 239942 396948 239944
rect 395337 239939 395403 239942
rect 396942 239940 396948 239942
rect 397012 239940 397018 240004
rect 580073 232386 580139 232389
rect 583520 232386 584960 232476
rect 580073 232384 584960 232386
rect 580073 232328 580078 232384
rect 580134 232328 584960 232384
rect 580073 232326 584960 232328
rect 580073 232323 580139 232326
rect 583520 232236 584960 232326
rect 394601 232114 394667 232117
rect 396758 232114 396764 232116
rect 394601 232112 396764 232114
rect 394601 232056 394606 232112
rect 394662 232056 396764 232112
rect 394601 232054 396764 232056
rect 394601 232051 394667 232054
rect 396758 232052 396764 232054
rect 396828 232052 396834 232116
rect 390369 231162 390435 231165
rect 396942 231162 396948 231164
rect 390369 231160 396948 231162
rect 390369 231104 390374 231160
rect 390430 231104 396948 231160
rect 390369 231102 396948 231104
rect 390369 231099 390435 231102
rect 396942 231100 396948 231102
rect 397012 231100 397018 231164
rect -960 227884 480 228124
rect 579797 219058 579863 219061
rect 583520 219058 584960 219148
rect 579797 219056 584960 219058
rect 579797 219000 579802 219056
rect 579858 219000 584960 219056
rect 579797 218998 584960 219000
rect 579797 218995 579863 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 3141 214978 3207 214981
rect -960 214976 3207 214978
rect -960 214920 3146 214976
rect 3202 214920 3207 214976
rect -960 214918 3207 214920
rect -960 214828 480 214918
rect 3141 214915 3207 214918
rect 579981 205730 580047 205733
rect 583520 205730 584960 205820
rect 579981 205728 584960 205730
rect 579981 205672 579986 205728
rect 580042 205672 584960 205728
rect 579981 205670 584960 205672
rect 579981 205667 580047 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3141 201922 3207 201925
rect -960 201920 3207 201922
rect -960 201864 3146 201920
rect 3202 201864 3207 201920
rect -960 201862 3207 201864
rect -960 201772 480 201862
rect 3141 201859 3207 201862
rect 138105 195938 138171 195941
rect 140405 195938 140471 195941
rect 138105 195936 140471 195938
rect 138105 195880 138110 195936
rect 138166 195880 140410 195936
rect 140466 195880 140471 195936
rect 138105 195878 140471 195880
rect 138105 195875 138171 195878
rect 140405 195875 140471 195878
rect 141417 195938 141483 195941
rect 160829 195938 160895 195941
rect 141417 195936 144194 195938
rect 141417 195880 141422 195936
rect 141478 195880 144194 195936
rect 141417 195878 144194 195880
rect 141417 195875 141483 195878
rect 144134 195644 144194 195878
rect 158854 195936 160895 195938
rect 158854 195928 160834 195936
rect 158854 195872 158902 195928
rect 158958 195880 160834 195928
rect 160890 195880 160895 195936
rect 158958 195878 160895 195880
rect 158958 195872 158963 195878
rect 160829 195875 160895 195878
rect 158854 195870 158963 195872
rect 158897 195867 158963 195870
rect 157149 195666 157215 195669
rect 155910 195664 157215 195666
rect 155910 195608 157154 195664
rect 157210 195608 157215 195664
rect 155910 195606 157215 195608
rect 139393 195530 139459 195533
rect 139393 195528 142170 195530
rect 139393 195472 139398 195528
rect 139454 195498 142170 195528
rect 139454 195472 142692 195498
rect 139393 195470 142692 195472
rect 139393 195467 139459 195470
rect 142110 195438 142692 195470
rect 155910 195340 155970 195606
rect 157149 195603 157215 195606
rect 143390 193292 143396 193356
rect 143460 193354 143466 193356
rect 155166 193354 155172 193356
rect 143460 193294 155172 193354
rect 143460 193292 143466 193294
rect 155166 193292 155172 193294
rect 155236 193292 155242 193356
rect 579889 192538 579955 192541
rect 583520 192538 584960 192628
rect 579889 192536 584960 192538
rect 579889 192480 579894 192536
rect 579950 192480 584960 192536
rect 579889 192478 584960 192480
rect 579889 192475 579955 192478
rect 583520 192388 584960 192478
rect 140865 191858 140931 191861
rect 143214 191858 143980 191900
rect 140865 191856 143980 191858
rect 140865 191800 140870 191856
rect 140926 191840 143980 191856
rect 140926 191800 143274 191840
rect 140865 191798 143274 191800
rect 140865 191795 140931 191798
rect 140773 191722 140839 191725
rect 143398 191722 143980 191760
rect 140773 191720 143980 191722
rect 140773 191664 140778 191720
rect 140834 191700 143980 191720
rect 140834 191664 143458 191700
rect 140773 191662 143458 191664
rect 140773 191659 140839 191662
rect 143574 191568 143580 191632
rect 143644 191630 143650 191632
rect 143644 191570 144164 191630
rect 143644 191568 143650 191570
rect 140957 190906 141023 190909
rect 144134 190906 144194 191460
rect 144361 191042 144427 191045
rect 144494 191042 144500 191044
rect 144361 191040 144500 191042
rect 144361 190984 144366 191040
rect 144422 190984 144500 191040
rect 144361 190982 144500 190984
rect 144361 190979 144427 190982
rect 144494 190980 144500 190982
rect 144564 190980 144570 191044
rect 140957 190904 144194 190906
rect 140957 190848 140962 190904
rect 141018 190848 144194 190904
rect 140957 190846 144194 190848
rect 140957 190843 141023 190846
rect 145833 189820 145899 189821
rect 145782 189818 145788 189820
rect 145742 189758 145788 189818
rect 145852 189816 145899 189820
rect 145894 189760 145899 189816
rect 145782 189756 145788 189758
rect 145852 189756 145899 189760
rect 145833 189755 145899 189756
rect 144494 189212 144500 189276
rect 144564 189274 144570 189276
rect 144821 189274 144887 189277
rect 144564 189272 144887 189274
rect 144564 189216 144826 189272
rect 144882 189216 144887 189272
rect 144564 189214 144887 189216
rect 144564 189212 144570 189214
rect 144821 189211 144887 189214
rect -960 188866 480 188956
rect 155166 188940 155172 189004
rect 155236 189002 155242 189004
rect 157333 189002 157399 189005
rect 155236 189000 157399 189002
rect 155236 188944 157338 189000
rect 157394 188944 157399 189000
rect 155236 188942 157399 188944
rect 155236 188940 155242 188942
rect 157333 188939 157399 188942
rect 3141 188866 3207 188869
rect -960 188864 3207 188866
rect -960 188808 3146 188864
rect 3202 188808 3207 188864
rect -960 188806 3207 188808
rect -960 188716 480 188806
rect 3141 188803 3207 188806
rect 140957 184378 141023 184381
rect 141182 184378 141188 184380
rect 140957 184376 141188 184378
rect 140957 184320 140962 184376
rect 141018 184320 141188 184376
rect 140957 184318 141188 184320
rect 140957 184315 141023 184318
rect 141182 184316 141188 184318
rect 141252 184316 141258 184380
rect 140773 184244 140839 184245
rect 140773 184240 140820 184244
rect 140884 184242 140890 184244
rect 140773 184184 140778 184240
rect 140773 184180 140820 184184
rect 140884 184182 140930 184242
rect 140884 184180 140890 184182
rect 140773 184179 140839 184180
rect 140865 184106 140931 184109
rect 142838 184106 142844 184108
rect 140865 184104 142844 184106
rect 140865 184048 140870 184104
rect 140926 184048 142844 184104
rect 140865 184046 142844 184048
rect 140865 184043 140931 184046
rect 142838 184044 142844 184046
rect 142908 184044 142914 184108
rect 144913 182066 144979 182069
rect 147254 182066 147260 182068
rect 144913 182064 147260 182066
rect 144913 182008 144918 182064
rect 144974 182008 147260 182064
rect 144913 182006 147260 182008
rect 144913 182003 144979 182006
rect 147254 182004 147260 182006
rect 147324 182004 147330 182068
rect 143390 181250 143396 181252
rect 141374 181190 143396 181250
rect 141233 181114 141299 181117
rect 141374 181114 141434 181190
rect 143390 181188 143396 181190
rect 143460 181188 143466 181252
rect 141233 181112 141434 181114
rect 141233 181056 141238 181112
rect 141294 181056 141434 181112
rect 141233 181054 141434 181056
rect 141233 181051 141299 181054
rect 143390 180916 143396 180980
rect 143460 180978 143466 180980
rect 144637 180978 144703 180981
rect 143460 180976 144703 180978
rect 143460 180920 144642 180976
rect 144698 180920 144703 180976
rect 143460 180918 144703 180920
rect 143460 180916 143466 180918
rect 144637 180915 144703 180918
rect 579981 179210 580047 179213
rect 583520 179210 584960 179300
rect 579981 179208 584960 179210
rect 579981 179152 579986 179208
rect 580042 179152 584960 179208
rect 579981 179150 584960 179152
rect 579981 179147 580047 179150
rect 142286 179012 142292 179076
rect 142356 179074 142362 179076
rect 142661 179074 142727 179077
rect 142356 179072 142727 179074
rect 142356 179016 142666 179072
rect 142722 179016 142727 179072
rect 583520 179060 584960 179150
rect 142356 179014 142727 179016
rect 142356 179012 142362 179014
rect 142661 179011 142727 179014
rect 142838 178876 142844 178940
rect 142908 178938 142914 178940
rect 144085 178938 144151 178941
rect 142908 178936 144151 178938
rect 142908 178880 144090 178936
rect 144146 178880 144151 178936
rect 142908 178878 144151 178880
rect 142908 178876 142914 178878
rect 144085 178875 144151 178878
rect 141182 178740 141188 178804
rect 141252 178802 141258 178804
rect 141693 178802 141759 178805
rect 141252 178800 141759 178802
rect 141252 178744 141698 178800
rect 141754 178744 141759 178800
rect 141252 178742 141759 178744
rect 141252 178740 141258 178742
rect 141693 178739 141759 178742
rect 140814 178604 140820 178668
rect 140884 178666 140890 178668
rect 141785 178666 141851 178669
rect 140884 178664 141851 178666
rect 140884 178608 141790 178664
rect 141846 178608 141851 178664
rect 140884 178606 141851 178608
rect 140884 178604 140890 178606
rect 141785 178603 141851 178606
rect 157793 178122 157859 178125
rect 158529 178122 158595 178125
rect 157793 178120 158595 178122
rect 157793 178064 157798 178120
rect 157854 178064 158534 178120
rect 158590 178064 158595 178120
rect 157793 178062 158595 178064
rect 157793 178059 157859 178062
rect 158529 178059 158595 178062
rect -960 175796 480 176036
rect 147254 174524 147260 174588
rect 147324 174586 147330 174588
rect 147489 174586 147555 174589
rect 147324 174584 147555 174586
rect 147324 174528 147494 174584
rect 147550 174528 147555 174584
rect 147324 174526 147555 174528
rect 147324 174524 147330 174526
rect 147489 174523 147555 174526
rect 579797 165882 579863 165885
rect 583520 165882 584960 165972
rect 579797 165880 584960 165882
rect 579797 165824 579802 165880
rect 579858 165824 584960 165880
rect 579797 165822 584960 165824
rect 579797 165819 579863 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3141 162890 3207 162893
rect -960 162888 3207 162890
rect -960 162832 3146 162888
rect 3202 162832 3207 162888
rect -960 162830 3207 162832
rect -960 162740 480 162830
rect 3141 162827 3207 162830
rect 580441 152690 580507 152693
rect 583520 152690 584960 152780
rect 580441 152688 584960 152690
rect 580441 152632 580446 152688
rect 580502 152632 584960 152688
rect 580441 152630 584960 152632
rect 580441 152627 580507 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3141 149834 3207 149837
rect -960 149832 3207 149834
rect -960 149776 3146 149832
rect 3202 149776 3207 149832
rect -960 149774 3207 149776
rect -960 149684 480 149774
rect 3141 149771 3207 149774
rect 579613 139362 579679 139365
rect 583520 139362 584960 139452
rect 579613 139360 584960 139362
rect 579613 139304 579618 139360
rect 579674 139304 584960 139360
rect 579613 139302 584960 139304
rect 579613 139299 579679 139302
rect 583520 139212 584960 139302
rect 139669 138002 139735 138005
rect 141918 138002 141924 138004
rect 139669 138000 141924 138002
rect 139669 137944 139674 138000
rect 139730 137944 141924 138000
rect 139669 137942 141924 137944
rect 139669 137939 139735 137942
rect 141918 137940 141924 137942
rect 141988 137940 141994 138004
rect 143574 137668 143580 137732
rect 143644 137730 143650 137732
rect 161565 137730 161631 137733
rect 143644 137728 161631 137730
rect 143644 137672 161570 137728
rect 161626 137672 161631 137728
rect 143644 137670 161631 137672
rect 143644 137668 143650 137670
rect 161565 137667 161631 137670
rect 146150 137532 146156 137596
rect 146220 137594 146226 137596
rect 167821 137594 167887 137597
rect 146220 137592 167887 137594
rect 146220 137536 167826 137592
rect 167882 137536 167887 137592
rect 146220 137534 167887 137536
rect 146220 137532 146226 137534
rect 167821 137531 167887 137534
rect 143390 137396 143396 137460
rect 143460 137458 143466 137460
rect 169385 137458 169451 137461
rect 143460 137456 169451 137458
rect 143460 137400 169390 137456
rect 169446 137400 169451 137456
rect 143460 137398 169451 137400
rect 143460 137396 143466 137398
rect 169385 137395 169451 137398
rect 114001 137322 114067 137325
rect 396574 137322 396580 137324
rect 114001 137320 396580 137322
rect 114001 137264 114006 137320
rect 114062 137264 396580 137320
rect 114001 137262 396580 137264
rect 114001 137259 114067 137262
rect 396574 137260 396580 137262
rect 396644 137260 396650 137324
rect -960 136778 480 136868
rect 3417 136778 3483 136781
rect -960 136776 3483 136778
rect -960 136720 3422 136776
rect 3478 136720 3483 136776
rect -960 136718 3483 136720
rect -960 136628 480 136718
rect 3417 136715 3483 136718
rect 115105 133242 115171 133245
rect 115105 133240 116226 133242
rect 115105 133184 115110 133240
rect 115166 133184 116226 133240
rect 115105 133182 116226 133184
rect 115105 133179 115171 133182
rect 116166 132600 116226 133182
rect 175598 132429 175658 132600
rect 175549 132424 175658 132429
rect 175549 132368 175554 132424
rect 175610 132368 175658 132424
rect 175549 132366 175658 132368
rect 175549 132363 175615 132366
rect 113725 131202 113791 131205
rect 178585 131202 178651 131205
rect 113725 131200 116226 131202
rect 113725 131144 113730 131200
rect 113786 131144 116226 131200
rect 113725 131142 116226 131144
rect 113725 131139 113791 131142
rect 116166 131104 116226 131142
rect 175782 131200 178651 131202
rect 175782 131144 178590 131200
rect 178646 131144 178651 131200
rect 175782 131142 178651 131144
rect 175782 131104 175842 131142
rect 178585 131139 178651 131142
rect 175365 129978 175431 129981
rect 175365 129976 175474 129978
rect 175365 129920 175370 129976
rect 175426 129920 175474 129976
rect 175365 129915 175474 129920
rect 175414 129608 175474 129915
rect 113725 129026 113791 129029
rect 116166 129026 116226 129608
rect 113725 129024 116226 129026
rect 113725 128968 113730 129024
rect 113786 128968 116226 129024
rect 113725 128966 116226 128968
rect 113725 128963 113791 128966
rect 175365 128346 175431 128349
rect 175365 128344 175474 128346
rect 175365 128288 175370 128344
rect 175426 128288 175474 128344
rect 175365 128283 175474 128288
rect 175414 128112 175474 128283
rect 113633 127530 113699 127533
rect 116166 127530 116226 128112
rect 113633 127528 116226 127530
rect 113633 127472 113638 127528
rect 113694 127472 116226 127528
rect 113633 127470 116226 127472
rect 113633 127467 113699 127470
rect 175641 126986 175707 126989
rect 175598 126984 175707 126986
rect 175598 126928 175646 126984
rect 175702 126928 175707 126984
rect 175598 126923 175707 126928
rect 113725 126850 113791 126853
rect 113725 126848 116226 126850
rect 113725 126792 113730 126848
rect 113786 126792 116226 126848
rect 113725 126790 116226 126792
rect 113725 126787 113791 126790
rect 116166 126616 116226 126790
rect 175598 126616 175658 126923
rect 579705 126034 579771 126037
rect 583520 126034 584960 126124
rect 579705 126032 584960 126034
rect 579705 125976 579710 126032
rect 579766 125976 584960 126032
rect 579705 125974 584960 125976
rect 579705 125971 579771 125974
rect 583520 125884 584960 125974
rect 178861 125490 178927 125493
rect 175782 125488 178927 125490
rect 175782 125432 178866 125488
rect 178922 125432 178927 125488
rect 175782 125430 178927 125432
rect 113541 125354 113607 125357
rect 113541 125352 116226 125354
rect 113541 125296 113546 125352
rect 113602 125296 116226 125352
rect 113541 125294 116226 125296
rect 113541 125291 113607 125294
rect 116166 125120 116226 125294
rect 175782 125120 175842 125430
rect 178861 125427 178927 125430
rect 178493 124130 178559 124133
rect 175782 124128 178559 124130
rect 175782 124072 178498 124128
rect 178554 124072 178559 124128
rect 175782 124070 178559 124072
rect 113725 123858 113791 123861
rect 113725 123856 116226 123858
rect -960 123572 480 123812
rect 113725 123800 113730 123856
rect 113786 123800 116226 123856
rect 113725 123798 116226 123800
rect 113725 123795 113791 123798
rect 116166 123624 116226 123798
rect 175782 123624 175842 124070
rect 178493 124067 178559 124070
rect 113357 122770 113423 122773
rect 113357 122768 116226 122770
rect 113357 122712 113362 122768
rect 113418 122712 116226 122768
rect 113357 122710 116226 122712
rect 113357 122707 113423 122710
rect 116166 122128 116226 122710
rect 178769 122498 178835 122501
rect 175782 122496 178835 122498
rect 175782 122440 178774 122496
rect 178830 122440 178835 122496
rect 175782 122438 178835 122440
rect 175782 122128 175842 122438
rect 178769 122435 178835 122438
rect 113725 121274 113791 121277
rect 177849 121274 177915 121277
rect 113725 121272 116226 121274
rect 113725 121216 113730 121272
rect 113786 121216 116226 121272
rect 113725 121214 116226 121216
rect 113725 121211 113791 121214
rect 116166 120632 116226 121214
rect 175782 121272 177915 121274
rect 175782 121216 177854 121272
rect 177910 121216 177915 121272
rect 175782 121214 177915 121216
rect 175782 120632 175842 121214
rect 177849 121211 177915 121214
rect 113725 119778 113791 119781
rect 178401 119778 178467 119781
rect 113725 119776 116226 119778
rect 113725 119720 113730 119776
rect 113786 119720 116226 119776
rect 113725 119718 116226 119720
rect 113725 119715 113791 119718
rect 116166 119136 116226 119718
rect 175782 119776 178467 119778
rect 175782 119720 178406 119776
rect 178462 119720 178467 119776
rect 175782 119718 178467 119720
rect 175782 119136 175842 119718
rect 178401 119715 178467 119718
rect 113633 118282 113699 118285
rect 178033 118282 178099 118285
rect 113633 118280 116226 118282
rect 113633 118224 113638 118280
rect 113694 118224 116226 118280
rect 113633 118222 116226 118224
rect 113633 118219 113699 118222
rect 116166 117640 116226 118222
rect 175782 118280 178099 118282
rect 175782 118224 178038 118280
rect 178094 118224 178099 118280
rect 175782 118222 178099 118224
rect 175782 117640 175842 118222
rect 178033 118219 178099 118222
rect 113725 116786 113791 116789
rect 178677 116786 178743 116789
rect 113725 116784 116226 116786
rect 113725 116728 113730 116784
rect 113786 116728 116226 116784
rect 113725 116726 116226 116728
rect 113725 116723 113791 116726
rect 116166 116144 116226 116726
rect 175782 116784 178743 116786
rect 175782 116728 178682 116784
rect 178738 116728 178743 116784
rect 175782 116726 178743 116728
rect 175782 116144 175842 116726
rect 178677 116723 178743 116726
rect 113725 115290 113791 115293
rect 178309 115290 178375 115293
rect 113725 115288 116226 115290
rect 113725 115232 113730 115288
rect 113786 115232 116226 115288
rect 113725 115230 116226 115232
rect 113725 115227 113791 115230
rect 116166 114648 116226 115230
rect 175782 115288 178375 115290
rect 175782 115232 178314 115288
rect 178370 115232 178375 115288
rect 175782 115230 178375 115232
rect 175782 114648 175842 115230
rect 178309 115227 178375 115230
rect 113725 113114 113791 113117
rect 116166 113114 116226 113152
rect 113725 113112 116226 113114
rect 113725 113056 113730 113112
rect 113786 113056 116226 113112
rect 113725 113054 116226 113056
rect 175782 113114 175842 113152
rect 178125 113114 178191 113117
rect 175782 113112 178191 113114
rect 175782 113056 178130 113112
rect 178186 113056 178191 113112
rect 175782 113054 178191 113056
rect 113725 113051 113791 113054
rect 178125 113051 178191 113054
rect 580533 112842 580599 112845
rect 583520 112842 584960 112932
rect 580533 112840 584960 112842
rect 580533 112784 580538 112840
rect 580594 112784 584960 112840
rect 580533 112782 584960 112784
rect 580533 112779 580599 112782
rect 583520 112692 584960 112782
rect 175457 111890 175523 111893
rect 175414 111888 175523 111890
rect 175414 111832 175462 111888
rect 175518 111832 175523 111888
rect 175414 111827 175523 111832
rect 113725 111754 113791 111757
rect 113725 111752 116226 111754
rect 113725 111696 113730 111752
rect 113786 111696 116226 111752
rect 113725 111694 116226 111696
rect 113725 111691 113791 111694
rect 116166 111656 116226 111694
rect 175414 111656 175474 111827
rect -960 110666 480 110756
rect 3785 110666 3851 110669
rect -960 110664 3851 110666
rect -960 110608 3790 110664
rect 3846 110608 3851 110664
rect -960 110606 3851 110608
rect -960 110516 480 110606
rect 3785 110603 3851 110606
rect 113725 110394 113791 110397
rect 178033 110394 178099 110397
rect 113725 110392 116226 110394
rect 113725 110336 113730 110392
rect 113786 110336 116226 110392
rect 113725 110334 116226 110336
rect 113725 110331 113791 110334
rect 116166 110160 116226 110334
rect 175782 110392 178099 110394
rect 175782 110336 178038 110392
rect 178094 110336 178099 110392
rect 175782 110334 178099 110336
rect 175782 110160 175842 110334
rect 178033 110331 178099 110334
rect 178217 109034 178283 109037
rect 175782 109032 178283 109034
rect 175782 108976 178222 109032
rect 178278 108976 178283 109032
rect 175782 108974 178283 108976
rect 113725 108898 113791 108901
rect 113725 108896 116226 108898
rect 113725 108840 113730 108896
rect 113786 108840 116226 108896
rect 113725 108838 116226 108840
rect 113725 108835 113791 108838
rect 116166 108664 116226 108838
rect 175782 108664 175842 108974
rect 178217 108971 178283 108974
rect 176745 107538 176811 107541
rect 175782 107536 176811 107538
rect 175782 107480 176750 107536
rect 176806 107480 176811 107536
rect 175782 107478 176811 107480
rect 113541 107402 113607 107405
rect 113541 107400 116226 107402
rect 113541 107344 113546 107400
rect 113602 107344 116226 107400
rect 113541 107342 116226 107344
rect 113541 107339 113607 107342
rect 116166 107168 116226 107342
rect 175782 107168 175842 107478
rect 176745 107475 176811 107478
rect 113725 106178 113791 106181
rect 113725 106176 116226 106178
rect 113725 106120 113730 106176
rect 113786 106120 116226 106176
rect 113725 106118 116226 106120
rect 113725 106115 113791 106118
rect 116166 105672 116226 106118
rect 178033 106042 178099 106045
rect 175782 106040 178099 106042
rect 175782 105984 178038 106040
rect 178094 105984 178099 106040
rect 175782 105982 178099 105984
rect 175782 105672 175842 105982
rect 178033 105979 178099 105982
rect 113357 104818 113423 104821
rect 113357 104816 116226 104818
rect 113357 104760 113362 104816
rect 113418 104760 116226 104816
rect 113357 104758 116226 104760
rect 113357 104755 113423 104758
rect 116166 104176 116226 104758
rect 178033 104546 178099 104549
rect 175782 104544 178099 104546
rect 175782 104488 178038 104544
rect 178094 104488 178099 104544
rect 175782 104486 178099 104488
rect 175782 104176 175842 104486
rect 178033 104483 178099 104486
rect 115289 103186 115355 103189
rect 115289 103184 116226 103186
rect 115289 103128 115294 103184
rect 115350 103128 116226 103184
rect 115289 103126 116226 103128
rect 115289 103123 115355 103126
rect 116166 102680 116226 103126
rect 178033 103050 178099 103053
rect 175782 103048 178099 103050
rect 175782 102992 178038 103048
rect 178094 102992 178099 103048
rect 175782 102990 178099 102992
rect 175782 102680 175842 102990
rect 178033 102987 178099 102990
rect 113817 101826 113883 101829
rect 113817 101824 116226 101826
rect 113817 101768 113822 101824
rect 113878 101768 116226 101824
rect 113817 101766 116226 101768
rect 113817 101763 113883 101766
rect 116166 101184 116226 101766
rect 178033 101690 178099 101693
rect 175782 101688 178099 101690
rect 175782 101632 178038 101688
rect 178094 101632 178099 101688
rect 175782 101630 178099 101632
rect 175782 101184 175842 101630
rect 178033 101627 178099 101630
rect 115933 100330 115999 100333
rect 115933 100328 116226 100330
rect 115933 100272 115938 100328
rect 115994 100272 116226 100328
rect 115933 100270 116226 100272
rect 115933 100267 115999 100270
rect 116166 99688 116226 100270
rect 178033 100194 178099 100197
rect 175782 100192 178099 100194
rect 175782 100136 178038 100192
rect 178094 100136 178099 100192
rect 175782 100134 178099 100136
rect 175782 99688 175842 100134
rect 178033 100131 178099 100134
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect 113909 98834 113975 98837
rect 178033 98834 178099 98837
rect 113909 98832 116226 98834
rect 113909 98776 113914 98832
rect 113970 98776 116226 98832
rect 113909 98774 116226 98776
rect 113909 98771 113975 98774
rect 116166 98192 116226 98774
rect 175782 98832 178099 98834
rect 175782 98776 178038 98832
rect 178094 98776 178099 98832
rect 175782 98774 178099 98776
rect 175782 98192 175842 98774
rect 178033 98771 178099 98774
rect -960 97610 480 97700
rect 3693 97610 3759 97613
rect -960 97608 3759 97610
rect -960 97552 3698 97608
rect 3754 97552 3759 97608
rect -960 97550 3759 97552
rect -960 97460 480 97550
rect 3693 97547 3759 97550
rect 178033 97338 178099 97341
rect 175782 97336 178099 97338
rect 175782 97280 178038 97336
rect 178094 97280 178099 97336
rect 175782 97278 178099 97280
rect 115657 96726 115723 96729
rect 115657 96724 116196 96726
rect 115657 96668 115662 96724
rect 115718 96668 116196 96724
rect 175782 96696 175842 97278
rect 178033 97275 178099 97278
rect 115657 96666 116196 96668
rect 115657 96663 115723 96666
rect 115565 95162 115631 95165
rect 116166 95162 116226 95200
rect 115565 95160 116226 95162
rect 115565 95104 115570 95160
rect 115626 95104 116226 95160
rect 115565 95102 116226 95104
rect 175782 95162 175842 95200
rect 178033 95162 178099 95165
rect 175782 95160 178099 95162
rect 175782 95104 178038 95160
rect 178094 95104 178099 95160
rect 175782 95102 178099 95104
rect 115565 95099 115631 95102
rect 178033 95099 178099 95102
rect 115473 93802 115539 93805
rect 178033 93802 178099 93805
rect 115473 93800 116226 93802
rect 115473 93744 115478 93800
rect 115534 93744 116226 93800
rect 115473 93742 116226 93744
rect 115473 93739 115539 93742
rect 116166 93704 116226 93742
rect 175782 93800 178099 93802
rect 175782 93744 178038 93800
rect 178094 93744 178099 93800
rect 175782 93742 178099 93744
rect 175782 93704 175842 93742
rect 178033 93739 178099 93742
rect 115381 92442 115447 92445
rect 115381 92440 116226 92442
rect 115381 92384 115386 92440
rect 115442 92384 116226 92440
rect 115381 92382 116226 92384
rect 115381 92379 115447 92382
rect 116166 92208 116226 92382
rect 178033 92306 178099 92309
rect 175782 92304 178099 92306
rect 175782 92248 178038 92304
rect 178094 92248 178099 92304
rect 175782 92246 178099 92248
rect 175782 92208 175842 92246
rect 178033 92243 178099 92246
rect 114001 91082 114067 91085
rect 114001 91080 116226 91082
rect 114001 91024 114006 91080
rect 114062 91024 116226 91080
rect 114001 91022 116226 91024
rect 114001 91019 114067 91022
rect 116166 90712 116226 91022
rect 178033 90946 178099 90949
rect 175782 90944 178099 90946
rect 175782 90888 178038 90944
rect 178094 90888 178099 90944
rect 175782 90886 178099 90888
rect 175782 90712 175842 90886
rect 178033 90883 178099 90886
rect 114093 89722 114159 89725
rect 114093 89720 116226 89722
rect 114093 89664 114098 89720
rect 114154 89664 116226 89720
rect 114093 89662 116226 89664
rect 114093 89659 114159 89662
rect 116166 89216 116226 89662
rect 178033 89450 178099 89453
rect 175782 89448 178099 89450
rect 175782 89392 178038 89448
rect 178094 89392 178099 89448
rect 175782 89390 178099 89392
rect 175782 89216 175842 89390
rect 178033 89387 178099 89390
rect 114185 88226 114251 88229
rect 114185 88224 116226 88226
rect 114185 88168 114190 88224
rect 114246 88168 116226 88224
rect 114185 88166 116226 88168
rect 114185 88163 114251 88166
rect 116166 87720 116226 88166
rect 178033 88090 178099 88093
rect 175782 88088 178099 88090
rect 175782 88032 178038 88088
rect 178094 88032 178099 88088
rect 175782 88030 178099 88032
rect 175782 87720 175842 88030
rect 178033 88027 178099 88030
rect 114277 86866 114343 86869
rect 114277 86864 116226 86866
rect 114277 86808 114282 86864
rect 114338 86808 116226 86864
rect 114277 86806 116226 86808
rect 114277 86803 114343 86806
rect 116166 86224 116226 86806
rect 178033 86594 178099 86597
rect 175782 86592 178099 86594
rect 175782 86536 178038 86592
rect 178094 86536 178099 86592
rect 175782 86534 178099 86536
rect 175782 86224 175842 86534
rect 178033 86531 178099 86534
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect 114369 85370 114435 85373
rect 114369 85368 116226 85370
rect 114369 85312 114374 85368
rect 114430 85312 116226 85368
rect 114369 85310 116226 85312
rect 114369 85307 114435 85310
rect -960 84690 480 84780
rect 116166 84728 116226 85310
rect 178033 85098 178099 85101
rect 175782 85096 178099 85098
rect 175782 85040 178038 85096
rect 178094 85040 178099 85096
rect 175782 85038 178099 85040
rect 175782 84728 175842 85038
rect 178033 85035 178099 85038
rect 3325 84690 3391 84693
rect -960 84688 3391 84690
rect -960 84632 3330 84688
rect 3386 84632 3391 84688
rect -960 84630 3391 84632
rect -960 84540 480 84630
rect 3325 84627 3391 84630
rect 178033 83738 178099 83741
rect 175782 83736 178099 83738
rect 175782 83680 178038 83736
rect 178094 83680 178099 83736
rect 175782 83678 178099 83680
rect 115841 83262 115907 83265
rect 115841 83260 116196 83262
rect 115841 83204 115846 83260
rect 115902 83204 116196 83260
rect 175782 83232 175842 83678
rect 178033 83675 178099 83678
rect 115841 83202 116196 83204
rect 115841 83199 115907 83202
rect 178033 82242 178099 82245
rect 175782 82240 178099 82242
rect 175782 82184 178038 82240
rect 178094 82184 178099 82240
rect 175782 82182 178099 82184
rect 115749 81766 115815 81769
rect 115749 81764 116196 81766
rect 115749 81708 115754 81764
rect 115810 81708 116196 81764
rect 175782 81736 175842 82182
rect 178033 82179 178099 82182
rect 115749 81706 116196 81708
rect 115749 81703 115815 81706
rect 114461 80882 114527 80885
rect 178677 80882 178743 80885
rect 114461 80880 116226 80882
rect 114461 80824 114466 80880
rect 114522 80824 116226 80880
rect 114461 80822 116226 80824
rect 114461 80819 114527 80822
rect 116166 80240 116226 80822
rect 175782 80880 178743 80882
rect 175782 80824 178682 80880
rect 178738 80824 178743 80880
rect 175782 80822 178743 80824
rect 175782 80240 175842 80822
rect 178677 80819 178743 80822
rect 116534 78437 116594 78744
rect 175782 78706 175842 78744
rect 178677 78706 178743 78709
rect 175782 78704 178743 78706
rect 175782 78648 178682 78704
rect 178738 78648 178743 78704
rect 175782 78646 178743 78648
rect 178677 78643 178743 78646
rect 116485 78432 116594 78437
rect 116485 78376 116490 78432
rect 116546 78376 116594 78432
rect 116485 78374 116594 78376
rect 116485 78371 116551 78374
rect 114369 76666 114435 76669
rect 116166 76666 116226 77248
rect 114369 76664 116226 76666
rect 114369 76608 114374 76664
rect 114430 76608 116226 76664
rect 114369 76606 116226 76608
rect 175782 76666 175842 77248
rect 178033 76666 178099 76669
rect 175782 76664 178099 76666
rect 175782 76608 178038 76664
rect 178094 76608 178099 76664
rect 175782 76606 178099 76608
rect 114369 76603 114435 76606
rect 178033 76603 178099 76606
rect 114461 75442 114527 75445
rect 116166 75442 116226 75752
rect 116485 75578 116551 75581
rect 175917 75578 175983 75581
rect 116485 75576 175983 75578
rect 116485 75520 116490 75576
rect 116546 75520 175922 75576
rect 175978 75520 175983 75576
rect 116485 75518 175983 75520
rect 116485 75515 116551 75518
rect 175917 75515 175983 75518
rect 114461 75440 116226 75442
rect 114461 75384 114466 75440
rect 114522 75384 116226 75440
rect 114461 75382 116226 75384
rect 114461 75379 114527 75382
rect 168414 75380 168420 75444
rect 168484 75442 168490 75444
rect 171409 75442 171475 75445
rect 168484 75440 171475 75442
rect 168484 75384 171414 75440
rect 171470 75384 171475 75440
rect 168484 75382 171475 75384
rect 168484 75380 168490 75382
rect 171409 75379 171475 75382
rect 103470 75246 122850 75306
rect 4981 75170 5047 75173
rect 103470 75170 103530 75246
rect 4981 75168 103530 75170
rect 4981 75112 4986 75168
rect 5042 75112 103530 75168
rect 4981 75110 103530 75112
rect 122790 75170 122850 75246
rect 167678 75244 167684 75308
rect 167748 75306 167754 75308
rect 168598 75306 168604 75308
rect 167748 75246 168604 75306
rect 167748 75244 167754 75246
rect 168598 75244 168604 75246
rect 168668 75244 168674 75308
rect 171685 75306 171751 75309
rect 168790 75304 171751 75306
rect 168790 75248 171690 75304
rect 171746 75248 171751 75304
rect 168790 75246 171751 75248
rect 168598 75170 168604 75172
rect 122790 75110 168604 75170
rect 4981 75107 5047 75110
rect 168598 75108 168604 75110
rect 168668 75108 168674 75172
rect 4797 75034 4863 75037
rect 168414 75034 168420 75036
rect 4797 75032 157350 75034
rect 4797 74976 4802 75032
rect 4858 74976 157350 75032
rect 4797 74974 157350 74976
rect 4797 74971 4863 74974
rect 157290 74762 157350 74974
rect 167502 74974 168420 75034
rect 167502 74901 167562 74974
rect 168414 74972 168420 74974
rect 168484 74972 168490 75036
rect 162393 74898 162459 74901
rect 162894 74898 162900 74900
rect 162393 74896 162900 74898
rect 162393 74840 162398 74896
rect 162454 74840 162900 74896
rect 162393 74838 162900 74840
rect 162393 74835 162459 74838
rect 162894 74836 162900 74838
rect 162964 74836 162970 74900
rect 167453 74896 167562 74901
rect 167453 74840 167458 74896
rect 167514 74840 167562 74896
rect 167453 74838 167562 74840
rect 167729 74898 167795 74901
rect 168790 74898 168850 75246
rect 171685 75243 171751 75246
rect 579613 75306 579679 75309
rect 580758 75306 580764 75308
rect 579613 75304 580764 75306
rect 579613 75248 579618 75304
rect 579674 75248 580764 75304
rect 579613 75246 580764 75248
rect 579613 75243 579679 75246
rect 580758 75244 580764 75246
rect 580828 75244 580834 75308
rect 167729 74896 168850 74898
rect 167729 74840 167734 74896
rect 167790 74840 168850 74896
rect 167729 74838 168850 74840
rect 168974 74974 176670 75034
rect 167453 74835 167519 74838
rect 167729 74835 167795 74838
rect 167494 74762 167500 74764
rect 157290 74702 167500 74762
rect 167494 74700 167500 74702
rect 167564 74700 167570 74764
rect 167637 74762 167703 74765
rect 168974 74762 169034 74974
rect 169150 74836 169156 74900
rect 169220 74898 169226 74900
rect 169477 74898 169543 74901
rect 169220 74896 169543 74898
rect 169220 74840 169482 74896
rect 169538 74840 169543 74896
rect 169220 74838 169543 74840
rect 169220 74836 169226 74838
rect 169477 74835 169543 74838
rect 169661 74898 169727 74901
rect 170397 74898 170463 74901
rect 169661 74896 170463 74898
rect 169661 74840 169666 74896
rect 169722 74840 170402 74896
rect 170458 74840 170463 74896
rect 169661 74838 170463 74840
rect 176610 74898 176670 74974
rect 396717 74898 396783 74901
rect 176610 74896 396783 74898
rect 176610 74840 396722 74896
rect 396778 74840 396783 74896
rect 176610 74838 396783 74840
rect 169661 74835 169727 74838
rect 170397 74835 170463 74838
rect 396717 74835 396783 74838
rect 167637 74760 169034 74762
rect 167637 74704 167642 74760
rect 167698 74704 169034 74760
rect 167637 74702 169034 74704
rect 169293 74764 169359 74765
rect 169293 74760 169340 74764
rect 169404 74762 169410 74764
rect 580257 74762 580323 74765
rect 169293 74704 169298 74760
rect 167637 74699 167703 74702
rect 169293 74700 169340 74704
rect 169404 74702 169450 74762
rect 169710 74760 580323 74762
rect 169710 74704 580262 74760
rect 580318 74704 580323 74760
rect 169710 74702 580323 74704
rect 169404 74700 169410 74702
rect 169293 74699 169359 74700
rect 151997 74626 152063 74629
rect 157517 74626 157583 74629
rect 151997 74624 157583 74626
rect 151997 74568 152002 74624
rect 152058 74568 157522 74624
rect 157578 74568 157583 74624
rect 151997 74566 157583 74568
rect 151997 74563 152063 74566
rect 157517 74563 157583 74566
rect 168097 74626 168163 74629
rect 169710 74626 169770 74702
rect 580257 74699 580323 74702
rect 168097 74624 169770 74626
rect 168097 74568 168102 74624
rect 168158 74568 169770 74624
rect 168097 74566 169770 74568
rect 171685 74626 171751 74629
rect 580901 74626 580967 74629
rect 171685 74624 580967 74626
rect 171685 74568 171690 74624
rect 171746 74568 580906 74624
rect 580962 74568 580967 74624
rect 171685 74566 580967 74568
rect 168097 74563 168163 74566
rect 171685 74563 171751 74566
rect 580901 74563 580967 74566
rect 3366 74428 3372 74492
rect 3436 74490 3442 74492
rect 167177 74490 167243 74493
rect 168189 74490 168255 74493
rect 3436 74430 167010 74490
rect 3436 74428 3442 74430
rect 3509 74354 3575 74357
rect 161657 74354 161723 74357
rect 162393 74354 162459 74357
rect 3509 74352 157350 74354
rect 3509 74296 3514 74352
rect 3570 74296 157350 74352
rect 3509 74294 157350 74296
rect 3509 74291 3575 74294
rect 157290 74218 157350 74294
rect 161657 74352 162459 74354
rect 161657 74296 161662 74352
rect 161718 74296 162398 74352
rect 162454 74296 162459 74352
rect 161657 74294 162459 74296
rect 166950 74354 167010 74430
rect 167177 74488 168255 74490
rect 167177 74432 167182 74488
rect 167238 74432 168194 74488
rect 168250 74432 168255 74488
rect 167177 74430 168255 74432
rect 167177 74427 167243 74430
rect 168189 74427 168255 74430
rect 169109 74354 169175 74357
rect 166950 74352 169175 74354
rect 166950 74296 169114 74352
rect 169170 74296 169175 74352
rect 166950 74294 169175 74296
rect 161657 74291 161723 74294
rect 162393 74291 162459 74294
rect 169109 74291 169175 74294
rect 167269 74218 167335 74221
rect 579889 74218 579955 74221
rect 157290 74158 167010 74218
rect 6913 74082 6979 74085
rect 166950 74082 167010 74158
rect 167269 74216 579955 74218
rect 167269 74160 167274 74216
rect 167330 74160 579894 74216
rect 579950 74160 579955 74216
rect 167269 74158 579955 74160
rect 167269 74155 167335 74158
rect 579889 74155 579955 74158
rect 169201 74082 169267 74085
rect 6913 74080 162226 74082
rect 6913 74024 6918 74080
rect 6974 74024 162226 74080
rect 6913 74022 162226 74024
rect 166950 74080 169267 74082
rect 166950 74024 169206 74080
rect 169262 74024 169267 74080
rect 166950 74022 169267 74024
rect 6913 74019 6979 74022
rect 4889 73946 4955 73949
rect 162166 73946 162226 74022
rect 169201 74019 169267 74022
rect 169017 73946 169083 73949
rect 4889 73944 157350 73946
rect 4889 73888 4894 73944
rect 4950 73888 157350 73944
rect 4889 73886 157350 73888
rect 162166 73944 169083 73946
rect 162166 73888 169022 73944
rect 169078 73888 169083 73944
rect 162166 73886 169083 73888
rect 4889 73883 4955 73886
rect 157290 73538 157350 73886
rect 169017 73883 169083 73886
rect 168189 73810 168255 73813
rect 580441 73810 580507 73813
rect 168189 73808 580507 73810
rect 168189 73752 168194 73808
rect 168250 73752 580446 73808
rect 580502 73752 580507 73808
rect 168189 73750 580507 73752
rect 168189 73747 168255 73750
rect 580441 73747 580507 73750
rect 167361 73674 167427 73677
rect 580073 73674 580139 73677
rect 167361 73672 580139 73674
rect 167361 73616 167366 73672
rect 167422 73616 580078 73672
rect 580134 73616 580139 73672
rect 167361 73614 580139 73616
rect 167361 73611 167427 73614
rect 580073 73611 580139 73614
rect 169385 73538 169451 73541
rect 157290 73536 169451 73538
rect 157290 73480 169390 73536
rect 169446 73480 169451 73536
rect 157290 73478 169451 73480
rect 169385 73475 169451 73478
rect 162393 73266 162459 73269
rect 162393 73264 166090 73266
rect 162393 73208 162398 73264
rect 162454 73208 166090 73264
rect 162393 73206 166090 73208
rect 162393 73203 162459 73206
rect 128537 73132 128603 73133
rect 128486 73130 128492 73132
rect 128446 73070 128492 73130
rect 128556 73128 128603 73132
rect 128598 73072 128603 73128
rect 128486 73068 128492 73070
rect 128556 73068 128603 73072
rect 128537 73067 128603 73068
rect 161289 73130 161355 73133
rect 162393 73130 162459 73133
rect 161289 73128 162459 73130
rect 161289 73072 161294 73128
rect 161350 73072 162398 73128
rect 162454 73072 162459 73128
rect 161289 73070 162459 73072
rect 161289 73067 161355 73070
rect 162393 73067 162459 73070
rect 163037 73130 163103 73133
rect 166030 73130 166090 73206
rect 167494 73130 167500 73132
rect 163037 73128 165906 73130
rect 163037 73072 163042 73128
rect 163098 73072 165906 73128
rect 163037 73070 165906 73072
rect 166030 73070 167500 73130
rect 163037 73067 163103 73070
rect 149462 72932 149468 72996
rect 149532 72994 149538 72996
rect 150157 72994 150223 72997
rect 149532 72992 150223 72994
rect 149532 72936 150162 72992
rect 150218 72936 150223 72992
rect 149532 72934 150223 72936
rect 149532 72932 149538 72934
rect 150157 72931 150223 72934
rect 153878 72932 153884 72996
rect 153948 72994 153954 72996
rect 154297 72994 154363 72997
rect 153948 72992 154363 72994
rect 153948 72936 154302 72992
rect 154358 72936 154363 72992
rect 153948 72934 154363 72936
rect 153948 72932 153954 72934
rect 154297 72931 154363 72934
rect 162158 72932 162164 72996
rect 162228 72994 162234 72996
rect 162577 72994 162643 72997
rect 162228 72992 162643 72994
rect 162228 72936 162582 72992
rect 162638 72936 162643 72992
rect 162228 72934 162643 72936
rect 162228 72932 162234 72934
rect 162577 72931 162643 72934
rect 163313 72994 163379 72997
rect 165846 72994 165906 73070
rect 167494 73068 167500 73070
rect 167564 73068 167570 73132
rect 168005 73130 168071 73133
rect 580349 73130 580415 73133
rect 168005 73128 580415 73130
rect 168005 73072 168010 73128
rect 168066 73072 580354 73128
rect 580410 73072 580415 73128
rect 168005 73070 580415 73072
rect 168005 73067 168071 73070
rect 580349 73067 580415 73070
rect 167678 72994 167684 72996
rect 163313 72992 165722 72994
rect 163313 72936 163318 72992
rect 163374 72936 165722 72992
rect 163313 72934 165722 72936
rect 165846 72934 167684 72994
rect 163313 72931 163379 72934
rect 148726 72796 148732 72860
rect 148796 72858 148802 72860
rect 148961 72858 149027 72861
rect 148796 72856 149027 72858
rect 148796 72800 148966 72856
rect 149022 72800 149027 72856
rect 148796 72798 149027 72800
rect 148796 72796 148802 72798
rect 148961 72795 149027 72798
rect 149830 72796 149836 72860
rect 149900 72858 149906 72860
rect 150341 72858 150407 72861
rect 149900 72856 150407 72858
rect 149900 72800 150346 72856
rect 150402 72800 150407 72856
rect 149900 72798 150407 72800
rect 149900 72796 149906 72798
rect 150341 72795 150407 72798
rect 151486 72796 151492 72860
rect 151556 72858 151562 72860
rect 151721 72858 151787 72861
rect 151556 72856 151787 72858
rect 151556 72800 151726 72856
rect 151782 72800 151787 72856
rect 151556 72798 151787 72800
rect 151556 72796 151562 72798
rect 151721 72795 151787 72798
rect 152774 72796 152780 72860
rect 152844 72858 152850 72860
rect 152917 72858 152983 72861
rect 152844 72856 152983 72858
rect 152844 72800 152922 72856
rect 152978 72800 152983 72856
rect 152844 72798 152983 72800
rect 152844 72796 152850 72798
rect 152917 72795 152983 72798
rect 154113 72858 154179 72861
rect 154430 72858 154436 72860
rect 154113 72856 154436 72858
rect 154113 72800 154118 72856
rect 154174 72800 154436 72856
rect 154113 72798 154436 72800
rect 154113 72795 154179 72798
rect 154430 72796 154436 72798
rect 154500 72796 154506 72860
rect 155534 72796 155540 72860
rect 155604 72858 155610 72860
rect 155769 72858 155835 72861
rect 155604 72856 155835 72858
rect 155604 72800 155774 72856
rect 155830 72800 155835 72856
rect 155604 72798 155835 72800
rect 155604 72796 155610 72798
rect 155769 72795 155835 72798
rect 156965 72858 157031 72861
rect 157190 72858 157196 72860
rect 156965 72856 157196 72858
rect 156965 72800 156970 72856
rect 157026 72800 157196 72856
rect 156965 72798 157196 72800
rect 156965 72795 157031 72798
rect 157190 72796 157196 72798
rect 157260 72796 157266 72860
rect 158294 72796 158300 72860
rect 158364 72858 158370 72860
rect 158621 72858 158687 72861
rect 158364 72856 158687 72858
rect 158364 72800 158626 72856
rect 158682 72800 158687 72856
rect 158364 72798 158687 72800
rect 158364 72796 158370 72798
rect 158621 72795 158687 72798
rect 158846 72796 158852 72860
rect 158916 72858 158922 72860
rect 159909 72858 159975 72861
rect 158916 72856 159975 72858
rect 158916 72800 159914 72856
rect 159970 72800 159975 72856
rect 158916 72798 159975 72800
rect 158916 72796 158922 72798
rect 159909 72795 159975 72798
rect 160686 72796 160692 72860
rect 160756 72858 160762 72860
rect 161197 72858 161263 72861
rect 160756 72856 161263 72858
rect 160756 72800 161202 72856
rect 161258 72800 161263 72856
rect 160756 72798 161263 72800
rect 160756 72796 160762 72798
rect 161197 72795 161263 72798
rect 162526 72796 162532 72860
rect 162596 72858 162602 72860
rect 162761 72858 162827 72861
rect 162596 72856 162827 72858
rect 162596 72800 162766 72856
rect 162822 72800 162827 72856
rect 162596 72798 162827 72800
rect 162596 72796 162602 72798
rect 162761 72795 162827 72798
rect 163262 72796 163268 72860
rect 163332 72858 163338 72860
rect 164049 72858 164115 72861
rect 163332 72856 164115 72858
rect 163332 72800 164054 72856
rect 164110 72800 164115 72856
rect 163332 72798 164115 72800
rect 163332 72796 163338 72798
rect 164049 72795 164115 72798
rect 165286 72796 165292 72860
rect 165356 72858 165362 72860
rect 165521 72858 165587 72861
rect 165356 72856 165587 72858
rect 165356 72800 165526 72856
rect 165582 72800 165587 72856
rect 165356 72798 165587 72800
rect 165662 72858 165722 72934
rect 167678 72932 167684 72934
rect 167748 72932 167754 72996
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 167862 72858 167868 72860
rect 165662 72798 167868 72858
rect 165356 72796 165362 72798
rect 165521 72795 165587 72798
rect 167862 72796 167868 72798
rect 167932 72796 167938 72860
rect 583520 72844 584960 72934
rect 148685 72722 148751 72725
rect 149973 72724 150039 72725
rect 148910 72722 148916 72724
rect 148685 72720 148916 72722
rect 148685 72664 148690 72720
rect 148746 72664 148916 72720
rect 148685 72662 148916 72664
rect 148685 72659 148751 72662
rect 148910 72660 148916 72662
rect 148980 72660 148986 72724
rect 149973 72720 150020 72724
rect 150084 72722 150090 72724
rect 151537 72722 151603 72725
rect 153009 72724 153075 72725
rect 151670 72722 151676 72724
rect 149973 72664 149978 72720
rect 149973 72660 150020 72664
rect 150084 72662 150130 72722
rect 151537 72720 151676 72722
rect 151537 72664 151542 72720
rect 151598 72664 151676 72720
rect 151537 72662 151676 72664
rect 150084 72660 150090 72662
rect 149973 72659 150039 72660
rect 151537 72659 151603 72662
rect 151670 72660 151676 72662
rect 151740 72660 151746 72724
rect 152958 72722 152964 72724
rect 152918 72662 152964 72722
rect 153028 72720 153075 72724
rect 153070 72664 153075 72720
rect 152958 72660 152964 72662
rect 153028 72660 153075 72664
rect 153009 72659 153075 72660
rect 154205 72724 154271 72725
rect 154205 72720 154252 72724
rect 154316 72722 154322 72724
rect 154205 72664 154210 72720
rect 154205 72660 154252 72664
rect 154316 72662 154362 72722
rect 154316 72660 154322 72662
rect 155718 72660 155724 72724
rect 155788 72722 155794 72724
rect 155861 72722 155927 72725
rect 156873 72724 156939 72725
rect 156822 72722 156828 72724
rect 155788 72720 155927 72722
rect 155788 72664 155866 72720
rect 155922 72664 155927 72720
rect 155788 72662 155927 72664
rect 156782 72662 156828 72722
rect 156892 72720 156939 72724
rect 156934 72664 156939 72720
rect 155788 72660 155794 72662
rect 154205 72659 154271 72660
rect 155861 72659 155927 72662
rect 156822 72660 156828 72662
rect 156892 72660 156939 72664
rect 157006 72660 157012 72724
rect 157076 72722 157082 72724
rect 157241 72722 157307 72725
rect 157076 72720 157307 72722
rect 157076 72664 157246 72720
rect 157302 72664 157307 72720
rect 157076 72662 157307 72664
rect 157076 72660 157082 72662
rect 156873 72659 156939 72660
rect 157241 72659 157307 72662
rect 158345 72722 158411 72725
rect 158478 72722 158484 72724
rect 158345 72720 158484 72722
rect 158345 72664 158350 72720
rect 158406 72664 158484 72720
rect 158345 72662 158484 72664
rect 158345 72659 158411 72662
rect 158478 72660 158484 72662
rect 158548 72660 158554 72724
rect 159030 72660 159036 72724
rect 159100 72722 159106 72724
rect 160001 72722 160067 72725
rect 159100 72720 160067 72722
rect 159100 72664 160006 72720
rect 160062 72664 160067 72720
rect 159100 72662 160067 72664
rect 159100 72660 159106 72662
rect 160001 72659 160067 72662
rect 160870 72660 160876 72724
rect 160940 72722 160946 72724
rect 161013 72722 161079 72725
rect 160940 72720 161079 72722
rect 160940 72664 161018 72720
rect 161074 72664 161079 72720
rect 160940 72662 161079 72664
rect 160940 72660 160946 72662
rect 161013 72659 161079 72662
rect 162485 72722 162551 72725
rect 162710 72722 162716 72724
rect 162485 72720 162716 72722
rect 162485 72664 162490 72720
rect 162546 72664 162716 72720
rect 162485 72662 162716 72664
rect 162485 72659 162551 72662
rect 162710 72660 162716 72662
rect 162780 72660 162786 72724
rect 163446 72660 163452 72724
rect 163516 72722 163522 72724
rect 163957 72722 164023 72725
rect 163516 72720 164023 72722
rect 163516 72664 163962 72720
rect 164018 72664 164023 72720
rect 163516 72662 164023 72664
rect 163516 72660 163522 72662
rect 163957 72659 164023 72662
rect 165102 72660 165108 72724
rect 165172 72722 165178 72724
rect 165245 72722 165311 72725
rect 165172 72720 165311 72722
rect 165172 72664 165250 72720
rect 165306 72664 165311 72720
rect 165172 72662 165311 72664
rect 165172 72660 165178 72662
rect 165245 72659 165311 72662
rect 166206 72660 166212 72724
rect 166276 72722 166282 72724
rect 166441 72722 166507 72725
rect 166809 72724 166875 72725
rect 166758 72722 166764 72724
rect 166276 72720 166507 72722
rect 166276 72664 166446 72720
rect 166502 72664 166507 72720
rect 166276 72662 166507 72664
rect 166718 72662 166764 72722
rect 166828 72720 166875 72724
rect 166870 72664 166875 72720
rect 166276 72660 166282 72662
rect 166441 72659 166507 72662
rect 166758 72660 166764 72662
rect 166828 72660 166875 72664
rect 166942 72660 166948 72724
rect 167012 72722 167018 72724
rect 404997 72722 405063 72725
rect 167012 72720 405063 72722
rect 167012 72664 405002 72720
rect 405058 72664 405063 72720
rect 167012 72662 405063 72664
rect 167012 72660 167018 72662
rect 166809 72659 166875 72660
rect 404997 72659 405063 72662
rect 22737 72586 22803 72589
rect 121913 72586 121979 72589
rect 22737 72584 121979 72586
rect 22737 72528 22742 72584
rect 22798 72528 121918 72584
rect 121974 72528 121979 72584
rect 22737 72526 121979 72528
rect 22737 72523 22803 72526
rect 121913 72523 121979 72526
rect 148358 72524 148364 72588
rect 148428 72586 148434 72588
rect 148869 72586 148935 72589
rect 148428 72584 148935 72586
rect 148428 72528 148874 72584
rect 148930 72528 148935 72584
rect 148428 72526 148935 72528
rect 148428 72524 148434 72526
rect 148869 72523 148935 72526
rect 149646 72524 149652 72588
rect 149716 72586 149722 72588
rect 150065 72586 150131 72589
rect 149716 72584 150131 72586
rect 149716 72528 150070 72584
rect 150126 72528 150131 72584
rect 149716 72526 150131 72528
rect 149716 72524 149722 72526
rect 150065 72523 150131 72526
rect 152406 72524 152412 72588
rect 152476 72586 152482 72588
rect 153101 72586 153167 72589
rect 152476 72584 153167 72586
rect 152476 72528 153106 72584
rect 153162 72528 153167 72584
rect 152476 72526 153167 72528
rect 152476 72524 152482 72526
rect 153101 72523 153167 72526
rect 154062 72524 154068 72588
rect 154132 72586 154138 72588
rect 154481 72586 154547 72589
rect 154132 72584 154547 72586
rect 154132 72528 154486 72584
rect 154542 72528 154547 72584
rect 154132 72526 154547 72528
rect 154132 72524 154138 72526
rect 154481 72523 154547 72526
rect 156638 72524 156644 72588
rect 156708 72586 156714 72588
rect 157057 72586 157123 72589
rect 156708 72584 157123 72586
rect 156708 72528 157062 72584
rect 157118 72528 157123 72584
rect 156708 72526 157123 72528
rect 156708 72524 156714 72526
rect 157057 72523 157123 72526
rect 158110 72524 158116 72588
rect 158180 72586 158186 72588
rect 158437 72586 158503 72589
rect 158180 72584 158503 72586
rect 158180 72528 158442 72584
rect 158498 72528 158503 72584
rect 158180 72526 158503 72528
rect 158180 72524 158186 72526
rect 158437 72523 158503 72526
rect 161054 72524 161060 72588
rect 161124 72586 161130 72588
rect 161381 72586 161447 72589
rect 161124 72584 161447 72586
rect 161124 72528 161386 72584
rect 161442 72528 161447 72584
rect 161124 72526 161447 72528
rect 161124 72524 161130 72526
rect 161381 72523 161447 72526
rect 162342 72524 162348 72588
rect 162412 72586 162418 72588
rect 162669 72586 162735 72589
rect 162412 72584 162735 72586
rect 162412 72528 162674 72584
rect 162730 72528 162735 72584
rect 162412 72526 162735 72528
rect 162412 72524 162418 72526
rect 162669 72523 162735 72526
rect 164918 72524 164924 72588
rect 164988 72586 164994 72588
rect 165429 72586 165495 72589
rect 164988 72584 165495 72586
rect 164988 72528 165434 72584
rect 165490 72528 165495 72584
rect 164988 72526 165495 72528
rect 164988 72524 164994 72526
rect 165429 72523 165495 72526
rect 166349 72586 166415 72589
rect 166574 72586 166580 72588
rect 166349 72584 166580 72586
rect 166349 72528 166354 72584
rect 166410 72528 166580 72584
rect 166349 72526 166580 72528
rect 166349 72523 166415 72526
rect 166574 72524 166580 72526
rect 166644 72524 166650 72588
rect 166809 72586 166875 72589
rect 480253 72586 480319 72589
rect 166809 72584 480319 72586
rect 166809 72528 166814 72584
rect 166870 72528 480258 72584
rect 480314 72528 480319 72584
rect 166809 72526 480319 72528
rect 166809 72523 166875 72526
rect 480253 72523 480319 72526
rect 148542 72388 148548 72452
rect 148612 72450 148618 72452
rect 148777 72450 148843 72453
rect 148612 72448 148843 72450
rect 148612 72392 148782 72448
rect 148838 72392 148843 72448
rect 148612 72390 148843 72392
rect 148612 72388 148618 72390
rect 148777 72387 148843 72390
rect 151302 72388 151308 72452
rect 151372 72450 151378 72452
rect 151629 72450 151695 72453
rect 151372 72448 151695 72450
rect 151372 72392 151634 72448
rect 151690 72392 151695 72448
rect 151372 72390 151695 72392
rect 151372 72388 151378 72390
rect 151629 72387 151695 72390
rect 152590 72388 152596 72452
rect 152660 72450 152666 72452
rect 152825 72450 152891 72453
rect 152660 72448 152891 72450
rect 152660 72392 152830 72448
rect 152886 72392 152891 72448
rect 152660 72390 152891 72392
rect 152660 72388 152666 72390
rect 152825 72387 152891 72390
rect 155677 72450 155743 72453
rect 157057 72450 157123 72453
rect 155677 72448 157123 72450
rect 155677 72392 155682 72448
rect 155738 72392 157062 72448
rect 157118 72392 157123 72448
rect 155677 72390 157123 72392
rect 155677 72387 155743 72390
rect 157057 72387 157123 72390
rect 158529 72450 158595 72453
rect 158662 72450 158668 72452
rect 158529 72448 158668 72450
rect 158529 72392 158534 72448
rect 158590 72392 158668 72448
rect 158529 72390 158668 72392
rect 158529 72387 158595 72390
rect 158662 72388 158668 72390
rect 158732 72388 158738 72452
rect 161105 72450 161171 72453
rect 161238 72450 161244 72452
rect 161105 72448 161244 72450
rect 161105 72392 161110 72448
rect 161166 72392 161244 72448
rect 161105 72390 161244 72392
rect 161105 72387 161171 72390
rect 161238 72388 161244 72390
rect 161308 72388 161314 72452
rect 162761 72450 162827 72453
rect 162894 72450 162900 72452
rect 162761 72448 162900 72450
rect 162761 72392 162766 72448
rect 162822 72392 162900 72448
rect 162761 72390 162900 72392
rect 162761 72387 162827 72390
rect 162894 72388 162900 72390
rect 162964 72388 162970 72452
rect 163630 72388 163636 72452
rect 163700 72450 163706 72452
rect 164141 72450 164207 72453
rect 163700 72448 164207 72450
rect 163700 72392 164146 72448
rect 164202 72392 164207 72448
rect 163700 72390 164207 72392
rect 163700 72388 163706 72390
rect 164141 72387 164207 72390
rect 165337 72450 165403 72453
rect 165470 72450 165476 72452
rect 165337 72448 165476 72450
rect 165337 72392 165342 72448
rect 165398 72392 165476 72448
rect 165337 72390 165476 72392
rect 165337 72387 165403 72390
rect 165470 72388 165476 72390
rect 165540 72388 165546 72452
rect 166390 72388 166396 72452
rect 166460 72450 166466 72452
rect 166533 72450 166599 72453
rect 498193 72450 498259 72453
rect 166460 72448 166599 72450
rect 166460 72392 166538 72448
rect 166594 72392 166599 72448
rect 166460 72390 166599 72392
rect 166460 72388 166466 72390
rect 166533 72387 166599 72390
rect 166950 72448 498259 72450
rect 166950 72392 498198 72448
rect 498254 72392 498259 72448
rect 166950 72390 498259 72392
rect 125685 72314 125751 72317
rect 126094 72314 126100 72316
rect 125685 72312 126100 72314
rect 125685 72256 125690 72312
rect 125746 72256 126100 72312
rect 125685 72254 126100 72256
rect 125685 72251 125751 72254
rect 126094 72252 126100 72254
rect 126164 72252 126170 72316
rect 142838 72252 142844 72316
rect 142908 72314 142914 72316
rect 143257 72314 143323 72317
rect 142908 72312 143323 72314
rect 142908 72256 143262 72312
rect 143318 72256 143323 72312
rect 142908 72254 143323 72256
rect 142908 72252 142914 72254
rect 143257 72251 143323 72254
rect 159633 72314 159699 72317
rect 161013 72314 161079 72317
rect 159633 72312 161079 72314
rect 159633 72256 159638 72312
rect 159694 72256 161018 72312
rect 161074 72256 161079 72312
rect 159633 72254 161079 72256
rect 159633 72251 159699 72254
rect 161013 72251 161079 72254
rect 124213 72178 124279 72181
rect 124622 72178 124628 72180
rect 124213 72176 124628 72178
rect 124213 72120 124218 72176
rect 124274 72120 124628 72176
rect 124213 72118 124628 72120
rect 124213 72115 124279 72118
rect 124622 72116 124628 72118
rect 124692 72116 124698 72180
rect 125542 72116 125548 72180
rect 125612 72178 125618 72180
rect 125777 72178 125843 72181
rect 125612 72176 125843 72178
rect 125612 72120 125782 72176
rect 125838 72120 125843 72176
rect 125612 72118 125843 72120
rect 125612 72116 125618 72118
rect 125777 72115 125843 72118
rect 128445 72178 128511 72181
rect 129038 72178 129044 72180
rect 128445 72176 129044 72178
rect 128445 72120 128450 72176
rect 128506 72120 129044 72176
rect 128445 72118 129044 72120
rect 128445 72115 128511 72118
rect 129038 72116 129044 72118
rect 129108 72116 129114 72180
rect 129733 72178 129799 72181
rect 129958 72178 129964 72180
rect 129733 72176 129964 72178
rect 129733 72120 129738 72176
rect 129794 72120 129964 72176
rect 129733 72118 129964 72120
rect 129733 72115 129799 72118
rect 129958 72116 129964 72118
rect 130028 72116 130034 72180
rect 133270 72116 133276 72180
rect 133340 72178 133346 72180
rect 133597 72178 133663 72181
rect 133340 72176 133663 72178
rect 133340 72120 133602 72176
rect 133658 72120 133663 72176
rect 133340 72118 133663 72120
rect 133340 72116 133346 72118
rect 133597 72115 133663 72118
rect 134742 72116 134748 72180
rect 134812 72178 134818 72180
rect 135069 72178 135135 72181
rect 134812 72176 135135 72178
rect 134812 72120 135074 72176
rect 135130 72120 135135 72176
rect 134812 72118 135135 72120
rect 134812 72116 134818 72118
rect 135069 72115 135135 72118
rect 136030 72116 136036 72180
rect 136100 72178 136106 72180
rect 136449 72178 136515 72181
rect 136100 72176 136515 72178
rect 136100 72120 136454 72176
rect 136510 72120 136515 72176
rect 136100 72118 136515 72120
rect 136100 72116 136106 72118
rect 136449 72115 136515 72118
rect 138974 72116 138980 72180
rect 139044 72178 139050 72180
rect 139301 72178 139367 72181
rect 139044 72176 139367 72178
rect 139044 72120 139306 72176
rect 139362 72120 139367 72176
rect 139044 72118 139367 72120
rect 139044 72116 139050 72118
rect 139301 72115 139367 72118
rect 140078 72116 140084 72180
rect 140148 72178 140154 72180
rect 140313 72178 140379 72181
rect 140148 72176 140379 72178
rect 140148 72120 140318 72176
rect 140374 72120 140379 72176
rect 140148 72118 140379 72120
rect 140148 72116 140154 72118
rect 140313 72115 140379 72118
rect 143022 72116 143028 72180
rect 143092 72178 143098 72180
rect 143349 72178 143415 72181
rect 143092 72176 143415 72178
rect 143092 72120 143354 72176
rect 143410 72120 143415 72176
rect 143092 72118 143415 72120
rect 143092 72116 143098 72118
rect 143349 72115 143415 72118
rect 144126 72116 144132 72180
rect 144196 72178 144202 72180
rect 144729 72178 144795 72181
rect 144196 72176 144795 72178
rect 144196 72120 144734 72176
rect 144790 72120 144795 72176
rect 144196 72118 144795 72120
rect 144196 72116 144202 72118
rect 144729 72115 144795 72118
rect 145230 72116 145236 72180
rect 145300 72178 145306 72180
rect 146017 72178 146083 72181
rect 145300 72176 146083 72178
rect 145300 72120 146022 72176
rect 146078 72120 146083 72176
rect 145300 72118 146083 72120
rect 145300 72116 145306 72118
rect 146017 72115 146083 72118
rect 146886 72116 146892 72180
rect 146956 72178 146962 72180
rect 147489 72178 147555 72181
rect 146956 72176 147555 72178
rect 146956 72120 147494 72176
rect 147550 72120 147555 72176
rect 146956 72118 147555 72120
rect 146956 72116 146962 72118
rect 147489 72115 147555 72118
rect 157149 72178 157215 72181
rect 157793 72178 157859 72181
rect 157149 72176 157859 72178
rect 157149 72120 157154 72176
rect 157210 72120 157798 72176
rect 157854 72120 157859 72176
rect 157149 72118 157859 72120
rect 157149 72115 157215 72118
rect 157793 72115 157859 72118
rect 160277 72178 160343 72181
rect 166950 72178 167010 72390
rect 498193 72387 498259 72390
rect 160277 72176 167010 72178
rect 160277 72120 160282 72176
rect 160338 72120 167010 72176
rect 160277 72118 167010 72120
rect 160277 72115 160343 72118
rect 121637 72044 121703 72045
rect 122833 72044 122899 72045
rect 121637 72042 121684 72044
rect 121592 72040 121684 72042
rect 121592 71984 121642 72040
rect 121592 71982 121684 71984
rect 121637 71980 121684 71982
rect 121748 71980 121754 72044
rect 122782 71980 122788 72044
rect 122852 72042 122899 72044
rect 122852 72040 122944 72042
rect 122894 71984 122944 72040
rect 122852 71982 122944 71984
rect 122852 71980 122899 71982
rect 124254 71980 124260 72044
rect 124324 72042 124330 72044
rect 124397 72042 124463 72045
rect 124324 72040 124463 72042
rect 124324 71984 124402 72040
rect 124458 71984 124463 72040
rect 124324 71982 124463 71984
rect 124324 71980 124330 71982
rect 121637 71979 121703 71980
rect 122833 71979 122899 71980
rect 124397 71979 124463 71982
rect 125593 72042 125659 72045
rect 125726 72042 125732 72044
rect 125593 72040 125732 72042
rect 125593 71984 125598 72040
rect 125654 71984 125732 72040
rect 125593 71982 125732 71984
rect 125593 71979 125659 71982
rect 125726 71980 125732 71982
rect 125796 71980 125802 72044
rect 127065 72042 127131 72045
rect 127198 72042 127204 72044
rect 127065 72040 127204 72042
rect 127065 71984 127070 72040
rect 127126 71984 127204 72040
rect 127065 71982 127204 71984
rect 127065 71979 127131 71982
rect 127198 71980 127204 71982
rect 127268 71980 127274 72044
rect 128353 72042 128419 72045
rect 128854 72042 128860 72044
rect 128353 72040 128860 72042
rect 128353 71984 128358 72040
rect 128414 71984 128860 72040
rect 128353 71982 128860 71984
rect 128353 71979 128419 71982
rect 128854 71980 128860 71982
rect 128924 71980 128930 72044
rect 130009 72042 130075 72045
rect 131205 72044 131271 72045
rect 130142 72042 130148 72044
rect 130009 72040 130148 72042
rect 130009 71984 130014 72040
rect 130070 71984 130148 72040
rect 130009 71982 130148 71984
rect 130009 71979 130075 71982
rect 130142 71980 130148 71982
rect 130212 71980 130218 72044
rect 131205 72042 131252 72044
rect 131160 72040 131252 72042
rect 131160 71984 131210 72040
rect 131160 71982 131252 71984
rect 131205 71980 131252 71982
rect 131316 71980 131322 72044
rect 131798 71980 131804 72044
rect 131868 72042 131874 72044
rect 132217 72042 132283 72045
rect 131868 72040 132283 72042
rect 131868 71984 132222 72040
rect 132278 71984 132283 72040
rect 131868 71982 132283 71984
rect 131868 71980 131874 71982
rect 131205 71979 131271 71980
rect 132217 71979 132283 71982
rect 133454 71980 133460 72044
rect 133524 72042 133530 72044
rect 133689 72042 133755 72045
rect 134977 72044 135043 72045
rect 134926 72042 134932 72044
rect 133524 72040 133755 72042
rect 133524 71984 133694 72040
rect 133750 71984 133755 72040
rect 133524 71982 133755 71984
rect 134886 71982 134932 72042
rect 134996 72040 135043 72044
rect 135038 71984 135043 72040
rect 133524 71980 133530 71982
rect 133689 71979 133755 71982
rect 134926 71980 134932 71982
rect 134996 71980 135043 71984
rect 136214 71980 136220 72044
rect 136284 72042 136290 72044
rect 136357 72042 136423 72045
rect 136284 72040 136423 72042
rect 136284 71984 136362 72040
rect 136418 71984 136423 72040
rect 136284 71982 136423 71984
rect 136284 71980 136290 71982
rect 134977 71979 135043 71980
rect 136357 71979 136423 71982
rect 137686 71980 137692 72044
rect 137756 72042 137762 72044
rect 137829 72042 137895 72045
rect 137756 72040 137895 72042
rect 137756 71984 137834 72040
rect 137890 71984 137895 72040
rect 137756 71982 137895 71984
rect 137756 71980 137762 71982
rect 137829 71979 137895 71982
rect 138790 71980 138796 72044
rect 138860 72042 138866 72044
rect 139025 72042 139091 72045
rect 138860 72040 139091 72042
rect 138860 71984 139030 72040
rect 139086 71984 139091 72040
rect 138860 71982 139091 71984
rect 138860 71980 138866 71982
rect 139025 71979 139091 71982
rect 140262 71980 140268 72044
rect 140332 72042 140338 72044
rect 140589 72042 140655 72045
rect 140332 72040 140655 72042
rect 140332 71984 140594 72040
rect 140650 71984 140655 72040
rect 140332 71982 140655 71984
rect 140332 71980 140338 71982
rect 140589 71979 140655 71982
rect 140814 71980 140820 72044
rect 140884 72042 140890 72044
rect 141969 72042 142035 72045
rect 140884 72040 142035 72042
rect 140884 71984 141974 72040
rect 142030 71984 142035 72040
rect 140884 71982 142035 71984
rect 140884 71980 140890 71982
rect 141969 71979 142035 71982
rect 143206 71980 143212 72044
rect 143276 72042 143282 72044
rect 143441 72042 143507 72045
rect 143276 72040 143507 72042
rect 143276 71984 143446 72040
rect 143502 71984 143507 72040
rect 143276 71982 143507 71984
rect 143276 71980 143282 71982
rect 143441 71979 143507 71982
rect 144494 71980 144500 72044
rect 144564 72042 144570 72044
rect 144637 72042 144703 72045
rect 144564 72040 144703 72042
rect 144564 71984 144642 72040
rect 144698 71984 144703 72040
rect 144564 71982 144703 71984
rect 144564 71980 144570 71982
rect 144637 71979 144703 71982
rect 145414 71980 145420 72044
rect 145484 72042 145490 72044
rect 146201 72042 146267 72045
rect 145484 72040 146267 72042
rect 145484 71984 146206 72040
rect 146262 71984 146267 72040
rect 145484 71982 146267 71984
rect 145484 71980 145490 71982
rect 146201 71979 146267 71982
rect 147070 71980 147076 72044
rect 147140 72042 147146 72044
rect 147397 72042 147463 72045
rect 147140 72040 147463 72042
rect 147140 71984 147402 72040
rect 147458 71984 147463 72040
rect 147140 71982 147463 71984
rect 147140 71980 147146 71982
rect 147397 71979 147463 71982
rect 158897 72042 158963 72045
rect 166809 72042 166875 72045
rect 158897 72040 166875 72042
rect 158897 71984 158902 72040
rect 158958 71984 166814 72040
rect 166870 71984 166875 72040
rect 158897 71982 166875 71984
rect 158897 71979 158963 71982
rect 166809 71979 166875 71982
rect 121545 71908 121611 71909
rect 121494 71906 121500 71908
rect 121454 71846 121500 71906
rect 121564 71904 121611 71908
rect 122925 71908 122991 71909
rect 124489 71908 124555 71909
rect 122925 71906 122972 71908
rect 121606 71848 121611 71904
rect 121494 71844 121500 71846
rect 121564 71844 121611 71848
rect 122880 71904 122972 71906
rect 122880 71848 122930 71904
rect 122880 71846 122972 71848
rect 121545 71843 121611 71844
rect 122925 71844 122972 71846
rect 123036 71844 123042 71908
rect 124438 71906 124444 71908
rect 124398 71846 124444 71906
rect 124508 71904 124555 71908
rect 125869 71908 125935 71909
rect 126973 71908 127039 71909
rect 128629 71908 128695 71909
rect 125869 71906 125916 71908
rect 124550 71848 124555 71904
rect 124438 71844 124444 71846
rect 124508 71844 124555 71848
rect 125824 71904 125916 71906
rect 125824 71848 125874 71904
rect 125824 71846 125916 71848
rect 122925 71843 122991 71844
rect 124489 71843 124555 71844
rect 125869 71844 125916 71846
rect 125980 71844 125986 71908
rect 126973 71906 127020 71908
rect 126928 71904 127020 71906
rect 126928 71848 126978 71904
rect 126928 71846 127020 71848
rect 126973 71844 127020 71846
rect 127084 71844 127090 71908
rect 128629 71906 128676 71908
rect 128584 71904 128676 71906
rect 128584 71848 128634 71904
rect 128584 71846 128676 71848
rect 128629 71844 128676 71846
rect 128740 71844 128746 71908
rect 129774 71844 129780 71908
rect 129844 71906 129850 71908
rect 129917 71906 129983 71909
rect 131113 71908 131179 71909
rect 131062 71906 131068 71908
rect 129844 71904 129983 71906
rect 129844 71848 129922 71904
rect 129978 71848 129983 71904
rect 129844 71846 129983 71848
rect 131022 71846 131068 71906
rect 131132 71904 131179 71908
rect 131174 71848 131179 71904
rect 129844 71844 129850 71846
rect 125869 71843 125935 71844
rect 126973 71843 127039 71844
rect 128629 71843 128695 71844
rect 129917 71843 129983 71846
rect 131062 71844 131068 71846
rect 131132 71844 131179 71848
rect 131982 71844 131988 71908
rect 132052 71906 132058 71908
rect 132401 71906 132467 71909
rect 132052 71904 132467 71906
rect 132052 71848 132406 71904
rect 132462 71848 132467 71904
rect 132052 71846 132467 71848
rect 132052 71844 132058 71846
rect 131113 71843 131179 71844
rect 132401 71843 132467 71846
rect 133638 71844 133644 71908
rect 133708 71906 133714 71908
rect 133781 71906 133847 71909
rect 135161 71908 135227 71909
rect 135110 71906 135116 71908
rect 133708 71904 133847 71906
rect 133708 71848 133786 71904
rect 133842 71848 133847 71904
rect 133708 71846 133847 71848
rect 135070 71846 135116 71906
rect 135180 71904 135227 71908
rect 135222 71848 135227 71904
rect 133708 71844 133714 71846
rect 133781 71843 133847 71846
rect 135110 71844 135116 71846
rect 135180 71844 135227 71848
rect 135846 71844 135852 71908
rect 135916 71906 135922 71908
rect 136173 71906 136239 71909
rect 135916 71904 136239 71906
rect 135916 71848 136178 71904
rect 136234 71848 136239 71904
rect 135916 71846 136239 71848
rect 135916 71844 135922 71846
rect 135161 71843 135227 71844
rect 136173 71843 136239 71846
rect 136398 71844 136404 71908
rect 136468 71906 136474 71908
rect 136541 71906 136607 71909
rect 137921 71908 137987 71909
rect 137870 71906 137876 71908
rect 136468 71904 136607 71906
rect 136468 71848 136546 71904
rect 136602 71848 136607 71904
rect 136468 71846 136607 71848
rect 137830 71846 137876 71906
rect 137940 71904 137987 71908
rect 137982 71848 137987 71904
rect 136468 71844 136474 71846
rect 136541 71843 136607 71846
rect 137870 71844 137876 71846
rect 137940 71844 137987 71848
rect 138606 71844 138612 71908
rect 138676 71906 138682 71908
rect 138933 71906 138999 71909
rect 139117 71908 139183 71909
rect 140405 71908 140471 71909
rect 140681 71908 140747 71909
rect 139117 71906 139164 71908
rect 138676 71904 138999 71906
rect 138676 71848 138938 71904
rect 138994 71848 138999 71904
rect 138676 71846 138999 71848
rect 139072 71904 139164 71906
rect 139072 71848 139122 71904
rect 139072 71846 139164 71848
rect 138676 71844 138682 71846
rect 137921 71843 137987 71844
rect 138933 71843 138999 71846
rect 139117 71844 139164 71846
rect 139228 71844 139234 71908
rect 140405 71906 140452 71908
rect 140360 71904 140452 71906
rect 140360 71848 140410 71904
rect 140360 71846 140452 71848
rect 140405 71844 140452 71846
rect 140516 71844 140522 71908
rect 140630 71844 140636 71908
rect 140700 71906 140747 71908
rect 140700 71904 140792 71906
rect 140742 71848 140792 71904
rect 140700 71846 140792 71848
rect 140700 71844 140747 71846
rect 140998 71844 141004 71908
rect 141068 71906 141074 71908
rect 142061 71906 142127 71909
rect 141068 71904 142127 71906
rect 141068 71848 142066 71904
rect 142122 71848 142127 71904
rect 141068 71846 142127 71848
rect 141068 71844 141074 71846
rect 139117 71843 139183 71844
rect 140405 71843 140471 71844
rect 140681 71843 140747 71844
rect 142061 71843 142127 71846
rect 143165 71906 143231 71909
rect 143390 71906 143396 71908
rect 143165 71904 143396 71906
rect 143165 71848 143170 71904
rect 143226 71848 143396 71904
rect 143165 71846 143396 71848
rect 143165 71843 143231 71846
rect 143390 71844 143396 71846
rect 143460 71844 143466 71908
rect 144310 71844 144316 71908
rect 144380 71906 144386 71908
rect 144545 71906 144611 71909
rect 144380 71904 144611 71906
rect 144380 71848 144550 71904
rect 144606 71848 144611 71904
rect 144380 71846 144611 71848
rect 144380 71844 144386 71846
rect 144545 71843 144611 71846
rect 144678 71844 144684 71908
rect 144748 71906 144754 71908
rect 144821 71906 144887 71909
rect 144748 71904 144887 71906
rect 144748 71848 144826 71904
rect 144882 71848 144887 71904
rect 144748 71846 144887 71848
rect 144748 71844 144754 71846
rect 144821 71843 144887 71846
rect 145598 71844 145604 71908
rect 145668 71906 145674 71908
rect 146109 71906 146175 71909
rect 147305 71908 147371 71909
rect 147254 71906 147260 71908
rect 145668 71904 146175 71906
rect 145668 71848 146114 71904
rect 146170 71848 146175 71904
rect 145668 71846 146175 71848
rect 147214 71846 147260 71906
rect 147324 71904 147371 71908
rect 147366 71848 147371 71904
rect 145668 71844 145674 71846
rect 146109 71843 146175 71846
rect 147254 71844 147260 71846
rect 147324 71844 147371 71848
rect 147438 71844 147444 71908
rect 147508 71906 147514 71908
rect 147581 71906 147647 71909
rect 147508 71904 147647 71906
rect 147508 71848 147586 71904
rect 147642 71848 147647 71904
rect 147508 71846 147647 71848
rect 147508 71844 147514 71846
rect 147305 71843 147371 71844
rect 147581 71843 147647 71846
rect 158805 71906 158871 71909
rect 166942 71906 166948 71908
rect 158805 71904 166948 71906
rect 158805 71848 158810 71904
rect 158866 71848 166948 71904
rect 158805 71846 166948 71848
rect 158805 71843 158871 71846
rect 166942 71844 166948 71846
rect 167012 71844 167018 71908
rect -960 71634 480 71724
rect 3509 71634 3575 71637
rect -960 71632 3575 71634
rect -960 71576 3514 71632
rect 3570 71576 3575 71632
rect -960 71574 3575 71576
rect -960 71484 480 71574
rect 3509 71571 3575 71574
rect 158662 65452 158668 65516
rect 158732 65514 158738 65516
rect 474733 65514 474799 65517
rect 158732 65512 474799 65514
rect 158732 65456 474738 65512
rect 474794 65456 474799 65512
rect 158732 65454 474799 65456
rect 158732 65452 158738 65454
rect 474733 65451 474799 65454
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3601 58578 3667 58581
rect -960 58576 3667 58578
rect -960 58520 3606 58576
rect 3662 58520 3667 58576
rect -960 58518 3667 58520
rect -960 58428 480 58518
rect 3601 58515 3667 58518
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3509 45522 3575 45525
rect -960 45520 3575 45522
rect -960 45464 3514 45520
rect 3570 45464 3575 45520
rect -960 45462 3575 45464
rect -960 45372 480 45462
rect 3509 45459 3575 45462
rect 144126 35260 144132 35324
rect 144196 35322 144202 35324
rect 298093 35322 298159 35325
rect 144196 35320 298159 35322
rect 144196 35264 298098 35320
rect 298154 35264 298159 35320
rect 144196 35262 298159 35264
rect 144196 35260 144202 35262
rect 298093 35259 298159 35262
rect 146886 35124 146892 35188
rect 146956 35186 146962 35188
rect 332593 35186 332659 35189
rect 146956 35184 332659 35186
rect 146956 35128 332598 35184
rect 332654 35128 332659 35184
rect 146956 35126 332659 35128
rect 146956 35124 146962 35126
rect 332593 35123 332659 35126
rect 137686 34036 137692 34100
rect 137756 34098 137762 34100
rect 209773 34098 209839 34101
rect 137756 34096 209839 34098
rect 137756 34040 209778 34096
rect 209834 34040 209839 34096
rect 137756 34038 209839 34040
rect 137756 34036 137762 34038
rect 209773 34035 209839 34038
rect 140078 33900 140084 33964
rect 140148 33962 140154 33964
rect 241513 33962 241579 33965
rect 140148 33960 241579 33962
rect 140148 33904 241518 33960
rect 241574 33904 241579 33960
rect 140148 33902 241579 33904
rect 140148 33900 140154 33902
rect 241513 33899 241579 33902
rect 140814 33764 140820 33828
rect 140884 33826 140890 33828
rect 262213 33826 262279 33829
rect 140884 33824 262279 33826
rect 140884 33768 262218 33824
rect 262274 33768 262279 33824
rect 140884 33766 262279 33768
rect 140884 33764 140890 33766
rect 262213 33763 262279 33766
rect 580257 33146 580323 33149
rect 583520 33146 584960 33236
rect 580257 33144 584960 33146
rect 580257 33088 580262 33144
rect 580318 33088 584960 33144
rect 580257 33086 584960 33088
rect 580257 33083 580323 33086
rect 583520 32996 584960 33086
rect 134742 32676 134748 32740
rect 134812 32738 134818 32740
rect 173893 32738 173959 32741
rect 134812 32736 173959 32738
rect 134812 32680 173898 32736
rect 173954 32680 173959 32736
rect 134812 32678 173959 32680
rect 134812 32676 134818 32678
rect 173893 32675 173959 32678
rect -960 32466 480 32556
rect 135846 32540 135852 32604
rect 135916 32602 135922 32604
rect 187693 32602 187759 32605
rect 135916 32600 187759 32602
rect 135916 32544 187698 32600
rect 187754 32544 187759 32600
rect 135916 32542 187759 32544
rect 135916 32540 135922 32542
rect 187693 32539 187759 32542
rect 2865 32466 2931 32469
rect -960 32464 2931 32466
rect -960 32408 2870 32464
rect 2926 32408 2931 32464
rect -960 32406 2931 32408
rect -960 32316 480 32406
rect 2865 32403 2931 32406
rect 136030 32404 136036 32468
rect 136100 32466 136106 32468
rect 191833 32466 191899 32469
rect 136100 32464 191899 32466
rect 136100 32408 191838 32464
rect 191894 32408 191899 32464
rect 136100 32406 191899 32408
rect 136100 32404 136106 32406
rect 191833 32403 191899 32406
rect 166206 31724 166212 31788
rect 166276 31786 166282 31788
rect 166901 31786 166967 31789
rect 166276 31784 166967 31786
rect 166276 31728 166906 31784
rect 166962 31728 166967 31784
rect 166276 31726 166967 31728
rect 166276 31724 166282 31726
rect 166901 31723 166967 31726
rect 163262 31180 163268 31244
rect 163332 31242 163338 31244
rect 445017 31242 445083 31245
rect 163332 31240 445083 31242
rect 163332 31184 445022 31240
rect 445078 31184 445083 31240
rect 163332 31182 445083 31184
rect 163332 31180 163338 31182
rect 445017 31179 445083 31182
rect 158110 31044 158116 31108
rect 158180 31106 158186 31108
rect 473353 31106 473419 31109
rect 158180 31104 473419 31106
rect 158180 31048 473358 31104
rect 473414 31048 473419 31104
rect 158180 31046 473419 31048
rect 158180 31044 158186 31046
rect 473353 31043 473419 31046
rect 158846 30908 158852 30972
rect 158916 30970 158922 30972
rect 492673 30970 492739 30973
rect 158916 30968 492739 30970
rect 158916 30912 492678 30968
rect 492734 30912 492739 30968
rect 158916 30910 492739 30912
rect 158916 30908 158922 30910
rect 492673 30907 492739 30910
rect 145230 29548 145236 29612
rect 145300 29610 145306 29612
rect 314653 29610 314719 29613
rect 145300 29608 314719 29610
rect 145300 29552 314658 29608
rect 314714 29552 314719 29608
rect 145300 29550 314719 29552
rect 145300 29548 145306 29550
rect 314653 29547 314719 29550
rect 136214 27100 136220 27164
rect 136284 27162 136290 27164
rect 190453 27162 190519 27165
rect 136284 27160 190519 27162
rect 136284 27104 190458 27160
rect 190514 27104 190519 27160
rect 136284 27102 190519 27104
rect 136284 27100 136290 27102
rect 190453 27099 190519 27102
rect 142838 26964 142844 27028
rect 142908 27026 142914 27028
rect 278773 27026 278839 27029
rect 142908 27024 278839 27026
rect 142908 26968 278778 27024
rect 278834 26968 278839 27024
rect 142908 26966 278839 26968
rect 142908 26964 142914 26966
rect 278773 26963 278839 26966
rect 149462 26828 149468 26892
rect 149532 26890 149538 26892
rect 367093 26890 367159 26893
rect 149532 26888 367159 26890
rect 149532 26832 367098 26888
rect 367154 26832 367159 26888
rect 149532 26830 367159 26832
rect 149532 26828 149538 26830
rect 367093 26827 367159 26830
rect 134926 25604 134932 25668
rect 134996 25666 135002 25668
rect 172513 25666 172579 25669
rect 134996 25664 172579 25666
rect 134996 25608 172518 25664
rect 172574 25608 172579 25664
rect 134996 25606 172579 25608
rect 134996 25604 135002 25606
rect 172513 25603 172579 25606
rect 156638 25468 156644 25532
rect 156708 25530 156714 25532
rect 456885 25530 456951 25533
rect 156708 25528 456951 25530
rect 156708 25472 456890 25528
rect 456946 25472 456951 25528
rect 156708 25470 456951 25472
rect 156708 25468 156714 25470
rect 456885 25467 456951 25470
rect 151302 24380 151308 24444
rect 151372 24442 151378 24444
rect 386413 24442 386479 24445
rect 151372 24440 386479 24442
rect 151372 24384 386418 24440
rect 386474 24384 386479 24440
rect 151372 24382 386479 24384
rect 151372 24380 151378 24382
rect 386413 24379 386479 24382
rect 162158 24244 162164 24308
rect 162228 24306 162234 24308
rect 527173 24306 527239 24309
rect 162228 24304 527239 24306
rect 162228 24248 527178 24304
rect 527234 24248 527239 24304
rect 162228 24246 527239 24248
rect 162228 24244 162234 24246
rect 527173 24243 527239 24246
rect 163446 24108 163452 24172
rect 163516 24170 163522 24172
rect 545113 24170 545179 24173
rect 163516 24168 545179 24170
rect 163516 24112 545118 24168
rect 545174 24112 545179 24168
rect 163516 24110 545179 24112
rect 163516 24108 163522 24110
rect 545113 24107 545179 24110
rect 156822 22748 156828 22812
rect 156892 22810 156898 22812
rect 454033 22810 454099 22813
rect 156892 22808 454099 22810
rect 156892 22752 454038 22808
rect 454094 22752 454099 22808
rect 156892 22750 454099 22752
rect 156892 22748 156898 22750
rect 454033 22747 454099 22750
rect 160686 22612 160692 22676
rect 160756 22674 160762 22676
rect 509233 22674 509299 22677
rect 160756 22672 509299 22674
rect 160756 22616 509238 22672
rect 509294 22616 509299 22672
rect 160756 22614 509299 22616
rect 160756 22612 160762 22614
rect 509233 22611 509299 22614
rect 148358 21524 148364 21588
rect 148428 21586 148434 21588
rect 350533 21586 350599 21589
rect 148428 21584 350599 21586
rect 148428 21528 350538 21584
rect 350594 21528 350599 21584
rect 148428 21526 350599 21528
rect 148428 21524 148434 21526
rect 350533 21523 350599 21526
rect 155534 21388 155540 21452
rect 155604 21450 155610 21452
rect 440233 21450 440299 21453
rect 155604 21448 440299 21450
rect 155604 21392 440238 21448
rect 440294 21392 440299 21448
rect 155604 21390 440299 21392
rect 155604 21388 155610 21390
rect 440233 21387 440299 21390
rect 158294 21252 158300 21316
rect 158364 21314 158370 21316
rect 476113 21314 476179 21317
rect 158364 21312 476179 21314
rect 158364 21256 476118 21312
rect 476174 21256 476179 21312
rect 158364 21254 476179 21256
rect 158364 21252 158370 21254
rect 476113 21251 476179 21254
rect 138606 20164 138612 20228
rect 138676 20226 138682 20228
rect 223573 20226 223639 20229
rect 138676 20224 223639 20226
rect 138676 20168 223578 20224
rect 223634 20168 223639 20224
rect 138676 20166 223639 20168
rect 138676 20164 138682 20166
rect 223573 20163 223639 20166
rect 140262 20028 140268 20092
rect 140332 20090 140338 20092
rect 244273 20090 244339 20093
rect 140332 20088 244339 20090
rect 140332 20032 244278 20088
rect 244334 20032 244339 20088
rect 140332 20030 244339 20032
rect 140332 20028 140338 20030
rect 244273 20027 244339 20030
rect 158478 19892 158484 19956
rect 158548 19954 158554 19956
rect 473445 19954 473511 19957
rect 158548 19952 473511 19954
rect 158548 19896 473450 19952
rect 473506 19896 473511 19952
rect 158548 19894 473511 19896
rect 158548 19892 158554 19894
rect 473445 19891 473511 19894
rect 580165 19818 580231 19821
rect 583520 19818 584960 19908
rect 580165 19816 584960 19818
rect 580165 19760 580170 19816
rect 580226 19760 584960 19816
rect 580165 19758 584960 19760
rect 580165 19755 580231 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 157190 18804 157196 18868
rect 157260 18866 157266 18868
rect 455413 18866 455479 18869
rect 157260 18864 455479 18866
rect 157260 18808 455418 18864
rect 455474 18808 455479 18864
rect 157260 18806 455479 18808
rect 157260 18804 157266 18806
rect 455413 18803 455479 18806
rect 157006 18668 157012 18732
rect 157076 18730 157082 18732
rect 458173 18730 458239 18733
rect 157076 18728 458239 18730
rect 157076 18672 458178 18728
rect 458234 18672 458239 18728
rect 157076 18670 458239 18672
rect 157076 18668 157082 18670
rect 458173 18667 458239 18670
rect 162342 18532 162348 18596
rect 162412 18594 162418 18596
rect 528553 18594 528619 18597
rect 162412 18592 528619 18594
rect 162412 18536 528558 18592
rect 528614 18536 528619 18592
rect 162412 18534 528619 18536
rect 162412 18532 162418 18534
rect 528553 18531 528619 18534
rect 145414 17580 145420 17644
rect 145484 17642 145490 17644
rect 316033 17642 316099 17645
rect 145484 17640 316099 17642
rect 145484 17584 316038 17640
rect 316094 17584 316099 17640
rect 145484 17582 316099 17584
rect 145484 17580 145490 17582
rect 316033 17579 316099 17582
rect 153878 17444 153884 17508
rect 153948 17506 153954 17508
rect 420913 17506 420979 17509
rect 153948 17504 420979 17506
rect 153948 17448 420918 17504
rect 420974 17448 420979 17504
rect 153948 17446 420979 17448
rect 153948 17444 153954 17446
rect 420913 17443 420979 17446
rect 154062 17308 154068 17372
rect 154132 17370 154138 17372
rect 423765 17370 423831 17373
rect 154132 17368 423831 17370
rect 154132 17312 423770 17368
rect 423826 17312 423831 17368
rect 154132 17310 423831 17312
rect 154132 17308 154138 17310
rect 423765 17307 423831 17310
rect 155718 17172 155724 17236
rect 155788 17234 155794 17236
rect 440325 17234 440391 17237
rect 155788 17232 440391 17234
rect 155788 17176 440330 17232
rect 440386 17176 440391 17232
rect 155788 17174 440391 17176
rect 155788 17172 155794 17174
rect 440325 17171 440391 17174
rect 144310 16220 144316 16284
rect 144380 16282 144386 16284
rect 295609 16282 295675 16285
rect 144380 16280 295675 16282
rect 144380 16224 295614 16280
rect 295670 16224 295675 16280
rect 144380 16222 295675 16224
rect 144380 16220 144386 16222
rect 295609 16219 295675 16222
rect 148542 16084 148548 16148
rect 148612 16146 148618 16148
rect 349153 16146 349219 16149
rect 148612 16144 349219 16146
rect 148612 16088 349158 16144
rect 349214 16088 349219 16144
rect 148612 16086 349219 16088
rect 148612 16084 148618 16086
rect 349153 16083 349219 16086
rect 152406 15948 152412 16012
rect 152476 16010 152482 16012
rect 406009 16010 406075 16013
rect 152476 16008 406075 16010
rect 152476 15952 406014 16008
rect 406070 15952 406075 16008
rect 152476 15950 406075 15952
rect 152476 15948 152482 15950
rect 406009 15947 406075 15950
rect 154246 15812 154252 15876
rect 154316 15874 154322 15876
rect 420177 15874 420243 15877
rect 154316 15872 420243 15874
rect 154316 15816 420182 15872
rect 420238 15816 420243 15872
rect 154316 15814 420243 15816
rect 154316 15812 154322 15814
rect 420177 15811 420243 15814
rect 140998 15132 141004 15196
rect 141068 15194 141074 15196
rect 264145 15194 264211 15197
rect 141068 15192 264211 15194
rect 141068 15136 264150 15192
rect 264206 15136 264211 15192
rect 141068 15134 264211 15136
rect 141068 15132 141074 15134
rect 264145 15131 264211 15134
rect 144494 14996 144500 15060
rect 144564 15058 144570 15060
rect 297265 15058 297331 15061
rect 144564 15056 297331 15058
rect 144564 15000 297270 15056
rect 297326 15000 297331 15056
rect 144564 14998 297331 15000
rect 144564 14996 144570 14998
rect 297265 14995 297331 14998
rect 145598 14860 145604 14924
rect 145668 14922 145674 14924
rect 316217 14922 316283 14925
rect 145668 14920 316283 14922
rect 145668 14864 316222 14920
rect 316278 14864 316283 14920
rect 145668 14862 316283 14864
rect 145668 14860 145674 14862
rect 316217 14859 316283 14862
rect 147070 14724 147076 14788
rect 147140 14786 147146 14788
rect 332685 14786 332751 14789
rect 147140 14784 332751 14786
rect 147140 14728 332690 14784
rect 332746 14728 332751 14784
rect 147140 14726 332751 14728
rect 147140 14724 147146 14726
rect 332685 14723 332751 14726
rect 151486 14588 151492 14652
rect 151556 14650 151562 14652
rect 387793 14650 387859 14653
rect 151556 14648 387859 14650
rect 151556 14592 387798 14648
rect 387854 14592 387859 14648
rect 151556 14590 387859 14592
rect 151556 14588 151562 14590
rect 387793 14587 387859 14590
rect 152590 14452 152596 14516
rect 152660 14514 152666 14516
rect 402513 14514 402579 14517
rect 152660 14512 402579 14514
rect 152660 14456 402518 14512
rect 402574 14456 402579 14512
rect 152660 14454 402579 14456
rect 152660 14452 152666 14454
rect 402513 14451 402579 14454
rect 140446 13636 140452 13700
rect 140516 13698 140522 13700
rect 242985 13698 243051 13701
rect 140516 13696 243051 13698
rect 140516 13640 242990 13696
rect 243046 13640 243051 13696
rect 140516 13638 243051 13640
rect 140516 13636 140522 13638
rect 242985 13635 243051 13638
rect 143022 13500 143028 13564
rect 143092 13562 143098 13564
rect 280705 13562 280771 13565
rect 143092 13560 280771 13562
rect 143092 13504 280710 13560
rect 280766 13504 280771 13560
rect 143092 13502 280771 13504
rect 143092 13500 143098 13502
rect 280705 13499 280771 13502
rect 149646 13364 149652 13428
rect 149716 13426 149722 13428
rect 365713 13426 365779 13429
rect 149716 13424 365779 13426
rect 149716 13368 365718 13424
rect 365774 13368 365779 13424
rect 149716 13366 365779 13368
rect 149716 13364 149722 13366
rect 365713 13363 365779 13366
rect 149830 13228 149836 13292
rect 149900 13290 149906 13292
rect 370129 13290 370195 13293
rect 149900 13288 370195 13290
rect 149900 13232 370134 13288
rect 370190 13232 370195 13288
rect 149900 13230 370195 13232
rect 149900 13228 149906 13230
rect 370129 13227 370195 13230
rect 154430 13092 154436 13156
rect 154500 13154 154506 13156
rect 418521 13154 418587 13157
rect 154500 13152 418587 13154
rect 154500 13096 418526 13152
rect 418582 13096 418587 13152
rect 154500 13094 418587 13096
rect 154500 13092 154506 13094
rect 418521 13091 418587 13094
rect 160870 12956 160876 13020
rect 160940 13018 160946 13020
rect 507209 13018 507275 13021
rect 160940 13016 507275 13018
rect 160940 12960 507214 13016
rect 507270 12960 507275 13016
rect 160940 12958 507275 12960
rect 160940 12956 160946 12958
rect 507209 12955 507275 12958
rect 138790 12820 138796 12884
rect 138860 12882 138866 12884
rect 225137 12882 225203 12885
rect 138860 12880 225203 12882
rect 138860 12824 225142 12880
rect 225198 12824 225203 12880
rect 138860 12822 225203 12824
rect 138860 12820 138866 12822
rect 225137 12819 225203 12822
rect 137870 12140 137876 12204
rect 137940 12202 137946 12204
rect 210969 12202 211035 12205
rect 137940 12200 211035 12202
rect 137940 12144 210974 12200
rect 211030 12144 211035 12200
rect 137940 12142 211035 12144
rect 137940 12140 137946 12142
rect 210969 12139 211035 12142
rect 148910 12004 148916 12068
rect 148980 12066 148986 12068
rect 349245 12066 349311 12069
rect 148980 12064 349311 12066
rect 148980 12008 349250 12064
rect 349306 12008 349311 12064
rect 148980 12006 349311 12008
rect 148980 12004 148986 12006
rect 349245 12003 349311 12006
rect 148726 11868 148732 11932
rect 148796 11930 148802 11932
rect 352833 11930 352899 11933
rect 148796 11928 352899 11930
rect 148796 11872 352838 11928
rect 352894 11872 352899 11928
rect 148796 11870 352899 11872
rect 148796 11868 148802 11870
rect 352833 11867 352899 11870
rect 150014 11732 150020 11796
rect 150084 11794 150090 11796
rect 365805 11794 365871 11797
rect 150084 11792 365871 11794
rect 150084 11736 365810 11792
rect 365866 11736 365871 11792
rect 150084 11734 365871 11736
rect 150084 11732 150090 11734
rect 365805 11731 365871 11734
rect 152774 11596 152780 11660
rect 152844 11658 152850 11660
rect 403617 11658 403683 11661
rect 152844 11656 403683 11658
rect 152844 11600 403622 11656
rect 403678 11600 403683 11656
rect 152844 11598 403683 11600
rect 152844 11596 152850 11598
rect 403617 11595 403683 11598
rect 89161 10434 89227 10437
rect 129038 10434 129044 10436
rect 89161 10432 129044 10434
rect 89161 10376 89166 10432
rect 89222 10376 129044 10432
rect 89161 10374 129044 10376
rect 89161 10371 89227 10374
rect 129038 10372 129044 10374
rect 129108 10372 129114 10436
rect 147254 10372 147260 10436
rect 147324 10434 147330 10436
rect 331213 10434 331279 10437
rect 147324 10432 331279 10434
rect 147324 10376 331218 10432
rect 331274 10376 331279 10432
rect 147324 10374 331279 10376
rect 147324 10372 147330 10374
rect 331213 10371 331279 10374
rect 71497 10298 71563 10301
rect 127198 10298 127204 10300
rect 71497 10296 127204 10298
rect 71497 10240 71502 10296
rect 71558 10240 127204 10296
rect 71497 10238 127204 10240
rect 71497 10235 71563 10238
rect 127198 10236 127204 10238
rect 127268 10236 127274 10300
rect 147438 10236 147444 10300
rect 147508 10298 147514 10300
rect 334617 10298 334683 10301
rect 147508 10296 334683 10298
rect 147508 10240 334622 10296
rect 334678 10240 334683 10296
rect 147508 10238 334683 10240
rect 147508 10236 147514 10238
rect 334617 10235 334683 10238
rect 109309 9482 109375 9485
rect 130142 9482 130148 9484
rect 109309 9480 130148 9482
rect 109309 9424 109314 9480
rect 109370 9424 130148 9480
rect 109309 9422 130148 9424
rect 109309 9419 109375 9422
rect 130142 9420 130148 9422
rect 130212 9420 130218 9484
rect 105721 9346 105787 9349
rect 129958 9346 129964 9348
rect 105721 9344 129964 9346
rect 105721 9288 105726 9344
rect 105782 9288 129964 9344
rect 105721 9286 129964 9288
rect 105721 9283 105787 9286
rect 129958 9284 129964 9286
rect 130028 9284 130034 9348
rect 53741 9210 53807 9213
rect 126094 9210 126100 9212
rect 53741 9208 126100 9210
rect 53741 9152 53746 9208
rect 53802 9152 126100 9208
rect 53741 9150 126100 9152
rect 53741 9147 53807 9150
rect 126094 9148 126100 9150
rect 126164 9148 126170 9212
rect 144678 9148 144684 9212
rect 144748 9210 144754 9212
rect 299657 9210 299723 9213
rect 144748 9208 299723 9210
rect 144748 9152 299662 9208
rect 299718 9152 299723 9208
rect 144748 9150 299723 9152
rect 144748 9148 144754 9150
rect 299657 9147 299723 9150
rect 38377 9074 38443 9077
rect 124438 9074 124444 9076
rect 38377 9072 124444 9074
rect 38377 9016 38382 9072
rect 38438 9016 124444 9072
rect 38377 9014 124444 9016
rect 38377 9011 38443 9014
rect 124438 9012 124444 9014
rect 124508 9012 124514 9076
rect 166574 9012 166580 9076
rect 166644 9074 166650 9076
rect 576301 9074 576367 9077
rect 166644 9072 576367 9074
rect 166644 9016 576306 9072
rect 576362 9016 576367 9072
rect 166644 9014 576367 9016
rect 166644 9012 166650 9014
rect 576301 9011 576367 9014
rect 34789 8938 34855 8941
rect 124622 8938 124628 8940
rect 34789 8936 124628 8938
rect 34789 8880 34794 8936
rect 34850 8880 124628 8936
rect 34789 8878 124628 8880
rect 34789 8875 34855 8878
rect 124622 8876 124628 8878
rect 124692 8876 124698 8940
rect 166390 8876 166396 8940
rect 166460 8938 166466 8940
rect 578601 8938 578667 8941
rect 166460 8936 578667 8938
rect 166460 8880 578606 8936
rect 578662 8880 578667 8936
rect 166460 8878 578667 8880
rect 166460 8876 166466 8878
rect 578601 8875 578667 8878
rect 135110 8060 135116 8124
rect 135180 8122 135186 8124
rect 169661 8122 169727 8125
rect 135180 8120 169727 8122
rect 135180 8064 169666 8120
rect 169722 8064 169727 8120
rect 135180 8062 169727 8064
rect 135180 8060 135186 8062
rect 169661 8059 169727 8062
rect 143390 7924 143396 7988
rect 143460 7986 143466 7988
rect 278313 7986 278379 7989
rect 143460 7984 278379 7986
rect 143460 7928 278318 7984
rect 278374 7928 278379 7984
rect 143460 7926 278379 7928
rect 143460 7924 143466 7926
rect 278313 7923 278379 7926
rect 91553 7850 91619 7853
rect 128670 7850 128676 7852
rect 91553 7848 128676 7850
rect 91553 7792 91558 7848
rect 91614 7792 128676 7848
rect 91553 7790 128676 7792
rect 91553 7787 91619 7790
rect 128670 7788 128676 7790
rect 128740 7788 128746 7852
rect 143206 7788 143212 7852
rect 143276 7850 143282 7852
rect 281901 7850 281967 7853
rect 143276 7848 281967 7850
rect 143276 7792 281906 7848
rect 281962 7792 281967 7848
rect 143276 7790 281967 7792
rect 143276 7788 143282 7790
rect 281901 7787 281967 7790
rect 87965 7714 88031 7717
rect 128854 7714 128860 7716
rect 87965 7712 128860 7714
rect 87965 7656 87970 7712
rect 88026 7656 128860 7712
rect 87965 7654 128860 7656
rect 87965 7651 88031 7654
rect 128854 7652 128860 7654
rect 128924 7652 128930 7716
rect 165102 7652 165108 7716
rect 165172 7714 165178 7716
rect 562041 7714 562107 7717
rect 165172 7712 562107 7714
rect 165172 7656 562046 7712
rect 562102 7656 562107 7712
rect 165172 7654 562107 7656
rect 165172 7652 165178 7654
rect 562041 7651 562107 7654
rect 70301 7578 70367 7581
rect 127014 7578 127020 7580
rect 70301 7576 127020 7578
rect 70301 7520 70306 7576
rect 70362 7520 127020 7576
rect 70301 7518 127020 7520
rect 70301 7515 70367 7518
rect 127014 7516 127020 7518
rect 127084 7516 127090 7580
rect 164918 7516 164924 7580
rect 164988 7578 164994 7580
rect 564433 7578 564499 7581
rect 164988 7576 564499 7578
rect 164988 7520 564438 7576
rect 564494 7520 564499 7576
rect 164988 7518 564499 7520
rect 164988 7516 164994 7518
rect 564433 7515 564499 7518
rect 139158 6836 139164 6900
rect 139228 6898 139234 6900
rect 226425 6898 226491 6901
rect 139228 6896 226491 6898
rect 139228 6840 226430 6896
rect 226486 6840 226491 6896
rect 139228 6838 226491 6840
rect 139228 6836 139234 6838
rect 226425 6835 226491 6838
rect 138974 6700 138980 6764
rect 139044 6762 139050 6764
rect 228725 6762 228791 6765
rect 139044 6760 228791 6762
rect 139044 6704 228730 6760
rect 228786 6704 228791 6760
rect 139044 6702 228791 6704
rect 139044 6700 139050 6702
rect 228725 6699 228791 6702
rect 108113 6626 108179 6629
rect 129774 6626 129780 6628
rect 108113 6624 129780 6626
rect -960 6490 480 6580
rect 108113 6568 108118 6624
rect 108174 6568 129780 6624
rect 108113 6566 129780 6568
rect 108113 6563 108179 6566
rect 129774 6564 129780 6566
rect 129844 6564 129850 6628
rect 140630 6564 140636 6628
rect 140700 6626 140706 6628
rect 246389 6626 246455 6629
rect 140700 6624 246455 6626
rect 140700 6568 246394 6624
rect 246450 6568 246455 6624
rect 140700 6566 246455 6568
rect 140700 6564 140706 6566
rect 246389 6563 246455 6566
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 3509 6490 3575 6493
rect -960 6488 3575 6490
rect -960 6432 3514 6488
rect 3570 6432 3575 6488
rect -960 6430 3575 6432
rect -960 6340 480 6430
rect 3509 6427 3575 6430
rect 56041 6490 56107 6493
rect 125910 6490 125916 6492
rect 56041 6488 125916 6490
rect 56041 6432 56046 6488
rect 56102 6432 125916 6488
rect 56041 6430 125916 6432
rect 56041 6427 56107 6430
rect 125910 6428 125916 6430
rect 125980 6428 125986 6492
rect 151670 6428 151676 6492
rect 151740 6490 151746 6492
rect 385953 6490 386019 6493
rect 151740 6488 386019 6490
rect 151740 6432 385958 6488
rect 386014 6432 386019 6488
rect 583520 6476 584960 6566
rect 151740 6430 386019 6432
rect 151740 6428 151746 6430
rect 385953 6427 386019 6430
rect 52545 6354 52611 6357
rect 125726 6354 125732 6356
rect 52545 6352 125732 6354
rect 52545 6296 52550 6352
rect 52606 6296 125732 6352
rect 52545 6294 125732 6296
rect 52545 6291 52611 6294
rect 125726 6292 125732 6294
rect 125796 6292 125802 6356
rect 162710 6292 162716 6356
rect 162780 6354 162786 6356
rect 526621 6354 526687 6357
rect 162780 6352 526687 6354
rect 162780 6296 526626 6352
rect 526682 6296 526687 6352
rect 162780 6294 526687 6296
rect 162780 6292 162786 6294
rect 526621 6291 526687 6294
rect 18229 6218 18295 6221
rect 122966 6218 122972 6220
rect 18229 6216 122972 6218
rect 18229 6160 18234 6216
rect 18290 6160 122972 6216
rect 18229 6158 122972 6160
rect 18229 6155 18295 6158
rect 122966 6156 122972 6158
rect 123036 6156 123042 6220
rect 162526 6156 162532 6220
rect 162596 6218 162602 6220
rect 530117 6218 530183 6221
rect 162596 6216 530183 6218
rect 162596 6160 530122 6216
rect 530178 6160 530183 6216
rect 162596 6158 530183 6160
rect 162596 6156 162602 6158
rect 530117 6155 530183 6158
rect 152958 5476 152964 5540
rect 153028 5538 153034 5540
rect 404813 5538 404879 5541
rect 153028 5536 404879 5538
rect 153028 5480 404818 5536
rect 404874 5480 404879 5536
rect 153028 5478 404879 5480
rect 153028 5476 153034 5478
rect 404813 5475 404879 5478
rect 161238 5340 161244 5404
rect 161308 5402 161314 5404
rect 508865 5402 508931 5405
rect 161308 5400 508931 5402
rect 161308 5344 508870 5400
rect 508926 5344 508931 5400
rect 161308 5342 508931 5344
rect 161308 5340 161314 5342
rect 508865 5339 508931 5342
rect 161054 5204 161060 5268
rect 161124 5266 161130 5268
rect 512453 5266 512519 5269
rect 161124 5264 512519 5266
rect 161124 5208 512458 5264
rect 512514 5208 512519 5264
rect 161124 5206 512519 5208
rect 161124 5204 161130 5206
rect 512453 5203 512519 5206
rect 163630 5068 163636 5132
rect 163700 5130 163706 5132
rect 547873 5130 547939 5133
rect 163700 5128 547939 5130
rect 163700 5072 547878 5128
rect 547934 5072 547939 5128
rect 163700 5070 547939 5072
rect 163700 5068 163706 5070
rect 547873 5067 547939 5070
rect 90357 4994 90423 4997
rect 128670 4994 128676 4996
rect 90357 4992 128676 4994
rect 90357 4936 90362 4992
rect 90418 4936 128676 4992
rect 90357 4934 128676 4936
rect 90357 4931 90423 4934
rect 128670 4932 128676 4934
rect 128740 4932 128746 4996
rect 133270 4932 133276 4996
rect 133340 4994 133346 4996
rect 155401 4994 155467 4997
rect 133340 4992 155467 4994
rect 133340 4936 155406 4992
rect 155462 4936 155467 4992
rect 133340 4934 155467 4936
rect 133340 4932 133346 4934
rect 155401 4931 155467 4934
rect 165470 4932 165476 4996
rect 165540 4994 165546 4996
rect 563237 4994 563303 4997
rect 165540 4992 563303 4994
rect 165540 4936 563242 4992
rect 563298 4936 563303 4992
rect 165540 4934 563303 4936
rect 165540 4932 165546 4934
rect 563237 4931 563303 4934
rect 37181 4858 37247 4861
rect 124254 4858 124260 4860
rect 37181 4856 124260 4858
rect 37181 4800 37186 4856
rect 37242 4800 124260 4856
rect 37181 4798 124260 4800
rect 37181 4795 37247 4798
rect 124254 4796 124260 4798
rect 124324 4796 124330 4860
rect 133454 4796 133460 4860
rect 133524 4858 133530 4860
rect 156597 4858 156663 4861
rect 133524 4856 156663 4858
rect 133524 4800 156602 4856
rect 156658 4800 156663 4856
rect 133524 4798 156663 4800
rect 133524 4796 133530 4798
rect 156597 4795 156663 4798
rect 165286 4796 165292 4860
rect 165356 4858 165362 4860
rect 565629 4858 565695 4861
rect 165356 4856 565695 4858
rect 165356 4800 565634 4856
rect 565690 4800 565695 4856
rect 165356 4798 565695 4800
rect 165356 4796 165362 4798
rect 565629 4795 565695 4798
rect 136398 4660 136404 4724
rect 136468 4722 136474 4724
rect 193305 4722 193371 4725
rect 136468 4720 193371 4722
rect 136468 4664 193310 4720
rect 193366 4664 193371 4720
rect 136468 4662 193371 4664
rect 136468 4660 136474 4662
rect 193305 4659 193371 4662
rect 159030 3980 159036 4044
rect 159100 4042 159106 4044
rect 494697 4042 494763 4045
rect 159100 4040 494763 4042
rect 159100 3984 494702 4040
rect 494758 3984 494763 4040
rect 159100 3982 494763 3984
rect 159100 3980 159106 3982
rect 494697 3979 494763 3982
rect 160829 3906 160895 3909
rect 505369 3906 505435 3909
rect 160829 3904 505435 3906
rect 160829 3848 160834 3904
rect 160890 3848 505374 3904
rect 505430 3848 505435 3904
rect 160829 3846 505435 3848
rect 160829 3843 160895 3846
rect 505369 3843 505435 3846
rect 54937 3770 55003 3773
rect 125542 3770 125548 3772
rect 54937 3768 125548 3770
rect 54937 3712 54942 3768
rect 54998 3712 125548 3768
rect 54937 3710 125548 3712
rect 54937 3707 55003 3710
rect 125542 3708 125548 3710
rect 125612 3708 125618 3772
rect 167494 3708 167500 3772
rect 167564 3770 167570 3772
rect 515949 3770 516015 3773
rect 167564 3768 516015 3770
rect 167564 3712 515954 3768
rect 516010 3712 516015 3768
rect 167564 3710 516015 3712
rect 167564 3708 167570 3710
rect 515949 3707 516015 3710
rect 17033 3634 17099 3637
rect 122598 3634 122604 3636
rect 17033 3632 122604 3634
rect 17033 3576 17038 3632
rect 17094 3576 122604 3632
rect 17033 3574 122604 3576
rect 17033 3571 17099 3574
rect 122598 3572 122604 3574
rect 122668 3572 122674 3636
rect 123477 3634 123543 3637
rect 131062 3634 131068 3636
rect 123477 3632 131068 3634
rect 123477 3576 123482 3632
rect 123538 3576 131068 3632
rect 123477 3574 131068 3576
rect 123477 3571 123543 3574
rect 131062 3572 131068 3574
rect 131132 3572 131138 3636
rect 131798 3572 131804 3636
rect 131868 3634 131874 3636
rect 137645 3634 137711 3637
rect 131868 3632 137711 3634
rect 131868 3576 137650 3632
rect 137706 3576 137711 3632
rect 131868 3574 137711 3576
rect 131868 3572 131874 3574
rect 137645 3571 137711 3574
rect 167678 3572 167684 3636
rect 167748 3634 167754 3636
rect 533705 3634 533771 3637
rect 167748 3632 533771 3634
rect 167748 3576 533710 3632
rect 533766 3576 533771 3632
rect 167748 3574 533771 3576
rect 167748 3572 167754 3574
rect 533705 3571 533771 3574
rect 1669 3498 1735 3501
rect 121678 3498 121684 3500
rect 1669 3496 121684 3498
rect 1669 3440 1674 3496
rect 1730 3440 121684 3496
rect 1669 3438 121684 3440
rect 1669 3435 1735 3438
rect 121678 3436 121684 3438
rect 121748 3436 121754 3500
rect 124673 3498 124739 3501
rect 131246 3498 131252 3500
rect 124673 3496 131252 3498
rect 124673 3440 124678 3496
rect 124734 3440 131252 3496
rect 124673 3438 131252 3440
rect 124673 3435 124739 3438
rect 131246 3436 131252 3438
rect 131316 3436 131322 3500
rect 131982 3436 131988 3500
rect 132052 3498 132058 3500
rect 140037 3498 140103 3501
rect 132052 3496 140103 3498
rect 132052 3440 140042 3496
rect 140098 3440 140103 3496
rect 132052 3438 140103 3440
rect 132052 3436 132058 3438
rect 140037 3435 140103 3438
rect 167862 3436 167868 3500
rect 167932 3498 167938 3500
rect 537201 3498 537267 3501
rect 167932 3496 537267 3498
rect 167932 3440 537206 3496
rect 537262 3440 537267 3496
rect 167932 3438 537267 3440
rect 167932 3436 167938 3438
rect 537201 3435 537267 3438
rect 565 3362 631 3365
rect 121494 3362 121500 3364
rect 565 3360 121500 3362
rect 565 3304 570 3360
rect 626 3304 121500 3360
rect 565 3302 121500 3304
rect 565 3299 631 3302
rect 121494 3300 121500 3302
rect 121564 3300 121570 3364
rect 133638 3300 133644 3364
rect 133708 3362 133714 3364
rect 157793 3362 157859 3365
rect 133708 3360 157859 3362
rect 133708 3304 157798 3360
rect 157854 3304 157859 3360
rect 133708 3302 157859 3304
rect 133708 3300 133714 3302
rect 157793 3299 157859 3302
rect 166758 3300 166764 3364
rect 166828 3362 166834 3364
rect 583385 3362 583451 3365
rect 166828 3360 583451 3362
rect 166828 3304 583390 3360
rect 583446 3304 583451 3360
rect 166828 3302 583451 3304
rect 166828 3300 166834 3302
rect 583385 3299 583451 3302
<< via3 >>
rect 580764 697172 580828 697236
rect 3372 658140 3436 658204
rect 396580 470596 396644 470660
rect 396764 240076 396828 240140
rect 396948 239940 397012 240004
rect 396764 232052 396828 232116
rect 396948 231100 397012 231164
rect 143396 193292 143460 193356
rect 155172 193292 155236 193356
rect 143580 191568 143644 191632
rect 144500 190980 144564 191044
rect 145788 189816 145852 189820
rect 145788 189760 145838 189816
rect 145838 189760 145852 189816
rect 145788 189756 145852 189760
rect 144500 189212 144564 189276
rect 155172 188940 155236 189004
rect 141188 184316 141252 184380
rect 140820 184240 140884 184244
rect 140820 184184 140834 184240
rect 140834 184184 140884 184240
rect 140820 184180 140884 184184
rect 142844 184044 142908 184108
rect 147260 182004 147324 182068
rect 143396 181188 143460 181252
rect 143396 180916 143460 180980
rect 142292 179012 142356 179076
rect 142844 178876 142908 178940
rect 141188 178740 141252 178804
rect 140820 178604 140884 178668
rect 147260 174524 147324 174588
rect 141924 137940 141988 138004
rect 143580 137668 143644 137732
rect 146156 137532 146220 137596
rect 143396 137396 143460 137460
rect 396580 137260 396644 137324
rect 168420 75380 168484 75444
rect 167684 75244 167748 75308
rect 168604 75244 168668 75308
rect 168604 75108 168668 75172
rect 168420 74972 168484 75036
rect 162900 74836 162964 74900
rect 580764 75244 580828 75308
rect 167500 74700 167564 74764
rect 169156 74836 169220 74900
rect 169340 74760 169404 74764
rect 169340 74704 169354 74760
rect 169354 74704 169404 74760
rect 169340 74700 169404 74704
rect 3372 74428 3436 74492
rect 128492 73128 128556 73132
rect 128492 73072 128542 73128
rect 128542 73072 128556 73128
rect 128492 73068 128556 73072
rect 149468 72932 149532 72996
rect 153884 72932 153948 72996
rect 162164 72932 162228 72996
rect 167500 73068 167564 73132
rect 148732 72796 148796 72860
rect 149836 72796 149900 72860
rect 151492 72796 151556 72860
rect 152780 72796 152844 72860
rect 154436 72796 154500 72860
rect 155540 72796 155604 72860
rect 157196 72796 157260 72860
rect 158300 72796 158364 72860
rect 158852 72796 158916 72860
rect 160692 72796 160756 72860
rect 162532 72796 162596 72860
rect 163268 72796 163332 72860
rect 165292 72796 165356 72860
rect 167684 72932 167748 72996
rect 167868 72796 167932 72860
rect 148916 72660 148980 72724
rect 150020 72720 150084 72724
rect 150020 72664 150034 72720
rect 150034 72664 150084 72720
rect 150020 72660 150084 72664
rect 151676 72660 151740 72724
rect 152964 72720 153028 72724
rect 152964 72664 153014 72720
rect 153014 72664 153028 72720
rect 152964 72660 153028 72664
rect 154252 72720 154316 72724
rect 154252 72664 154266 72720
rect 154266 72664 154316 72720
rect 154252 72660 154316 72664
rect 155724 72660 155788 72724
rect 156828 72720 156892 72724
rect 156828 72664 156878 72720
rect 156878 72664 156892 72720
rect 156828 72660 156892 72664
rect 157012 72660 157076 72724
rect 158484 72660 158548 72724
rect 159036 72660 159100 72724
rect 160876 72660 160940 72724
rect 162716 72660 162780 72724
rect 163452 72660 163516 72724
rect 165108 72660 165172 72724
rect 166212 72660 166276 72724
rect 166764 72720 166828 72724
rect 166764 72664 166814 72720
rect 166814 72664 166828 72720
rect 166764 72660 166828 72664
rect 166948 72660 167012 72724
rect 148364 72524 148428 72588
rect 149652 72524 149716 72588
rect 152412 72524 152476 72588
rect 154068 72524 154132 72588
rect 156644 72524 156708 72588
rect 158116 72524 158180 72588
rect 161060 72524 161124 72588
rect 162348 72524 162412 72588
rect 164924 72524 164988 72588
rect 166580 72524 166644 72588
rect 148548 72388 148612 72452
rect 151308 72388 151372 72452
rect 152596 72388 152660 72452
rect 158668 72388 158732 72452
rect 161244 72388 161308 72452
rect 162900 72388 162964 72452
rect 163636 72388 163700 72452
rect 165476 72388 165540 72452
rect 166396 72388 166460 72452
rect 126100 72252 126164 72316
rect 142844 72252 142908 72316
rect 124628 72116 124692 72180
rect 125548 72116 125612 72180
rect 129044 72116 129108 72180
rect 129964 72116 130028 72180
rect 133276 72116 133340 72180
rect 134748 72116 134812 72180
rect 136036 72116 136100 72180
rect 138980 72116 139044 72180
rect 140084 72116 140148 72180
rect 143028 72116 143092 72180
rect 144132 72116 144196 72180
rect 145236 72116 145300 72180
rect 146892 72116 146956 72180
rect 121684 72040 121748 72044
rect 121684 71984 121698 72040
rect 121698 71984 121748 72040
rect 121684 71980 121748 71984
rect 122788 72040 122852 72044
rect 122788 71984 122838 72040
rect 122838 71984 122852 72040
rect 122788 71980 122852 71984
rect 124260 71980 124324 72044
rect 125732 71980 125796 72044
rect 127204 71980 127268 72044
rect 128860 71980 128924 72044
rect 130148 71980 130212 72044
rect 131252 72040 131316 72044
rect 131252 71984 131266 72040
rect 131266 71984 131316 72040
rect 131252 71980 131316 71984
rect 131804 71980 131868 72044
rect 133460 71980 133524 72044
rect 134932 72040 134996 72044
rect 134932 71984 134982 72040
rect 134982 71984 134996 72040
rect 134932 71980 134996 71984
rect 136220 71980 136284 72044
rect 137692 71980 137756 72044
rect 138796 71980 138860 72044
rect 140268 71980 140332 72044
rect 140820 71980 140884 72044
rect 143212 71980 143276 72044
rect 144500 71980 144564 72044
rect 145420 71980 145484 72044
rect 147076 71980 147140 72044
rect 121500 71904 121564 71908
rect 121500 71848 121550 71904
rect 121550 71848 121564 71904
rect 121500 71844 121564 71848
rect 122972 71904 123036 71908
rect 122972 71848 122986 71904
rect 122986 71848 123036 71904
rect 122972 71844 123036 71848
rect 124444 71904 124508 71908
rect 124444 71848 124494 71904
rect 124494 71848 124508 71904
rect 124444 71844 124508 71848
rect 125916 71904 125980 71908
rect 125916 71848 125930 71904
rect 125930 71848 125980 71904
rect 125916 71844 125980 71848
rect 127020 71904 127084 71908
rect 127020 71848 127034 71904
rect 127034 71848 127084 71904
rect 127020 71844 127084 71848
rect 128676 71904 128740 71908
rect 128676 71848 128690 71904
rect 128690 71848 128740 71904
rect 128676 71844 128740 71848
rect 129780 71844 129844 71908
rect 131068 71904 131132 71908
rect 131068 71848 131118 71904
rect 131118 71848 131132 71904
rect 131068 71844 131132 71848
rect 131988 71844 132052 71908
rect 133644 71844 133708 71908
rect 135116 71904 135180 71908
rect 135116 71848 135166 71904
rect 135166 71848 135180 71904
rect 135116 71844 135180 71848
rect 135852 71844 135916 71908
rect 136404 71844 136468 71908
rect 137876 71904 137940 71908
rect 137876 71848 137926 71904
rect 137926 71848 137940 71904
rect 137876 71844 137940 71848
rect 138612 71844 138676 71908
rect 139164 71904 139228 71908
rect 139164 71848 139178 71904
rect 139178 71848 139228 71904
rect 139164 71844 139228 71848
rect 140452 71904 140516 71908
rect 140452 71848 140466 71904
rect 140466 71848 140516 71904
rect 140452 71844 140516 71848
rect 140636 71904 140700 71908
rect 140636 71848 140686 71904
rect 140686 71848 140700 71904
rect 140636 71844 140700 71848
rect 141004 71844 141068 71908
rect 143396 71844 143460 71908
rect 144316 71844 144380 71908
rect 144684 71844 144748 71908
rect 145604 71844 145668 71908
rect 147260 71904 147324 71908
rect 147260 71848 147310 71904
rect 147310 71848 147324 71904
rect 147260 71844 147324 71848
rect 147444 71844 147508 71908
rect 166948 71844 167012 71908
rect 158668 65452 158732 65516
rect 144132 35260 144196 35324
rect 146892 35124 146956 35188
rect 137692 34036 137756 34100
rect 140084 33900 140148 33964
rect 140820 33764 140884 33828
rect 134748 32676 134812 32740
rect 135852 32540 135916 32604
rect 136036 32404 136100 32468
rect 166212 31724 166276 31788
rect 163268 31180 163332 31244
rect 158116 31044 158180 31108
rect 158852 30908 158916 30972
rect 145236 29548 145300 29612
rect 136220 27100 136284 27164
rect 142844 26964 142908 27028
rect 149468 26828 149532 26892
rect 134932 25604 134996 25668
rect 156644 25468 156708 25532
rect 151308 24380 151372 24444
rect 162164 24244 162228 24308
rect 163452 24108 163516 24172
rect 156828 22748 156892 22812
rect 160692 22612 160756 22676
rect 148364 21524 148428 21588
rect 155540 21388 155604 21452
rect 158300 21252 158364 21316
rect 138612 20164 138676 20228
rect 140268 20028 140332 20092
rect 158484 19892 158548 19956
rect 157196 18804 157260 18868
rect 157012 18668 157076 18732
rect 162348 18532 162412 18596
rect 145420 17580 145484 17644
rect 153884 17444 153948 17508
rect 154068 17308 154132 17372
rect 155724 17172 155788 17236
rect 144316 16220 144380 16284
rect 148548 16084 148612 16148
rect 152412 15948 152476 16012
rect 154252 15812 154316 15876
rect 141004 15132 141068 15196
rect 144500 14996 144564 15060
rect 145604 14860 145668 14924
rect 147076 14724 147140 14788
rect 151492 14588 151556 14652
rect 152596 14452 152660 14516
rect 140452 13636 140516 13700
rect 143028 13500 143092 13564
rect 149652 13364 149716 13428
rect 149836 13228 149900 13292
rect 154436 13092 154500 13156
rect 160876 12956 160940 13020
rect 138796 12820 138860 12884
rect 137876 12140 137940 12204
rect 148916 12004 148980 12068
rect 148732 11868 148796 11932
rect 150020 11732 150084 11796
rect 152780 11596 152844 11660
rect 129044 10372 129108 10436
rect 147260 10372 147324 10436
rect 127204 10236 127268 10300
rect 147444 10236 147508 10300
rect 130148 9420 130212 9484
rect 129964 9284 130028 9348
rect 126100 9148 126164 9212
rect 144684 9148 144748 9212
rect 124444 9012 124508 9076
rect 166580 9012 166644 9076
rect 124628 8876 124692 8940
rect 166396 8876 166460 8940
rect 135116 8060 135180 8124
rect 143396 7924 143460 7988
rect 128676 7788 128740 7852
rect 143212 7788 143276 7852
rect 128860 7652 128924 7716
rect 165108 7652 165172 7716
rect 127020 7516 127084 7580
rect 164924 7516 164988 7580
rect 139164 6836 139228 6900
rect 138980 6700 139044 6764
rect 129780 6564 129844 6628
rect 140636 6564 140700 6628
rect 125916 6428 125980 6492
rect 151676 6428 151740 6492
rect 125732 6292 125796 6356
rect 162716 6292 162780 6356
rect 122972 6156 123036 6220
rect 162532 6156 162596 6220
rect 152964 5476 153028 5540
rect 161244 5340 161308 5404
rect 161060 5204 161124 5268
rect 163636 5068 163700 5132
rect 128676 4932 128740 4996
rect 133276 4932 133340 4996
rect 165476 4932 165540 4996
rect 124260 4796 124324 4860
rect 133460 4796 133524 4860
rect 165292 4796 165356 4860
rect 136404 4660 136468 4724
rect 159036 3980 159100 4044
rect 125548 3708 125612 3772
rect 167500 3708 167564 3772
rect 122604 3572 122668 3636
rect 131068 3572 131132 3636
rect 131804 3572 131868 3636
rect 167684 3572 167748 3636
rect 121684 3436 121748 3500
rect 131252 3436 131316 3500
rect 131988 3436 132052 3500
rect 167868 3436 167932 3500
rect 121500 3300 121564 3364
rect 133644 3300 133708 3364
rect 166764 3300 166828 3364
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 682954 -8106 711002
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 -8106 682954
rect -8726 682634 -8106 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 -8106 682634
rect -8726 646954 -8106 682398
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 -8106 646954
rect -8726 646634 -8106 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 -8106 646634
rect -8726 610954 -8106 646398
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 -8106 610954
rect -8726 610634 -8106 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 -8106 610634
rect -8726 574954 -8106 610398
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 -8106 574954
rect -8726 574634 -8106 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 -8106 574634
rect -8726 538954 -8106 574398
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 -8106 538954
rect -8726 538634 -8106 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 -8106 538634
rect -8726 502954 -8106 538398
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 -8106 502954
rect -8726 502634 -8106 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 -8106 502634
rect -8726 466954 -8106 502398
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 -8106 466954
rect -8726 466634 -8106 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 -8106 466634
rect -8726 430954 -8106 466398
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 -8106 430954
rect -8726 430634 -8106 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 -8106 430634
rect -8726 394954 -8106 430398
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 -8106 394954
rect -8726 394634 -8106 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 -8106 394634
rect -8726 358954 -8106 394398
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 -8106 358954
rect -8726 358634 -8106 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 -8106 358634
rect -8726 322954 -8106 358398
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 -8106 322954
rect -8726 322634 -8106 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 -8106 322634
rect -8726 286954 -8106 322398
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 -8106 286954
rect -8726 286634 -8106 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 -8106 286634
rect -8726 250954 -8106 286398
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 -8106 250954
rect -8726 250634 -8106 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 -8106 250634
rect -8726 214954 -8106 250398
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 -8106 214954
rect -8726 214634 -8106 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 -8106 214634
rect -8726 178954 -8106 214398
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 -8106 178954
rect -8726 178634 -8106 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 -8106 178634
rect -8726 142954 -8106 178398
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 -8106 142954
rect -8726 142634 -8106 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 -8106 142634
rect -8726 106954 -8106 142398
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 -8106 106954
rect -8726 106634 -8106 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 -8106 106634
rect -8726 70954 -8106 106398
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 -8106 70954
rect -8726 70634 -8106 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 -8106 70634
rect -8726 34954 -8106 70398
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 -8106 34954
rect -8726 34634 -8106 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 -8106 34634
rect -8726 -7066 -8106 34398
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 678454 -7146 710042
rect -7766 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 -7146 678454
rect -7766 678134 -7146 678218
rect -7766 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 -7146 678134
rect -7766 642454 -7146 677898
rect -7766 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 -7146 642454
rect -7766 642134 -7146 642218
rect -7766 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 -7146 642134
rect -7766 606454 -7146 641898
rect -7766 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 -7146 606454
rect -7766 606134 -7146 606218
rect -7766 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 -7146 606134
rect -7766 570454 -7146 605898
rect -7766 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 -7146 570454
rect -7766 570134 -7146 570218
rect -7766 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 -7146 570134
rect -7766 534454 -7146 569898
rect -7766 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 -7146 534454
rect -7766 534134 -7146 534218
rect -7766 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 -7146 534134
rect -7766 498454 -7146 533898
rect -7766 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 -7146 498454
rect -7766 498134 -7146 498218
rect -7766 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 -7146 498134
rect -7766 462454 -7146 497898
rect -7766 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 -7146 462454
rect -7766 462134 -7146 462218
rect -7766 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 -7146 462134
rect -7766 426454 -7146 461898
rect -7766 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 -7146 426454
rect -7766 426134 -7146 426218
rect -7766 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 -7146 426134
rect -7766 390454 -7146 425898
rect -7766 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 -7146 390454
rect -7766 390134 -7146 390218
rect -7766 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 -7146 390134
rect -7766 354454 -7146 389898
rect -7766 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 -7146 354454
rect -7766 354134 -7146 354218
rect -7766 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 -7146 354134
rect -7766 318454 -7146 353898
rect -7766 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 -7146 318454
rect -7766 318134 -7146 318218
rect -7766 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 -7146 318134
rect -7766 282454 -7146 317898
rect -7766 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 -7146 282454
rect -7766 282134 -7146 282218
rect -7766 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 -7146 282134
rect -7766 246454 -7146 281898
rect -7766 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 -7146 246454
rect -7766 246134 -7146 246218
rect -7766 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 -7146 246134
rect -7766 210454 -7146 245898
rect -7766 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 -7146 210454
rect -7766 210134 -7146 210218
rect -7766 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 -7146 210134
rect -7766 174454 -7146 209898
rect -7766 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 -7146 174454
rect -7766 174134 -7146 174218
rect -7766 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 -7146 174134
rect -7766 138454 -7146 173898
rect -7766 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 -7146 138454
rect -7766 138134 -7146 138218
rect -7766 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 -7146 138134
rect -7766 102454 -7146 137898
rect -7766 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 -7146 102454
rect -7766 102134 -7146 102218
rect -7766 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 -7146 102134
rect -7766 66454 -7146 101898
rect -7766 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 -7146 66454
rect -7766 66134 -7146 66218
rect -7766 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 -7146 66134
rect -7766 30454 -7146 65898
rect -7766 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 -7146 30454
rect -7766 30134 -7146 30218
rect -7766 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 -7146 30134
rect -7766 -6106 -7146 29898
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 673954 -6186 709082
rect -6806 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 -6186 673954
rect -6806 673634 -6186 673718
rect -6806 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 -6186 673634
rect -6806 637954 -6186 673398
rect -6806 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 -6186 637954
rect -6806 637634 -6186 637718
rect -6806 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 -6186 637634
rect -6806 601954 -6186 637398
rect -6806 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 -6186 601954
rect -6806 601634 -6186 601718
rect -6806 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 -6186 601634
rect -6806 565954 -6186 601398
rect -6806 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 -6186 565954
rect -6806 565634 -6186 565718
rect -6806 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 -6186 565634
rect -6806 529954 -6186 565398
rect -6806 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 -6186 529954
rect -6806 529634 -6186 529718
rect -6806 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 -6186 529634
rect -6806 493954 -6186 529398
rect -6806 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 -6186 493954
rect -6806 493634 -6186 493718
rect -6806 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 -6186 493634
rect -6806 457954 -6186 493398
rect -6806 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 -6186 457954
rect -6806 457634 -6186 457718
rect -6806 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 -6186 457634
rect -6806 421954 -6186 457398
rect -6806 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 -6186 421954
rect -6806 421634 -6186 421718
rect -6806 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 -6186 421634
rect -6806 385954 -6186 421398
rect -6806 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 -6186 385954
rect -6806 385634 -6186 385718
rect -6806 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 -6186 385634
rect -6806 349954 -6186 385398
rect -6806 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 -6186 349954
rect -6806 349634 -6186 349718
rect -6806 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 -6186 349634
rect -6806 313954 -6186 349398
rect -6806 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 -6186 313954
rect -6806 313634 -6186 313718
rect -6806 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 -6186 313634
rect -6806 277954 -6186 313398
rect -6806 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 -6186 277954
rect -6806 277634 -6186 277718
rect -6806 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 -6186 277634
rect -6806 241954 -6186 277398
rect -6806 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 -6186 241954
rect -6806 241634 -6186 241718
rect -6806 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 -6186 241634
rect -6806 205954 -6186 241398
rect -6806 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 -6186 205954
rect -6806 205634 -6186 205718
rect -6806 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 -6186 205634
rect -6806 169954 -6186 205398
rect -6806 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 -6186 169954
rect -6806 169634 -6186 169718
rect -6806 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 -6186 169634
rect -6806 133954 -6186 169398
rect -6806 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 -6186 133954
rect -6806 133634 -6186 133718
rect -6806 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 -6186 133634
rect -6806 97954 -6186 133398
rect -6806 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 -6186 97954
rect -6806 97634 -6186 97718
rect -6806 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 -6186 97634
rect -6806 61954 -6186 97398
rect -6806 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 -6186 61954
rect -6806 61634 -6186 61718
rect -6806 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 -6186 61634
rect -6806 25954 -6186 61398
rect -6806 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 -6186 25954
rect -6806 25634 -6186 25718
rect -6806 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 -6186 25634
rect -6806 -5146 -6186 25398
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 669454 -5226 708122
rect -5846 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 -5226 669454
rect -5846 669134 -5226 669218
rect -5846 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 -5226 669134
rect -5846 633454 -5226 668898
rect -5846 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 -5226 633454
rect -5846 633134 -5226 633218
rect -5846 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 -5226 633134
rect -5846 597454 -5226 632898
rect -5846 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 -5226 597454
rect -5846 597134 -5226 597218
rect -5846 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 -5226 597134
rect -5846 561454 -5226 596898
rect -5846 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 -5226 561454
rect -5846 561134 -5226 561218
rect -5846 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 -5226 561134
rect -5846 525454 -5226 560898
rect -5846 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 -5226 525454
rect -5846 525134 -5226 525218
rect -5846 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 -5226 525134
rect -5846 489454 -5226 524898
rect -5846 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 -5226 489454
rect -5846 489134 -5226 489218
rect -5846 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 -5226 489134
rect -5846 453454 -5226 488898
rect -5846 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 -5226 453454
rect -5846 453134 -5226 453218
rect -5846 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 -5226 453134
rect -5846 417454 -5226 452898
rect -5846 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 -5226 417454
rect -5846 417134 -5226 417218
rect -5846 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 -5226 417134
rect -5846 381454 -5226 416898
rect -5846 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 -5226 381454
rect -5846 381134 -5226 381218
rect -5846 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 -5226 381134
rect -5846 345454 -5226 380898
rect -5846 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 -5226 345454
rect -5846 345134 -5226 345218
rect -5846 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 -5226 345134
rect -5846 309454 -5226 344898
rect -5846 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 -5226 309454
rect -5846 309134 -5226 309218
rect -5846 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 -5226 309134
rect -5846 273454 -5226 308898
rect -5846 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 -5226 273454
rect -5846 273134 -5226 273218
rect -5846 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 -5226 273134
rect -5846 237454 -5226 272898
rect -5846 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 -5226 237454
rect -5846 237134 -5226 237218
rect -5846 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 -5226 237134
rect -5846 201454 -5226 236898
rect -5846 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 -5226 201454
rect -5846 201134 -5226 201218
rect -5846 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 -5226 201134
rect -5846 165454 -5226 200898
rect -5846 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 -5226 165454
rect -5846 165134 -5226 165218
rect -5846 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 -5226 165134
rect -5846 129454 -5226 164898
rect -5846 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 -5226 129454
rect -5846 129134 -5226 129218
rect -5846 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 -5226 129134
rect -5846 93454 -5226 128898
rect -5846 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 -5226 93454
rect -5846 93134 -5226 93218
rect -5846 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 -5226 93134
rect -5846 57454 -5226 92898
rect -5846 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 -5226 57454
rect -5846 57134 -5226 57218
rect -5846 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 -5226 57134
rect -5846 21454 -5226 56898
rect -5846 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 -5226 21454
rect -5846 21134 -5226 21218
rect -5846 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 -5226 21134
rect -5846 -4186 -5226 20898
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 700954 -4266 707162
rect -4886 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 -4266 700954
rect -4886 700634 -4266 700718
rect -4886 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 -4266 700634
rect -4886 664954 -4266 700398
rect -4886 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 -4266 664954
rect -4886 664634 -4266 664718
rect -4886 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 -4266 664634
rect -4886 628954 -4266 664398
rect -4886 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 -4266 628954
rect -4886 628634 -4266 628718
rect -4886 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 -4266 628634
rect -4886 592954 -4266 628398
rect -4886 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 -4266 592954
rect -4886 592634 -4266 592718
rect -4886 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 -4266 592634
rect -4886 556954 -4266 592398
rect -4886 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 -4266 556954
rect -4886 556634 -4266 556718
rect -4886 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 -4266 556634
rect -4886 520954 -4266 556398
rect -4886 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 -4266 520954
rect -4886 520634 -4266 520718
rect -4886 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 -4266 520634
rect -4886 484954 -4266 520398
rect -4886 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 -4266 484954
rect -4886 484634 -4266 484718
rect -4886 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 -4266 484634
rect -4886 448954 -4266 484398
rect -4886 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 -4266 448954
rect -4886 448634 -4266 448718
rect -4886 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 -4266 448634
rect -4886 412954 -4266 448398
rect -4886 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 -4266 412954
rect -4886 412634 -4266 412718
rect -4886 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 -4266 412634
rect -4886 376954 -4266 412398
rect -4886 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 -4266 376954
rect -4886 376634 -4266 376718
rect -4886 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 -4266 376634
rect -4886 340954 -4266 376398
rect -4886 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 -4266 340954
rect -4886 340634 -4266 340718
rect -4886 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 -4266 340634
rect -4886 304954 -4266 340398
rect -4886 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 -4266 304954
rect -4886 304634 -4266 304718
rect -4886 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 -4266 304634
rect -4886 268954 -4266 304398
rect -4886 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 -4266 268954
rect -4886 268634 -4266 268718
rect -4886 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 -4266 268634
rect -4886 232954 -4266 268398
rect -4886 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 -4266 232954
rect -4886 232634 -4266 232718
rect -4886 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 -4266 232634
rect -4886 196954 -4266 232398
rect -4886 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 -4266 196954
rect -4886 196634 -4266 196718
rect -4886 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 -4266 196634
rect -4886 160954 -4266 196398
rect -4886 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 -4266 160954
rect -4886 160634 -4266 160718
rect -4886 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 -4266 160634
rect -4886 124954 -4266 160398
rect -4886 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 -4266 124954
rect -4886 124634 -4266 124718
rect -4886 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 -4266 124634
rect -4886 88954 -4266 124398
rect -4886 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 -4266 88954
rect -4886 88634 -4266 88718
rect -4886 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 -4266 88634
rect -4886 52954 -4266 88398
rect -4886 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 -4266 52954
rect -4886 52634 -4266 52718
rect -4886 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 -4266 52634
rect -4886 16954 -4266 52398
rect -4886 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 -4266 16954
rect -4886 16634 -4266 16718
rect -4886 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 -4266 16634
rect -4886 -3226 -4266 16398
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 696454 -3306 706202
rect -3926 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 -3306 696454
rect -3926 696134 -3306 696218
rect -3926 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 -3306 696134
rect -3926 660454 -3306 695898
rect -3926 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 -3306 660454
rect -3926 660134 -3306 660218
rect -3926 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 -3306 660134
rect -3926 624454 -3306 659898
rect -3926 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 -3306 624454
rect -3926 624134 -3306 624218
rect -3926 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 -3306 624134
rect -3926 588454 -3306 623898
rect -3926 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 -3306 588454
rect -3926 588134 -3306 588218
rect -3926 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 -3306 588134
rect -3926 552454 -3306 587898
rect -3926 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 -3306 552454
rect -3926 552134 -3306 552218
rect -3926 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 -3306 552134
rect -3926 516454 -3306 551898
rect -3926 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 -3306 516454
rect -3926 516134 -3306 516218
rect -3926 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 -3306 516134
rect -3926 480454 -3306 515898
rect -3926 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 -3306 480454
rect -3926 480134 -3306 480218
rect -3926 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 -3306 480134
rect -3926 444454 -3306 479898
rect -3926 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 -3306 444454
rect -3926 444134 -3306 444218
rect -3926 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 -3306 444134
rect -3926 408454 -3306 443898
rect -3926 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 -3306 408454
rect -3926 408134 -3306 408218
rect -3926 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 -3306 408134
rect -3926 372454 -3306 407898
rect -3926 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 -3306 372454
rect -3926 372134 -3306 372218
rect -3926 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 -3306 372134
rect -3926 336454 -3306 371898
rect -3926 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 -3306 336454
rect -3926 336134 -3306 336218
rect -3926 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 -3306 336134
rect -3926 300454 -3306 335898
rect -3926 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 -3306 300454
rect -3926 300134 -3306 300218
rect -3926 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 -3306 300134
rect -3926 264454 -3306 299898
rect -3926 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 -3306 264454
rect -3926 264134 -3306 264218
rect -3926 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 -3306 264134
rect -3926 228454 -3306 263898
rect -3926 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 -3306 228454
rect -3926 228134 -3306 228218
rect -3926 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 -3306 228134
rect -3926 192454 -3306 227898
rect -3926 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 -3306 192454
rect -3926 192134 -3306 192218
rect -3926 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 -3306 192134
rect -3926 156454 -3306 191898
rect -3926 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 -3306 156454
rect -3926 156134 -3306 156218
rect -3926 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 -3306 156134
rect -3926 120454 -3306 155898
rect -3926 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 -3306 120454
rect -3926 120134 -3306 120218
rect -3926 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 -3306 120134
rect -3926 84454 -3306 119898
rect -3926 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 -3306 84454
rect -3926 84134 -3306 84218
rect -3926 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 -3306 84134
rect -3926 48454 -3306 83898
rect -3926 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 -3306 48454
rect -3926 48134 -3306 48218
rect -3926 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 -3306 48134
rect -3926 12454 -3306 47898
rect -3926 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 -3306 12454
rect -3926 12134 -3306 12218
rect -3926 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 -3306 12134
rect -3926 -2266 -3306 11898
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691954 -2346 705242
rect -2966 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 -2346 691954
rect -2966 691634 -2346 691718
rect -2966 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 -2346 691634
rect -2966 655954 -2346 691398
rect -2966 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 -2346 655954
rect -2966 655634 -2346 655718
rect -2966 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 -2346 655634
rect -2966 619954 -2346 655398
rect -2966 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 -2346 619954
rect -2966 619634 -2346 619718
rect -2966 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 -2346 619634
rect -2966 583954 -2346 619398
rect -2966 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 -2346 583954
rect -2966 583634 -2346 583718
rect -2966 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 -2346 583634
rect -2966 547954 -2346 583398
rect -2966 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 -2346 547954
rect -2966 547634 -2346 547718
rect -2966 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 -2346 547634
rect -2966 511954 -2346 547398
rect -2966 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 -2346 511954
rect -2966 511634 -2346 511718
rect -2966 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 -2346 511634
rect -2966 475954 -2346 511398
rect -2966 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 -2346 475954
rect -2966 475634 -2346 475718
rect -2966 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 -2346 475634
rect -2966 439954 -2346 475398
rect -2966 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 -2346 439954
rect -2966 439634 -2346 439718
rect -2966 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 -2346 439634
rect -2966 403954 -2346 439398
rect -2966 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 -2346 403954
rect -2966 403634 -2346 403718
rect -2966 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 -2346 403634
rect -2966 367954 -2346 403398
rect -2966 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 -2346 367954
rect -2966 367634 -2346 367718
rect -2966 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 -2346 367634
rect -2966 331954 -2346 367398
rect -2966 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 -2346 331954
rect -2966 331634 -2346 331718
rect -2966 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 -2346 331634
rect -2966 295954 -2346 331398
rect -2966 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 -2346 295954
rect -2966 295634 -2346 295718
rect -2966 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 -2346 295634
rect -2966 259954 -2346 295398
rect -2966 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 -2346 259954
rect -2966 259634 -2346 259718
rect -2966 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 -2346 259634
rect -2966 223954 -2346 259398
rect -2966 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 -2346 223954
rect -2966 223634 -2346 223718
rect -2966 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 -2346 223634
rect -2966 187954 -2346 223398
rect -2966 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 -2346 187954
rect -2966 187634 -2346 187718
rect -2966 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 -2346 187634
rect -2966 151954 -2346 187398
rect -2966 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 -2346 151954
rect -2966 151634 -2346 151718
rect -2966 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 -2346 151634
rect -2966 115954 -2346 151398
rect -2966 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 -2346 115954
rect -2966 115634 -2346 115718
rect -2966 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 -2346 115634
rect -2966 79954 -2346 115398
rect -2966 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 -2346 79954
rect -2966 79634 -2346 79718
rect -2966 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 -2346 79634
rect -2966 43954 -2346 79398
rect -2966 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 -2346 43954
rect -2966 43634 -2346 43718
rect -2966 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 -2346 43634
rect -2966 7954 -2346 43398
rect -2966 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 -2346 7954
rect -2966 7634 -2346 7718
rect -2966 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 -2346 7634
rect -2966 -1306 -2346 7398
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 6294 705798 6914 711590
rect 6294 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 6914 705798
rect 6294 705478 6914 705562
rect 6294 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 6914 705478
rect 6294 691954 6914 705242
rect 6294 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 6914 691954
rect 6294 691634 6914 691718
rect 6294 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 6914 691634
rect 3371 658204 3437 658205
rect 3371 658140 3372 658204
rect 3436 658140 3437 658204
rect 3371 658139 3437 658140
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 3374 74493 3434 658139
rect 6294 655954 6914 691398
rect 6294 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 6914 655954
rect 6294 655634 6914 655718
rect 6294 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 6914 655634
rect 6294 619954 6914 655398
rect 6294 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 6914 619954
rect 6294 619634 6914 619718
rect 6294 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 6914 619634
rect 6294 583954 6914 619398
rect 6294 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 6914 583954
rect 6294 583634 6914 583718
rect 6294 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 6914 583634
rect 6294 547954 6914 583398
rect 6294 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 6914 547954
rect 6294 547634 6914 547718
rect 6294 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 6914 547634
rect 6294 511954 6914 547398
rect 6294 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 6914 511954
rect 6294 511634 6914 511718
rect 6294 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 6914 511634
rect 6294 475954 6914 511398
rect 6294 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 6914 475954
rect 6294 475634 6914 475718
rect 6294 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 6914 475634
rect 6294 439954 6914 475398
rect 6294 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 6914 439954
rect 6294 439634 6914 439718
rect 6294 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 6914 439634
rect 6294 403954 6914 439398
rect 6294 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 6914 403954
rect 6294 403634 6914 403718
rect 6294 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 6914 403634
rect 6294 367954 6914 403398
rect 6294 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 6914 367954
rect 6294 367634 6914 367718
rect 6294 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 6914 367634
rect 6294 331954 6914 367398
rect 6294 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 6914 331954
rect 6294 331634 6914 331718
rect 6294 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 6914 331634
rect 6294 295954 6914 331398
rect 6294 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 6914 295954
rect 6294 295634 6914 295718
rect 6294 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 6914 295634
rect 6294 259954 6914 295398
rect 6294 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 6914 259954
rect 6294 259634 6914 259718
rect 6294 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 6914 259634
rect 6294 223954 6914 259398
rect 6294 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 6914 223954
rect 6294 223634 6914 223718
rect 6294 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 6914 223634
rect 6294 187954 6914 223398
rect 6294 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 6914 187954
rect 6294 187634 6914 187718
rect 6294 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 6914 187634
rect 6294 151954 6914 187398
rect 6294 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 6914 151954
rect 6294 151634 6914 151718
rect 6294 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 6914 151634
rect 6294 115954 6914 151398
rect 6294 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 6914 115954
rect 6294 115634 6914 115718
rect 6294 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 6914 115634
rect 6294 79954 6914 115398
rect 6294 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 6914 79954
rect 6294 79634 6914 79718
rect 6294 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 6914 79634
rect 3371 74492 3437 74493
rect 3371 74428 3372 74492
rect 3436 74428 3437 74492
rect 3371 74427 3437 74428
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 6294 43954 6914 79398
rect 6294 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 6914 43954
rect 6294 43634 6914 43718
rect 6294 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 6914 43634
rect 6294 7954 6914 43398
rect 6294 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 6914 7954
rect 6294 7634 6914 7718
rect 6294 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 6914 7634
rect 6294 -1306 6914 7398
rect 6294 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 6914 -1306
rect 6294 -1626 6914 -1542
rect 6294 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 6914 -1626
rect 6294 -7654 6914 -1862
rect 10794 706758 11414 711590
rect 10794 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 11414 706758
rect 10794 706438 11414 706522
rect 10794 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 11414 706438
rect 10794 696454 11414 706202
rect 10794 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 11414 696454
rect 10794 696134 11414 696218
rect 10794 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 11414 696134
rect 10794 660454 11414 695898
rect 10794 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 11414 660454
rect 10794 660134 11414 660218
rect 10794 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 11414 660134
rect 10794 624454 11414 659898
rect 10794 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 11414 624454
rect 10794 624134 11414 624218
rect 10794 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 11414 624134
rect 10794 588454 11414 623898
rect 10794 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 11414 588454
rect 10794 588134 11414 588218
rect 10794 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 11414 588134
rect 10794 552454 11414 587898
rect 10794 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 11414 552454
rect 10794 552134 11414 552218
rect 10794 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 11414 552134
rect 10794 516454 11414 551898
rect 10794 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 11414 516454
rect 10794 516134 11414 516218
rect 10794 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 11414 516134
rect 10794 480454 11414 515898
rect 10794 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 11414 480454
rect 10794 480134 11414 480218
rect 10794 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 11414 480134
rect 10794 444454 11414 479898
rect 10794 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 11414 444454
rect 10794 444134 11414 444218
rect 10794 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 11414 444134
rect 10794 408454 11414 443898
rect 10794 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 11414 408454
rect 10794 408134 11414 408218
rect 10794 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 11414 408134
rect 10794 372454 11414 407898
rect 10794 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 11414 372454
rect 10794 372134 11414 372218
rect 10794 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 11414 372134
rect 10794 336454 11414 371898
rect 10794 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 11414 336454
rect 10794 336134 11414 336218
rect 10794 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 11414 336134
rect 10794 300454 11414 335898
rect 10794 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 11414 300454
rect 10794 300134 11414 300218
rect 10794 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 11414 300134
rect 10794 264454 11414 299898
rect 10794 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 11414 264454
rect 10794 264134 11414 264218
rect 10794 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 11414 264134
rect 10794 228454 11414 263898
rect 10794 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 11414 228454
rect 10794 228134 11414 228218
rect 10794 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 11414 228134
rect 10794 192454 11414 227898
rect 10794 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 11414 192454
rect 10794 192134 11414 192218
rect 10794 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 11414 192134
rect 10794 156454 11414 191898
rect 10794 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 11414 156454
rect 10794 156134 11414 156218
rect 10794 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 11414 156134
rect 10794 120454 11414 155898
rect 10794 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 11414 120454
rect 10794 120134 11414 120218
rect 10794 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 11414 120134
rect 10794 84454 11414 119898
rect 10794 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 11414 84454
rect 10794 84134 11414 84218
rect 10794 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 11414 84134
rect 10794 48454 11414 83898
rect 10794 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 11414 48454
rect 10794 48134 11414 48218
rect 10794 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 11414 48134
rect 10794 12454 11414 47898
rect 10794 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 11414 12454
rect 10794 12134 11414 12218
rect 10794 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 11414 12134
rect 10794 -2266 11414 11898
rect 10794 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 11414 -2266
rect 10794 -2586 11414 -2502
rect 10794 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 11414 -2586
rect 10794 -7654 11414 -2822
rect 15294 707718 15914 711590
rect 15294 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 15914 707718
rect 15294 707398 15914 707482
rect 15294 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 15914 707398
rect 15294 700954 15914 707162
rect 15294 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 15914 700954
rect 15294 700634 15914 700718
rect 15294 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 15914 700634
rect 15294 664954 15914 700398
rect 15294 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 15914 664954
rect 15294 664634 15914 664718
rect 15294 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 15914 664634
rect 15294 628954 15914 664398
rect 15294 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 15914 628954
rect 15294 628634 15914 628718
rect 15294 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 15914 628634
rect 15294 592954 15914 628398
rect 15294 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 15914 592954
rect 15294 592634 15914 592718
rect 15294 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 15914 592634
rect 15294 556954 15914 592398
rect 15294 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 15914 556954
rect 15294 556634 15914 556718
rect 15294 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 15914 556634
rect 15294 520954 15914 556398
rect 15294 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 15914 520954
rect 15294 520634 15914 520718
rect 15294 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 15914 520634
rect 15294 484954 15914 520398
rect 15294 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 15914 484954
rect 15294 484634 15914 484718
rect 15294 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 15914 484634
rect 15294 448954 15914 484398
rect 15294 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 15914 448954
rect 15294 448634 15914 448718
rect 15294 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 15914 448634
rect 15294 412954 15914 448398
rect 15294 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 15914 412954
rect 15294 412634 15914 412718
rect 15294 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 15914 412634
rect 15294 376954 15914 412398
rect 15294 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 15914 376954
rect 15294 376634 15914 376718
rect 15294 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 15914 376634
rect 15294 340954 15914 376398
rect 15294 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 15914 340954
rect 15294 340634 15914 340718
rect 15294 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 15914 340634
rect 15294 304954 15914 340398
rect 15294 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 15914 304954
rect 15294 304634 15914 304718
rect 15294 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 15914 304634
rect 15294 268954 15914 304398
rect 15294 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 15914 268954
rect 15294 268634 15914 268718
rect 15294 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 15914 268634
rect 15294 232954 15914 268398
rect 15294 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 15914 232954
rect 15294 232634 15914 232718
rect 15294 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 15914 232634
rect 15294 196954 15914 232398
rect 15294 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 15914 196954
rect 15294 196634 15914 196718
rect 15294 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 15914 196634
rect 15294 160954 15914 196398
rect 15294 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 15914 160954
rect 15294 160634 15914 160718
rect 15294 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 15914 160634
rect 15294 124954 15914 160398
rect 15294 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 15914 124954
rect 15294 124634 15914 124718
rect 15294 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 15914 124634
rect 15294 88954 15914 124398
rect 15294 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 15914 88954
rect 15294 88634 15914 88718
rect 15294 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 15914 88634
rect 15294 52954 15914 88398
rect 15294 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 15914 52954
rect 15294 52634 15914 52718
rect 15294 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 15914 52634
rect 15294 16954 15914 52398
rect 15294 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 15914 16954
rect 15294 16634 15914 16718
rect 15294 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 15914 16634
rect 15294 -3226 15914 16398
rect 15294 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 15914 -3226
rect 15294 -3546 15914 -3462
rect 15294 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 15914 -3546
rect 15294 -7654 15914 -3782
rect 19794 708678 20414 711590
rect 19794 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 20414 708678
rect 19794 708358 20414 708442
rect 19794 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 20414 708358
rect 19794 669454 20414 708122
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -4186 20414 20898
rect 19794 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 20414 -4186
rect 19794 -4506 20414 -4422
rect 19794 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 20414 -4506
rect 19794 -7654 20414 -4742
rect 24294 709638 24914 711590
rect 24294 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 24914 709638
rect 24294 709318 24914 709402
rect 24294 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 24914 709318
rect 24294 673954 24914 709082
rect 24294 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 24914 673954
rect 24294 673634 24914 673718
rect 24294 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 24914 673634
rect 24294 637954 24914 673398
rect 24294 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 24914 637954
rect 24294 637634 24914 637718
rect 24294 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 24914 637634
rect 24294 601954 24914 637398
rect 24294 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 24914 601954
rect 24294 601634 24914 601718
rect 24294 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 24914 601634
rect 24294 565954 24914 601398
rect 24294 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 24914 565954
rect 24294 565634 24914 565718
rect 24294 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 24914 565634
rect 24294 529954 24914 565398
rect 24294 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 24914 529954
rect 24294 529634 24914 529718
rect 24294 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 24914 529634
rect 24294 493954 24914 529398
rect 24294 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 24914 493954
rect 24294 493634 24914 493718
rect 24294 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 24914 493634
rect 24294 457954 24914 493398
rect 24294 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 24914 457954
rect 24294 457634 24914 457718
rect 24294 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 24914 457634
rect 24294 421954 24914 457398
rect 24294 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 24914 421954
rect 24294 421634 24914 421718
rect 24294 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 24914 421634
rect 24294 385954 24914 421398
rect 24294 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 24914 385954
rect 24294 385634 24914 385718
rect 24294 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 24914 385634
rect 24294 349954 24914 385398
rect 24294 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 24914 349954
rect 24294 349634 24914 349718
rect 24294 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 24914 349634
rect 24294 313954 24914 349398
rect 24294 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 24914 313954
rect 24294 313634 24914 313718
rect 24294 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 24914 313634
rect 24294 277954 24914 313398
rect 24294 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 24914 277954
rect 24294 277634 24914 277718
rect 24294 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 24914 277634
rect 24294 241954 24914 277398
rect 24294 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 24914 241954
rect 24294 241634 24914 241718
rect 24294 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 24914 241634
rect 24294 205954 24914 241398
rect 24294 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 24914 205954
rect 24294 205634 24914 205718
rect 24294 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 24914 205634
rect 24294 169954 24914 205398
rect 24294 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 24914 169954
rect 24294 169634 24914 169718
rect 24294 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 24914 169634
rect 24294 133954 24914 169398
rect 24294 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 24914 133954
rect 24294 133634 24914 133718
rect 24294 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 24914 133634
rect 24294 97954 24914 133398
rect 24294 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 24914 97954
rect 24294 97634 24914 97718
rect 24294 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 24914 97634
rect 24294 61954 24914 97398
rect 24294 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 24914 61954
rect 24294 61634 24914 61718
rect 24294 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 24914 61634
rect 24294 25954 24914 61398
rect 24294 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 24914 25954
rect 24294 25634 24914 25718
rect 24294 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 24914 25634
rect 24294 -5146 24914 25398
rect 24294 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 24914 -5146
rect 24294 -5466 24914 -5382
rect 24294 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 24914 -5466
rect 24294 -7654 24914 -5702
rect 28794 710598 29414 711590
rect 28794 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 29414 710598
rect 28794 710278 29414 710362
rect 28794 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 29414 710278
rect 28794 678454 29414 710042
rect 28794 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 29414 678454
rect 28794 678134 29414 678218
rect 28794 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 29414 678134
rect 28794 642454 29414 677898
rect 28794 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 29414 642454
rect 28794 642134 29414 642218
rect 28794 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 29414 642134
rect 28794 606454 29414 641898
rect 28794 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 29414 606454
rect 28794 606134 29414 606218
rect 28794 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 29414 606134
rect 28794 570454 29414 605898
rect 28794 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 29414 570454
rect 28794 570134 29414 570218
rect 28794 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 29414 570134
rect 28794 534454 29414 569898
rect 28794 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 29414 534454
rect 28794 534134 29414 534218
rect 28794 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 29414 534134
rect 28794 498454 29414 533898
rect 28794 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 29414 498454
rect 28794 498134 29414 498218
rect 28794 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 29414 498134
rect 28794 462454 29414 497898
rect 28794 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 29414 462454
rect 28794 462134 29414 462218
rect 28794 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 29414 462134
rect 28794 426454 29414 461898
rect 28794 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 29414 426454
rect 28794 426134 29414 426218
rect 28794 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 29414 426134
rect 28794 390454 29414 425898
rect 28794 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 29414 390454
rect 28794 390134 29414 390218
rect 28794 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 29414 390134
rect 28794 354454 29414 389898
rect 28794 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 29414 354454
rect 28794 354134 29414 354218
rect 28794 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 29414 354134
rect 28794 318454 29414 353898
rect 28794 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 29414 318454
rect 28794 318134 29414 318218
rect 28794 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 29414 318134
rect 28794 282454 29414 317898
rect 28794 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 29414 282454
rect 28794 282134 29414 282218
rect 28794 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 29414 282134
rect 28794 246454 29414 281898
rect 28794 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 29414 246454
rect 28794 246134 29414 246218
rect 28794 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 29414 246134
rect 28794 210454 29414 245898
rect 28794 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 29414 210454
rect 28794 210134 29414 210218
rect 28794 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 29414 210134
rect 28794 174454 29414 209898
rect 28794 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 29414 174454
rect 28794 174134 29414 174218
rect 28794 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 29414 174134
rect 28794 138454 29414 173898
rect 28794 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 29414 138454
rect 28794 138134 29414 138218
rect 28794 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 29414 138134
rect 28794 102454 29414 137898
rect 28794 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 29414 102454
rect 28794 102134 29414 102218
rect 28794 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 29414 102134
rect 28794 66454 29414 101898
rect 28794 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 29414 66454
rect 28794 66134 29414 66218
rect 28794 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 29414 66134
rect 28794 30454 29414 65898
rect 28794 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 29414 30454
rect 28794 30134 29414 30218
rect 28794 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 29414 30134
rect 28794 -6106 29414 29898
rect 28794 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 29414 -6106
rect 28794 -6426 29414 -6342
rect 28794 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 29414 -6426
rect 28794 -7654 29414 -6662
rect 33294 711558 33914 711590
rect 33294 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 33914 711558
rect 33294 711238 33914 711322
rect 33294 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 33914 711238
rect 33294 682954 33914 711002
rect 33294 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 33914 682954
rect 33294 682634 33914 682718
rect 33294 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 33914 682634
rect 33294 646954 33914 682398
rect 33294 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 33914 646954
rect 33294 646634 33914 646718
rect 33294 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 33914 646634
rect 33294 610954 33914 646398
rect 33294 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 33914 610954
rect 33294 610634 33914 610718
rect 33294 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 33914 610634
rect 33294 574954 33914 610398
rect 33294 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 33914 574954
rect 33294 574634 33914 574718
rect 33294 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 33914 574634
rect 33294 538954 33914 574398
rect 33294 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 33914 538954
rect 33294 538634 33914 538718
rect 33294 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 33914 538634
rect 33294 502954 33914 538398
rect 33294 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 33914 502954
rect 33294 502634 33914 502718
rect 33294 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 33914 502634
rect 33294 466954 33914 502398
rect 33294 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 33914 466954
rect 33294 466634 33914 466718
rect 33294 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 33914 466634
rect 33294 430954 33914 466398
rect 33294 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 33914 430954
rect 33294 430634 33914 430718
rect 33294 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 33914 430634
rect 33294 394954 33914 430398
rect 33294 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 33914 394954
rect 33294 394634 33914 394718
rect 33294 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 33914 394634
rect 33294 358954 33914 394398
rect 33294 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 33914 358954
rect 33294 358634 33914 358718
rect 33294 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 33914 358634
rect 33294 322954 33914 358398
rect 33294 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 33914 322954
rect 33294 322634 33914 322718
rect 33294 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 33914 322634
rect 33294 286954 33914 322398
rect 33294 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 33914 286954
rect 33294 286634 33914 286718
rect 33294 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 33914 286634
rect 33294 250954 33914 286398
rect 33294 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 33914 250954
rect 33294 250634 33914 250718
rect 33294 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 33914 250634
rect 33294 214954 33914 250398
rect 33294 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 33914 214954
rect 33294 214634 33914 214718
rect 33294 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 33914 214634
rect 33294 178954 33914 214398
rect 33294 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 33914 178954
rect 33294 178634 33914 178718
rect 33294 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 33914 178634
rect 33294 142954 33914 178398
rect 33294 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 33914 142954
rect 33294 142634 33914 142718
rect 33294 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 33914 142634
rect 33294 106954 33914 142398
rect 33294 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 33914 106954
rect 33294 106634 33914 106718
rect 33294 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 33914 106634
rect 33294 70954 33914 106398
rect 33294 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 33914 70954
rect 33294 70634 33914 70718
rect 33294 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 33914 70634
rect 33294 34954 33914 70398
rect 33294 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 33914 34954
rect 33294 34634 33914 34718
rect 33294 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 33914 34634
rect 33294 -7066 33914 34398
rect 33294 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 33914 -7066
rect 33294 -7386 33914 -7302
rect 33294 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 33914 -7386
rect 33294 -7654 33914 -7622
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 42294 705798 42914 711590
rect 42294 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 42914 705798
rect 42294 705478 42914 705562
rect 42294 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 42914 705478
rect 42294 691954 42914 705242
rect 42294 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 42914 691954
rect 42294 691634 42914 691718
rect 42294 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 42914 691634
rect 42294 655954 42914 691398
rect 42294 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 42914 655954
rect 42294 655634 42914 655718
rect 42294 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 42914 655634
rect 42294 619954 42914 655398
rect 42294 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 42914 619954
rect 42294 619634 42914 619718
rect 42294 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 42914 619634
rect 42294 583954 42914 619398
rect 42294 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 42914 583954
rect 42294 583634 42914 583718
rect 42294 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 42914 583634
rect 42294 547954 42914 583398
rect 42294 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 42914 547954
rect 42294 547634 42914 547718
rect 42294 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 42914 547634
rect 42294 511954 42914 547398
rect 42294 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 42914 511954
rect 42294 511634 42914 511718
rect 42294 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 42914 511634
rect 42294 475954 42914 511398
rect 42294 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 42914 475954
rect 42294 475634 42914 475718
rect 42294 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 42914 475634
rect 42294 439954 42914 475398
rect 42294 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 42914 439954
rect 42294 439634 42914 439718
rect 42294 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 42914 439634
rect 42294 403954 42914 439398
rect 42294 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 42914 403954
rect 42294 403634 42914 403718
rect 42294 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 42914 403634
rect 42294 367954 42914 403398
rect 42294 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 42914 367954
rect 42294 367634 42914 367718
rect 42294 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 42914 367634
rect 42294 331954 42914 367398
rect 42294 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 42914 331954
rect 42294 331634 42914 331718
rect 42294 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 42914 331634
rect 42294 295954 42914 331398
rect 42294 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 42914 295954
rect 42294 295634 42914 295718
rect 42294 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 42914 295634
rect 42294 259954 42914 295398
rect 42294 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 42914 259954
rect 42294 259634 42914 259718
rect 42294 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 42914 259634
rect 42294 223954 42914 259398
rect 46794 706758 47414 711590
rect 46794 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 47414 706758
rect 46794 706438 47414 706522
rect 46794 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 47414 706438
rect 46794 696454 47414 706202
rect 46794 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 47414 696454
rect 46794 696134 47414 696218
rect 46794 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 47414 696134
rect 46794 660454 47414 695898
rect 46794 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 47414 660454
rect 46794 660134 47414 660218
rect 46794 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 47414 660134
rect 46794 624454 47414 659898
rect 46794 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 47414 624454
rect 46794 624134 47414 624218
rect 46794 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 47414 624134
rect 46794 588454 47414 623898
rect 46794 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 47414 588454
rect 46794 588134 47414 588218
rect 46794 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 47414 588134
rect 46794 552454 47414 587898
rect 46794 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 47414 552454
rect 46794 552134 47414 552218
rect 46794 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 47414 552134
rect 46794 516454 47414 551898
rect 46794 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 47414 516454
rect 46794 516134 47414 516218
rect 46794 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 47414 516134
rect 46794 480454 47414 515898
rect 46794 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 47414 480454
rect 46794 480134 47414 480218
rect 46794 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 47414 480134
rect 46794 444454 47414 479898
rect 46794 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 47414 444454
rect 46794 444134 47414 444218
rect 46794 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 47414 444134
rect 46794 408454 47414 443898
rect 46794 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 47414 408454
rect 46794 408134 47414 408218
rect 46794 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 47414 408134
rect 46794 372454 47414 407898
rect 46794 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 47414 372454
rect 46794 372134 47414 372218
rect 46794 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 47414 372134
rect 46794 336454 47414 371898
rect 46794 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 47414 336454
rect 46794 336134 47414 336218
rect 46794 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 47414 336134
rect 46794 300454 47414 335898
rect 46794 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 47414 300454
rect 46794 300134 47414 300218
rect 46794 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 47414 300134
rect 46794 264454 47414 299898
rect 46794 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 47414 264454
rect 46794 264134 47414 264218
rect 46794 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 47414 264134
rect 46794 248684 47414 263898
rect 51294 707718 51914 711590
rect 51294 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 51914 707718
rect 51294 707398 51914 707482
rect 51294 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 51914 707398
rect 51294 700954 51914 707162
rect 51294 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 51914 700954
rect 51294 700634 51914 700718
rect 51294 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 51914 700634
rect 51294 664954 51914 700398
rect 51294 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 51914 664954
rect 51294 664634 51914 664718
rect 51294 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 51914 664634
rect 51294 628954 51914 664398
rect 51294 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 51914 628954
rect 51294 628634 51914 628718
rect 51294 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 51914 628634
rect 51294 592954 51914 628398
rect 51294 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 51914 592954
rect 51294 592634 51914 592718
rect 51294 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 51914 592634
rect 51294 556954 51914 592398
rect 51294 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 51914 556954
rect 51294 556634 51914 556718
rect 51294 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 51914 556634
rect 51294 520954 51914 556398
rect 51294 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 51914 520954
rect 51294 520634 51914 520718
rect 51294 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 51914 520634
rect 51294 484954 51914 520398
rect 51294 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 51914 484954
rect 51294 484634 51914 484718
rect 51294 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 51914 484634
rect 51294 448954 51914 484398
rect 51294 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 51914 448954
rect 51294 448634 51914 448718
rect 51294 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 51914 448634
rect 51294 412954 51914 448398
rect 51294 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 51914 412954
rect 51294 412634 51914 412718
rect 51294 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 51914 412634
rect 51294 376954 51914 412398
rect 51294 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 51914 376954
rect 51294 376634 51914 376718
rect 51294 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 51914 376634
rect 51294 340954 51914 376398
rect 51294 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 51914 340954
rect 51294 340634 51914 340718
rect 51294 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 51914 340634
rect 51294 304954 51914 340398
rect 51294 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 51914 304954
rect 51294 304634 51914 304718
rect 51294 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 51914 304634
rect 51294 268954 51914 304398
rect 51294 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 51914 268954
rect 51294 268634 51914 268718
rect 51294 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 51914 268634
rect 51294 248684 51914 268398
rect 55794 708678 56414 711590
rect 55794 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 56414 708678
rect 55794 708358 56414 708442
rect 55794 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 56414 708358
rect 55794 669454 56414 708122
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 248684 56414 272898
rect 60294 709638 60914 711590
rect 60294 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 60914 709638
rect 60294 709318 60914 709402
rect 60294 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 60914 709318
rect 60294 673954 60914 709082
rect 60294 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 60914 673954
rect 60294 673634 60914 673718
rect 60294 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 60914 673634
rect 60294 637954 60914 673398
rect 60294 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 60914 637954
rect 60294 637634 60914 637718
rect 60294 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 60914 637634
rect 60294 601954 60914 637398
rect 60294 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 60914 601954
rect 60294 601634 60914 601718
rect 60294 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 60914 601634
rect 60294 565954 60914 601398
rect 60294 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 60914 565954
rect 60294 565634 60914 565718
rect 60294 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 60914 565634
rect 60294 529954 60914 565398
rect 60294 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 60914 529954
rect 60294 529634 60914 529718
rect 60294 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 60914 529634
rect 60294 493954 60914 529398
rect 60294 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 60914 493954
rect 60294 493634 60914 493718
rect 60294 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 60914 493634
rect 60294 457954 60914 493398
rect 60294 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 60914 457954
rect 60294 457634 60914 457718
rect 60294 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 60914 457634
rect 60294 421954 60914 457398
rect 60294 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 60914 421954
rect 60294 421634 60914 421718
rect 60294 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 60914 421634
rect 60294 385954 60914 421398
rect 60294 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 60914 385954
rect 60294 385634 60914 385718
rect 60294 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 60914 385634
rect 60294 349954 60914 385398
rect 60294 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 60914 349954
rect 60294 349634 60914 349718
rect 60294 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 60914 349634
rect 60294 313954 60914 349398
rect 60294 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 60914 313954
rect 60294 313634 60914 313718
rect 60294 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 60914 313634
rect 60294 277954 60914 313398
rect 60294 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 60914 277954
rect 60294 277634 60914 277718
rect 60294 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 60914 277634
rect 60294 248684 60914 277398
rect 64794 710598 65414 711590
rect 64794 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 65414 710598
rect 64794 710278 65414 710362
rect 64794 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 65414 710278
rect 64794 678454 65414 710042
rect 64794 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 65414 678454
rect 64794 678134 65414 678218
rect 64794 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 65414 678134
rect 64794 642454 65414 677898
rect 64794 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 65414 642454
rect 64794 642134 65414 642218
rect 64794 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 65414 642134
rect 64794 606454 65414 641898
rect 64794 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 65414 606454
rect 64794 606134 65414 606218
rect 64794 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 65414 606134
rect 64794 570454 65414 605898
rect 64794 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 65414 570454
rect 64794 570134 65414 570218
rect 64794 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 65414 570134
rect 64794 534454 65414 569898
rect 64794 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 65414 534454
rect 64794 534134 65414 534218
rect 64794 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 65414 534134
rect 64794 498454 65414 533898
rect 64794 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 65414 498454
rect 64794 498134 65414 498218
rect 64794 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 65414 498134
rect 64794 462454 65414 497898
rect 64794 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 65414 462454
rect 64794 462134 65414 462218
rect 64794 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 65414 462134
rect 64794 426454 65414 461898
rect 64794 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 65414 426454
rect 64794 426134 65414 426218
rect 64794 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 65414 426134
rect 64794 390454 65414 425898
rect 64794 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 65414 390454
rect 64794 390134 65414 390218
rect 64794 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 65414 390134
rect 64794 354454 65414 389898
rect 64794 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 65414 354454
rect 64794 354134 65414 354218
rect 64794 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 65414 354134
rect 64794 318454 65414 353898
rect 64794 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 65414 318454
rect 64794 318134 65414 318218
rect 64794 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 65414 318134
rect 64794 282454 65414 317898
rect 64794 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 65414 282454
rect 64794 282134 65414 282218
rect 64794 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 65414 282134
rect 64794 248684 65414 281898
rect 69294 711558 69914 711590
rect 69294 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 69914 711558
rect 69294 711238 69914 711322
rect 69294 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 69914 711238
rect 69294 682954 69914 711002
rect 69294 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 69914 682954
rect 69294 682634 69914 682718
rect 69294 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 69914 682634
rect 69294 646954 69914 682398
rect 69294 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 69914 646954
rect 69294 646634 69914 646718
rect 69294 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 69914 646634
rect 69294 610954 69914 646398
rect 69294 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 69914 610954
rect 69294 610634 69914 610718
rect 69294 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 69914 610634
rect 69294 574954 69914 610398
rect 69294 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 69914 574954
rect 69294 574634 69914 574718
rect 69294 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 69914 574634
rect 69294 538954 69914 574398
rect 69294 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 69914 538954
rect 69294 538634 69914 538718
rect 69294 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 69914 538634
rect 69294 502954 69914 538398
rect 69294 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 69914 502954
rect 69294 502634 69914 502718
rect 69294 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 69914 502634
rect 69294 466954 69914 502398
rect 69294 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 69914 466954
rect 69294 466634 69914 466718
rect 69294 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 69914 466634
rect 69294 430954 69914 466398
rect 69294 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 69914 430954
rect 69294 430634 69914 430718
rect 69294 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 69914 430634
rect 69294 394954 69914 430398
rect 69294 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 69914 394954
rect 69294 394634 69914 394718
rect 69294 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 69914 394634
rect 69294 358954 69914 394398
rect 69294 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 69914 358954
rect 69294 358634 69914 358718
rect 69294 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 69914 358634
rect 69294 322954 69914 358398
rect 69294 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 69914 322954
rect 69294 322634 69914 322718
rect 69294 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 69914 322634
rect 69294 286954 69914 322398
rect 69294 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 69914 286954
rect 69294 286634 69914 286718
rect 69294 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 69914 286634
rect 69294 250954 69914 286398
rect 69294 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 69914 250954
rect 69294 250634 69914 250718
rect 69294 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 69914 250634
rect 69294 248684 69914 250398
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 248684 74414 254898
rect 78294 705798 78914 711590
rect 78294 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 78914 705798
rect 78294 705478 78914 705562
rect 78294 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 78914 705478
rect 78294 691954 78914 705242
rect 78294 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 78914 691954
rect 78294 691634 78914 691718
rect 78294 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 78914 691634
rect 78294 655954 78914 691398
rect 78294 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 78914 655954
rect 78294 655634 78914 655718
rect 78294 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 78914 655634
rect 78294 619954 78914 655398
rect 78294 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 78914 619954
rect 78294 619634 78914 619718
rect 78294 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 78914 619634
rect 78294 583954 78914 619398
rect 78294 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 78914 583954
rect 78294 583634 78914 583718
rect 78294 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 78914 583634
rect 78294 547954 78914 583398
rect 78294 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 78914 547954
rect 78294 547634 78914 547718
rect 78294 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 78914 547634
rect 78294 511954 78914 547398
rect 78294 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 78914 511954
rect 78294 511634 78914 511718
rect 78294 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 78914 511634
rect 78294 475954 78914 511398
rect 78294 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 78914 475954
rect 78294 475634 78914 475718
rect 78294 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 78914 475634
rect 78294 439954 78914 475398
rect 78294 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 78914 439954
rect 78294 439634 78914 439718
rect 78294 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 78914 439634
rect 78294 403954 78914 439398
rect 78294 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 78914 403954
rect 78294 403634 78914 403718
rect 78294 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 78914 403634
rect 78294 367954 78914 403398
rect 78294 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 78914 367954
rect 78294 367634 78914 367718
rect 78294 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 78914 367634
rect 78294 331954 78914 367398
rect 78294 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 78914 331954
rect 78294 331634 78914 331718
rect 78294 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 78914 331634
rect 78294 295954 78914 331398
rect 78294 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 78914 295954
rect 78294 295634 78914 295718
rect 78294 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 78914 295634
rect 78294 259954 78914 295398
rect 78294 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 78914 259954
rect 78294 259634 78914 259718
rect 78294 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 78914 259634
rect 78294 248684 78914 259398
rect 82794 706758 83414 711590
rect 82794 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 83414 706758
rect 82794 706438 83414 706522
rect 82794 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 83414 706438
rect 82794 696454 83414 706202
rect 82794 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 83414 696454
rect 82794 696134 83414 696218
rect 82794 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 83414 696134
rect 82794 660454 83414 695898
rect 82794 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 83414 660454
rect 82794 660134 83414 660218
rect 82794 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 83414 660134
rect 82794 624454 83414 659898
rect 82794 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 83414 624454
rect 82794 624134 83414 624218
rect 82794 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 83414 624134
rect 82794 588454 83414 623898
rect 82794 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 83414 588454
rect 82794 588134 83414 588218
rect 82794 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 83414 588134
rect 82794 552454 83414 587898
rect 82794 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 83414 552454
rect 82794 552134 83414 552218
rect 82794 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 83414 552134
rect 82794 516454 83414 551898
rect 82794 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 83414 516454
rect 82794 516134 83414 516218
rect 82794 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 83414 516134
rect 82794 480454 83414 515898
rect 82794 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 83414 480454
rect 82794 480134 83414 480218
rect 82794 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 83414 480134
rect 82794 444454 83414 479898
rect 82794 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 83414 444454
rect 82794 444134 83414 444218
rect 82794 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 83414 444134
rect 82794 408454 83414 443898
rect 82794 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 83414 408454
rect 82794 408134 83414 408218
rect 82794 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 83414 408134
rect 82794 372454 83414 407898
rect 82794 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 83414 372454
rect 82794 372134 83414 372218
rect 82794 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 83414 372134
rect 82794 336454 83414 371898
rect 82794 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 83414 336454
rect 82794 336134 83414 336218
rect 82794 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 83414 336134
rect 82794 300454 83414 335898
rect 82794 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 83414 300454
rect 82794 300134 83414 300218
rect 82794 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 83414 300134
rect 82794 264454 83414 299898
rect 82794 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 83414 264454
rect 82794 264134 83414 264218
rect 82794 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 83414 264134
rect 82794 248684 83414 263898
rect 87294 707718 87914 711590
rect 87294 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 87914 707718
rect 87294 707398 87914 707482
rect 87294 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 87914 707398
rect 87294 700954 87914 707162
rect 87294 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 87914 700954
rect 87294 700634 87914 700718
rect 87294 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 87914 700634
rect 87294 664954 87914 700398
rect 87294 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 87914 664954
rect 87294 664634 87914 664718
rect 87294 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 87914 664634
rect 87294 628954 87914 664398
rect 87294 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 87914 628954
rect 87294 628634 87914 628718
rect 87294 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 87914 628634
rect 87294 592954 87914 628398
rect 87294 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 87914 592954
rect 87294 592634 87914 592718
rect 87294 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 87914 592634
rect 87294 556954 87914 592398
rect 87294 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 87914 556954
rect 87294 556634 87914 556718
rect 87294 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 87914 556634
rect 87294 520954 87914 556398
rect 87294 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 87914 520954
rect 87294 520634 87914 520718
rect 87294 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 87914 520634
rect 87294 484954 87914 520398
rect 87294 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 87914 484954
rect 87294 484634 87914 484718
rect 87294 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 87914 484634
rect 87294 448954 87914 484398
rect 87294 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 87914 448954
rect 87294 448634 87914 448718
rect 87294 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 87914 448634
rect 87294 412954 87914 448398
rect 87294 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 87914 412954
rect 87294 412634 87914 412718
rect 87294 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 87914 412634
rect 87294 376954 87914 412398
rect 87294 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 87914 376954
rect 87294 376634 87914 376718
rect 87294 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 87914 376634
rect 87294 340954 87914 376398
rect 87294 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 87914 340954
rect 87294 340634 87914 340718
rect 87294 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 87914 340634
rect 87294 304954 87914 340398
rect 87294 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 87914 304954
rect 87294 304634 87914 304718
rect 87294 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 87914 304634
rect 87294 268954 87914 304398
rect 87294 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 87914 268954
rect 87294 268634 87914 268718
rect 87294 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 87914 268634
rect 87294 248684 87914 268398
rect 91794 708678 92414 711590
rect 91794 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 92414 708678
rect 91794 708358 92414 708442
rect 91794 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 92414 708358
rect 91794 669454 92414 708122
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 273454 92414 308898
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 248684 92414 272898
rect 96294 709638 96914 711590
rect 96294 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 96914 709638
rect 96294 709318 96914 709402
rect 96294 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 96914 709318
rect 96294 673954 96914 709082
rect 96294 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 96914 673954
rect 96294 673634 96914 673718
rect 96294 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 96914 673634
rect 96294 637954 96914 673398
rect 96294 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 96914 637954
rect 96294 637634 96914 637718
rect 96294 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 96914 637634
rect 96294 601954 96914 637398
rect 96294 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 96914 601954
rect 96294 601634 96914 601718
rect 96294 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 96914 601634
rect 96294 565954 96914 601398
rect 96294 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 96914 565954
rect 96294 565634 96914 565718
rect 96294 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 96914 565634
rect 96294 529954 96914 565398
rect 96294 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 96914 529954
rect 96294 529634 96914 529718
rect 96294 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 96914 529634
rect 96294 493954 96914 529398
rect 96294 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 96914 493954
rect 96294 493634 96914 493718
rect 96294 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 96914 493634
rect 96294 457954 96914 493398
rect 96294 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 96914 457954
rect 96294 457634 96914 457718
rect 96294 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 96914 457634
rect 96294 421954 96914 457398
rect 96294 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 96914 421954
rect 96294 421634 96914 421718
rect 96294 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 96914 421634
rect 96294 385954 96914 421398
rect 96294 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 96914 385954
rect 96294 385634 96914 385718
rect 96294 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 96914 385634
rect 96294 349954 96914 385398
rect 96294 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 96914 349954
rect 96294 349634 96914 349718
rect 96294 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 96914 349634
rect 96294 313954 96914 349398
rect 96294 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 96914 313954
rect 96294 313634 96914 313718
rect 96294 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 96914 313634
rect 96294 277954 96914 313398
rect 96294 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 96914 277954
rect 96294 277634 96914 277718
rect 96294 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 96914 277634
rect 96294 248684 96914 277398
rect 100794 710598 101414 711590
rect 100794 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 101414 710598
rect 100794 710278 101414 710362
rect 100794 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 101414 710278
rect 100794 678454 101414 710042
rect 100794 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 101414 678454
rect 100794 678134 101414 678218
rect 100794 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 101414 678134
rect 100794 642454 101414 677898
rect 100794 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 101414 642454
rect 100794 642134 101414 642218
rect 100794 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 101414 642134
rect 100794 606454 101414 641898
rect 100794 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 101414 606454
rect 100794 606134 101414 606218
rect 100794 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 101414 606134
rect 100794 570454 101414 605898
rect 100794 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 101414 570454
rect 100794 570134 101414 570218
rect 100794 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 101414 570134
rect 100794 534454 101414 569898
rect 100794 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 101414 534454
rect 100794 534134 101414 534218
rect 100794 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 101414 534134
rect 100794 498454 101414 533898
rect 100794 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 101414 498454
rect 100794 498134 101414 498218
rect 100794 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 101414 498134
rect 100794 462454 101414 497898
rect 100794 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 101414 462454
rect 100794 462134 101414 462218
rect 100794 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 101414 462134
rect 100794 426454 101414 461898
rect 100794 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 101414 426454
rect 100794 426134 101414 426218
rect 100794 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 101414 426134
rect 100794 390454 101414 425898
rect 100794 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 101414 390454
rect 100794 390134 101414 390218
rect 100794 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 101414 390134
rect 100794 354454 101414 389898
rect 100794 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 101414 354454
rect 100794 354134 101414 354218
rect 100794 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 101414 354134
rect 100794 318454 101414 353898
rect 100794 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 101414 318454
rect 100794 318134 101414 318218
rect 100794 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 101414 318134
rect 100794 282454 101414 317898
rect 100794 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 101414 282454
rect 100794 282134 101414 282218
rect 100794 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 101414 282134
rect 100794 248684 101414 281898
rect 105294 711558 105914 711590
rect 105294 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 105914 711558
rect 105294 711238 105914 711322
rect 105294 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 105914 711238
rect 105294 682954 105914 711002
rect 105294 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 105914 682954
rect 105294 682634 105914 682718
rect 105294 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 105914 682634
rect 105294 646954 105914 682398
rect 105294 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 105914 646954
rect 105294 646634 105914 646718
rect 105294 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 105914 646634
rect 105294 610954 105914 646398
rect 105294 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 105914 610954
rect 105294 610634 105914 610718
rect 105294 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 105914 610634
rect 105294 574954 105914 610398
rect 105294 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 105914 574954
rect 105294 574634 105914 574718
rect 105294 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 105914 574634
rect 105294 538954 105914 574398
rect 105294 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 105914 538954
rect 105294 538634 105914 538718
rect 105294 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 105914 538634
rect 105294 502954 105914 538398
rect 105294 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 105914 502954
rect 105294 502634 105914 502718
rect 105294 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 105914 502634
rect 105294 466954 105914 502398
rect 105294 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 105914 466954
rect 105294 466634 105914 466718
rect 105294 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 105914 466634
rect 105294 430954 105914 466398
rect 105294 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 105914 430954
rect 105294 430634 105914 430718
rect 105294 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 105914 430634
rect 105294 394954 105914 430398
rect 105294 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 105914 394954
rect 105294 394634 105914 394718
rect 105294 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 105914 394634
rect 105294 358954 105914 394398
rect 105294 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 105914 358954
rect 105294 358634 105914 358718
rect 105294 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 105914 358634
rect 105294 322954 105914 358398
rect 105294 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 105914 322954
rect 105294 322634 105914 322718
rect 105294 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 105914 322634
rect 105294 286954 105914 322398
rect 105294 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 105914 286954
rect 105294 286634 105914 286718
rect 105294 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 105914 286634
rect 105294 250954 105914 286398
rect 105294 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 105914 250954
rect 105294 250634 105914 250718
rect 105294 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 105914 250634
rect 105294 248684 105914 250398
rect 109794 704838 110414 711590
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 248684 110414 254898
rect 114294 705798 114914 711590
rect 114294 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 114914 705798
rect 114294 705478 114914 705562
rect 114294 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 114914 705478
rect 114294 691954 114914 705242
rect 114294 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 114914 691954
rect 114294 691634 114914 691718
rect 114294 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 114914 691634
rect 114294 655954 114914 691398
rect 114294 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 114914 655954
rect 114294 655634 114914 655718
rect 114294 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 114914 655634
rect 114294 619954 114914 655398
rect 114294 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 114914 619954
rect 114294 619634 114914 619718
rect 114294 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 114914 619634
rect 114294 583954 114914 619398
rect 114294 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 114914 583954
rect 114294 583634 114914 583718
rect 114294 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 114914 583634
rect 114294 547954 114914 583398
rect 114294 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 114914 547954
rect 114294 547634 114914 547718
rect 114294 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 114914 547634
rect 114294 511954 114914 547398
rect 114294 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 114914 511954
rect 114294 511634 114914 511718
rect 114294 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 114914 511634
rect 114294 475954 114914 511398
rect 114294 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 114914 475954
rect 114294 475634 114914 475718
rect 114294 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 114914 475634
rect 114294 439954 114914 475398
rect 114294 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 114914 439954
rect 114294 439634 114914 439718
rect 114294 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 114914 439634
rect 114294 403954 114914 439398
rect 114294 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 114914 403954
rect 114294 403634 114914 403718
rect 114294 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 114914 403634
rect 114294 367954 114914 403398
rect 114294 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 114914 367954
rect 114294 367634 114914 367718
rect 114294 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 114914 367634
rect 114294 331954 114914 367398
rect 114294 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 114914 331954
rect 114294 331634 114914 331718
rect 114294 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 114914 331634
rect 114294 295954 114914 331398
rect 114294 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 114914 295954
rect 114294 295634 114914 295718
rect 114294 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 114914 295634
rect 114294 259954 114914 295398
rect 114294 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 114914 259954
rect 114294 259634 114914 259718
rect 114294 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 114914 259634
rect 114294 248684 114914 259398
rect 118794 706758 119414 711590
rect 118794 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 119414 706758
rect 118794 706438 119414 706522
rect 118794 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 119414 706438
rect 118794 696454 119414 706202
rect 118794 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 119414 696454
rect 118794 696134 119414 696218
rect 118794 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 119414 696134
rect 118794 660454 119414 695898
rect 118794 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 119414 660454
rect 118794 660134 119414 660218
rect 118794 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 119414 660134
rect 118794 624454 119414 659898
rect 118794 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 119414 624454
rect 118794 624134 119414 624218
rect 118794 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 119414 624134
rect 118794 588454 119414 623898
rect 118794 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 119414 588454
rect 118794 588134 119414 588218
rect 118794 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 119414 588134
rect 118794 552454 119414 587898
rect 118794 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 119414 552454
rect 118794 552134 119414 552218
rect 118794 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 119414 552134
rect 118794 516454 119414 551898
rect 118794 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 119414 516454
rect 118794 516134 119414 516218
rect 118794 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 119414 516134
rect 118794 480454 119414 515898
rect 118794 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 119414 480454
rect 118794 480134 119414 480218
rect 118794 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 119414 480134
rect 118794 444454 119414 479898
rect 118794 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 119414 444454
rect 118794 444134 119414 444218
rect 118794 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 119414 444134
rect 118794 408454 119414 443898
rect 118794 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 119414 408454
rect 118794 408134 119414 408218
rect 118794 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 119414 408134
rect 118794 372454 119414 407898
rect 118794 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 119414 372454
rect 118794 372134 119414 372218
rect 118794 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 119414 372134
rect 118794 336454 119414 371898
rect 118794 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 119414 336454
rect 118794 336134 119414 336218
rect 118794 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 119414 336134
rect 118794 300454 119414 335898
rect 118794 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 119414 300454
rect 118794 300134 119414 300218
rect 118794 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 119414 300134
rect 118794 264454 119414 299898
rect 118794 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 119414 264454
rect 118794 264134 119414 264218
rect 118794 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 119414 264134
rect 118794 248684 119414 263898
rect 123294 707718 123914 711590
rect 123294 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 123914 707718
rect 123294 707398 123914 707482
rect 123294 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 123914 707398
rect 123294 700954 123914 707162
rect 123294 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 123914 700954
rect 123294 700634 123914 700718
rect 123294 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 123914 700634
rect 123294 664954 123914 700398
rect 123294 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 123914 664954
rect 123294 664634 123914 664718
rect 123294 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 123914 664634
rect 123294 628954 123914 664398
rect 123294 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 123914 628954
rect 123294 628634 123914 628718
rect 123294 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 123914 628634
rect 123294 592954 123914 628398
rect 123294 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 123914 592954
rect 123294 592634 123914 592718
rect 123294 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 123914 592634
rect 123294 556954 123914 592398
rect 123294 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 123914 556954
rect 123294 556634 123914 556718
rect 123294 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 123914 556634
rect 123294 520954 123914 556398
rect 123294 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 123914 520954
rect 123294 520634 123914 520718
rect 123294 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 123914 520634
rect 123294 484954 123914 520398
rect 123294 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 123914 484954
rect 123294 484634 123914 484718
rect 123294 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 123914 484634
rect 123294 448954 123914 484398
rect 123294 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 123914 448954
rect 123294 448634 123914 448718
rect 123294 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 123914 448634
rect 123294 412954 123914 448398
rect 123294 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 123914 412954
rect 123294 412634 123914 412718
rect 123294 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 123914 412634
rect 123294 376954 123914 412398
rect 123294 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 123914 376954
rect 123294 376634 123914 376718
rect 123294 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 123914 376634
rect 123294 340954 123914 376398
rect 123294 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 123914 340954
rect 123294 340634 123914 340718
rect 123294 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 123914 340634
rect 123294 304954 123914 340398
rect 123294 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 123914 304954
rect 123294 304634 123914 304718
rect 123294 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 123914 304634
rect 123294 268954 123914 304398
rect 123294 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 123914 268954
rect 123294 268634 123914 268718
rect 123294 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 123914 268634
rect 123294 248684 123914 268398
rect 127794 708678 128414 711590
rect 127794 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 128414 708678
rect 127794 708358 128414 708442
rect 127794 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 128414 708358
rect 127794 669454 128414 708122
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 248684 128414 272898
rect 132294 709638 132914 711590
rect 132294 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 132914 709638
rect 132294 709318 132914 709402
rect 132294 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 132914 709318
rect 132294 673954 132914 709082
rect 132294 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 132914 673954
rect 132294 673634 132914 673718
rect 132294 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 132914 673634
rect 132294 637954 132914 673398
rect 132294 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 132914 637954
rect 132294 637634 132914 637718
rect 132294 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 132914 637634
rect 132294 601954 132914 637398
rect 132294 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 132914 601954
rect 132294 601634 132914 601718
rect 132294 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 132914 601634
rect 132294 565954 132914 601398
rect 132294 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 132914 565954
rect 132294 565634 132914 565718
rect 132294 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 132914 565634
rect 132294 529954 132914 565398
rect 132294 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 132914 529954
rect 132294 529634 132914 529718
rect 132294 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 132914 529634
rect 132294 493954 132914 529398
rect 132294 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 132914 493954
rect 132294 493634 132914 493718
rect 132294 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 132914 493634
rect 132294 457954 132914 493398
rect 132294 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 132914 457954
rect 132294 457634 132914 457718
rect 132294 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 132914 457634
rect 132294 421954 132914 457398
rect 132294 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 132914 421954
rect 132294 421634 132914 421718
rect 132294 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 132914 421634
rect 132294 385954 132914 421398
rect 132294 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 132914 385954
rect 132294 385634 132914 385718
rect 132294 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 132914 385634
rect 132294 349954 132914 385398
rect 132294 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 132914 349954
rect 132294 349634 132914 349718
rect 132294 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 132914 349634
rect 132294 313954 132914 349398
rect 132294 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 132914 313954
rect 132294 313634 132914 313718
rect 132294 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 132914 313634
rect 132294 277954 132914 313398
rect 132294 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 132914 277954
rect 132294 277634 132914 277718
rect 132294 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 132914 277634
rect 132294 248684 132914 277398
rect 136794 710598 137414 711590
rect 136794 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 137414 710598
rect 136794 710278 137414 710362
rect 136794 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 137414 710278
rect 136794 678454 137414 710042
rect 136794 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 137414 678454
rect 136794 678134 137414 678218
rect 136794 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 137414 678134
rect 136794 642454 137414 677898
rect 136794 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 137414 642454
rect 136794 642134 137414 642218
rect 136794 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 137414 642134
rect 136794 606454 137414 641898
rect 136794 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 137414 606454
rect 136794 606134 137414 606218
rect 136794 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 137414 606134
rect 136794 570454 137414 605898
rect 136794 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 137414 570454
rect 136794 570134 137414 570218
rect 136794 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 137414 570134
rect 136794 534454 137414 569898
rect 136794 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 137414 534454
rect 136794 534134 137414 534218
rect 136794 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 137414 534134
rect 136794 498454 137414 533898
rect 136794 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 137414 498454
rect 136794 498134 137414 498218
rect 136794 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 137414 498134
rect 136794 462454 137414 497898
rect 136794 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 137414 462454
rect 136794 462134 137414 462218
rect 136794 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 137414 462134
rect 136794 426454 137414 461898
rect 136794 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 137414 426454
rect 136794 426134 137414 426218
rect 136794 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 137414 426134
rect 136794 390454 137414 425898
rect 136794 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 137414 390454
rect 136794 390134 137414 390218
rect 136794 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 137414 390134
rect 136794 354454 137414 389898
rect 136794 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 137414 354454
rect 136794 354134 137414 354218
rect 136794 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 137414 354134
rect 136794 318454 137414 353898
rect 136794 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 137414 318454
rect 136794 318134 137414 318218
rect 136794 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 137414 318134
rect 136794 282454 137414 317898
rect 136794 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 137414 282454
rect 136794 282134 137414 282218
rect 136794 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 137414 282134
rect 136794 248684 137414 281898
rect 141294 711558 141914 711590
rect 141294 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 141914 711558
rect 141294 711238 141914 711322
rect 141294 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 141914 711238
rect 141294 682954 141914 711002
rect 141294 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 141914 682954
rect 141294 682634 141914 682718
rect 141294 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 141914 682634
rect 141294 646954 141914 682398
rect 141294 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 141914 646954
rect 141294 646634 141914 646718
rect 141294 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 141914 646634
rect 141294 610954 141914 646398
rect 141294 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 141914 610954
rect 141294 610634 141914 610718
rect 141294 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 141914 610634
rect 141294 574954 141914 610398
rect 141294 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 141914 574954
rect 141294 574634 141914 574718
rect 141294 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 141914 574634
rect 141294 538954 141914 574398
rect 141294 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 141914 538954
rect 141294 538634 141914 538718
rect 141294 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 141914 538634
rect 141294 502954 141914 538398
rect 141294 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 141914 502954
rect 141294 502634 141914 502718
rect 141294 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 141914 502634
rect 141294 466954 141914 502398
rect 141294 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 141914 466954
rect 141294 466634 141914 466718
rect 141294 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 141914 466634
rect 141294 430954 141914 466398
rect 141294 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 141914 430954
rect 141294 430634 141914 430718
rect 141294 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 141914 430634
rect 141294 394954 141914 430398
rect 141294 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 141914 394954
rect 141294 394634 141914 394718
rect 141294 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 141914 394634
rect 141294 358954 141914 394398
rect 141294 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 141914 358954
rect 141294 358634 141914 358718
rect 141294 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 141914 358634
rect 141294 322954 141914 358398
rect 141294 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 141914 322954
rect 141294 322634 141914 322718
rect 141294 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 141914 322634
rect 141294 286954 141914 322398
rect 141294 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 141914 286954
rect 141294 286634 141914 286718
rect 141294 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 141914 286634
rect 141294 250954 141914 286398
rect 141294 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 141914 250954
rect 141294 250634 141914 250718
rect 141294 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 141914 250634
rect 141294 248684 141914 250398
rect 145794 704838 146414 711590
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 248684 146414 254898
rect 150294 705798 150914 711590
rect 150294 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 150914 705798
rect 150294 705478 150914 705562
rect 150294 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 150914 705478
rect 150294 691954 150914 705242
rect 150294 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 150914 691954
rect 150294 691634 150914 691718
rect 150294 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 150914 691634
rect 150294 655954 150914 691398
rect 150294 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 150914 655954
rect 150294 655634 150914 655718
rect 150294 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 150914 655634
rect 150294 619954 150914 655398
rect 150294 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 150914 619954
rect 150294 619634 150914 619718
rect 150294 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 150914 619634
rect 150294 583954 150914 619398
rect 150294 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 150914 583954
rect 150294 583634 150914 583718
rect 150294 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 150914 583634
rect 150294 547954 150914 583398
rect 150294 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 150914 547954
rect 150294 547634 150914 547718
rect 150294 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 150914 547634
rect 150294 511954 150914 547398
rect 150294 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 150914 511954
rect 150294 511634 150914 511718
rect 150294 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 150914 511634
rect 150294 475954 150914 511398
rect 150294 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 150914 475954
rect 150294 475634 150914 475718
rect 150294 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 150914 475634
rect 150294 439954 150914 475398
rect 150294 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 150914 439954
rect 150294 439634 150914 439718
rect 150294 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 150914 439634
rect 150294 403954 150914 439398
rect 150294 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 150914 403954
rect 150294 403634 150914 403718
rect 150294 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 150914 403634
rect 150294 367954 150914 403398
rect 150294 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 150914 367954
rect 150294 367634 150914 367718
rect 150294 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 150914 367634
rect 150294 331954 150914 367398
rect 150294 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 150914 331954
rect 150294 331634 150914 331718
rect 150294 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 150914 331634
rect 150294 295954 150914 331398
rect 150294 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 150914 295954
rect 150294 295634 150914 295718
rect 150294 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 150914 295634
rect 150294 259954 150914 295398
rect 150294 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 150914 259954
rect 150294 259634 150914 259718
rect 150294 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 150914 259634
rect 150294 248684 150914 259398
rect 154794 706758 155414 711590
rect 154794 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 155414 706758
rect 154794 706438 155414 706522
rect 154794 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 155414 706438
rect 154794 696454 155414 706202
rect 154794 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 155414 696454
rect 154794 696134 155414 696218
rect 154794 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 155414 696134
rect 154794 660454 155414 695898
rect 154794 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 155414 660454
rect 154794 660134 155414 660218
rect 154794 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 155414 660134
rect 154794 624454 155414 659898
rect 154794 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 155414 624454
rect 154794 624134 155414 624218
rect 154794 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 155414 624134
rect 154794 588454 155414 623898
rect 154794 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 155414 588454
rect 154794 588134 155414 588218
rect 154794 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 155414 588134
rect 154794 552454 155414 587898
rect 154794 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 155414 552454
rect 154794 552134 155414 552218
rect 154794 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 155414 552134
rect 154794 516454 155414 551898
rect 154794 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 155414 516454
rect 154794 516134 155414 516218
rect 154794 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 155414 516134
rect 154794 480454 155414 515898
rect 154794 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 155414 480454
rect 154794 480134 155414 480218
rect 154794 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 155414 480134
rect 154794 444454 155414 479898
rect 154794 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 155414 444454
rect 154794 444134 155414 444218
rect 154794 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 155414 444134
rect 154794 408454 155414 443898
rect 154794 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 155414 408454
rect 154794 408134 155414 408218
rect 154794 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 155414 408134
rect 154794 372454 155414 407898
rect 154794 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 155414 372454
rect 154794 372134 155414 372218
rect 154794 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 155414 372134
rect 154794 336454 155414 371898
rect 154794 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 155414 336454
rect 154794 336134 155414 336218
rect 154794 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 155414 336134
rect 154794 300454 155414 335898
rect 154794 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 155414 300454
rect 154794 300134 155414 300218
rect 154794 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 155414 300134
rect 154794 264454 155414 299898
rect 154794 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 155414 264454
rect 154794 264134 155414 264218
rect 154794 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 155414 264134
rect 154794 248684 155414 263898
rect 159294 707718 159914 711590
rect 159294 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 159914 707718
rect 159294 707398 159914 707482
rect 159294 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 159914 707398
rect 159294 700954 159914 707162
rect 159294 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 159914 700954
rect 159294 700634 159914 700718
rect 159294 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 159914 700634
rect 159294 664954 159914 700398
rect 159294 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 159914 664954
rect 159294 664634 159914 664718
rect 159294 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 159914 664634
rect 159294 628954 159914 664398
rect 159294 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 159914 628954
rect 159294 628634 159914 628718
rect 159294 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 159914 628634
rect 159294 592954 159914 628398
rect 159294 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 159914 592954
rect 159294 592634 159914 592718
rect 159294 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 159914 592634
rect 159294 556954 159914 592398
rect 159294 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 159914 556954
rect 159294 556634 159914 556718
rect 159294 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 159914 556634
rect 159294 520954 159914 556398
rect 159294 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 159914 520954
rect 159294 520634 159914 520718
rect 159294 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 159914 520634
rect 159294 484954 159914 520398
rect 159294 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 159914 484954
rect 159294 484634 159914 484718
rect 159294 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 159914 484634
rect 159294 448954 159914 484398
rect 159294 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 159914 448954
rect 159294 448634 159914 448718
rect 159294 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 159914 448634
rect 159294 412954 159914 448398
rect 159294 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 159914 412954
rect 159294 412634 159914 412718
rect 159294 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 159914 412634
rect 159294 376954 159914 412398
rect 159294 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 159914 376954
rect 159294 376634 159914 376718
rect 159294 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 159914 376634
rect 159294 340954 159914 376398
rect 159294 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 159914 340954
rect 159294 340634 159914 340718
rect 159294 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 159914 340634
rect 159294 304954 159914 340398
rect 159294 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 159914 304954
rect 159294 304634 159914 304718
rect 159294 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 159914 304634
rect 159294 268954 159914 304398
rect 159294 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 159914 268954
rect 159294 268634 159914 268718
rect 159294 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 159914 268634
rect 159294 248684 159914 268398
rect 163794 708678 164414 711590
rect 163794 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 164414 708678
rect 163794 708358 164414 708442
rect 163794 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 164414 708358
rect 163794 669454 164414 708122
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 248684 164414 272898
rect 168294 709638 168914 711590
rect 168294 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 168914 709638
rect 168294 709318 168914 709402
rect 168294 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 168914 709318
rect 168294 673954 168914 709082
rect 168294 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 168914 673954
rect 168294 673634 168914 673718
rect 168294 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 168914 673634
rect 168294 637954 168914 673398
rect 168294 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 168914 637954
rect 168294 637634 168914 637718
rect 168294 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 168914 637634
rect 168294 601954 168914 637398
rect 168294 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 168914 601954
rect 168294 601634 168914 601718
rect 168294 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 168914 601634
rect 168294 565954 168914 601398
rect 168294 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 168914 565954
rect 168294 565634 168914 565718
rect 168294 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 168914 565634
rect 168294 529954 168914 565398
rect 168294 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 168914 529954
rect 168294 529634 168914 529718
rect 168294 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 168914 529634
rect 168294 493954 168914 529398
rect 168294 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 168914 493954
rect 168294 493634 168914 493718
rect 168294 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 168914 493634
rect 168294 457954 168914 493398
rect 168294 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 168914 457954
rect 168294 457634 168914 457718
rect 168294 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 168914 457634
rect 168294 421954 168914 457398
rect 168294 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 168914 421954
rect 168294 421634 168914 421718
rect 168294 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 168914 421634
rect 168294 385954 168914 421398
rect 168294 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 168914 385954
rect 168294 385634 168914 385718
rect 168294 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 168914 385634
rect 168294 349954 168914 385398
rect 168294 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 168914 349954
rect 168294 349634 168914 349718
rect 168294 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 168914 349634
rect 168294 313954 168914 349398
rect 168294 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 168914 313954
rect 168294 313634 168914 313718
rect 168294 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 168914 313634
rect 168294 277954 168914 313398
rect 168294 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 168914 277954
rect 168294 277634 168914 277718
rect 168294 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 168914 277634
rect 168294 248684 168914 277398
rect 172794 710598 173414 711590
rect 172794 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 173414 710598
rect 172794 710278 173414 710362
rect 172794 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 173414 710278
rect 172794 678454 173414 710042
rect 172794 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 173414 678454
rect 172794 678134 173414 678218
rect 172794 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 173414 678134
rect 172794 642454 173414 677898
rect 172794 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 173414 642454
rect 172794 642134 173414 642218
rect 172794 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 173414 642134
rect 172794 606454 173414 641898
rect 172794 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 173414 606454
rect 172794 606134 173414 606218
rect 172794 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 173414 606134
rect 172794 570454 173414 605898
rect 172794 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 173414 570454
rect 172794 570134 173414 570218
rect 172794 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 173414 570134
rect 172794 534454 173414 569898
rect 172794 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 173414 534454
rect 172794 534134 173414 534218
rect 172794 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 173414 534134
rect 172794 498454 173414 533898
rect 172794 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 173414 498454
rect 172794 498134 173414 498218
rect 172794 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 173414 498134
rect 172794 462454 173414 497898
rect 172794 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 173414 462454
rect 172794 462134 173414 462218
rect 172794 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 173414 462134
rect 172794 426454 173414 461898
rect 172794 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 173414 426454
rect 172794 426134 173414 426218
rect 172794 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 173414 426134
rect 172794 390454 173414 425898
rect 172794 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 173414 390454
rect 172794 390134 173414 390218
rect 172794 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 173414 390134
rect 172794 354454 173414 389898
rect 172794 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 173414 354454
rect 172794 354134 173414 354218
rect 172794 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 173414 354134
rect 172794 318454 173414 353898
rect 172794 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 173414 318454
rect 172794 318134 173414 318218
rect 172794 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 173414 318134
rect 172794 282454 173414 317898
rect 172794 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 173414 282454
rect 172794 282134 173414 282218
rect 172794 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 173414 282134
rect 172794 248684 173414 281898
rect 177294 711558 177914 711590
rect 177294 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 177914 711558
rect 177294 711238 177914 711322
rect 177294 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 177914 711238
rect 177294 682954 177914 711002
rect 177294 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 177914 682954
rect 177294 682634 177914 682718
rect 177294 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 177914 682634
rect 177294 646954 177914 682398
rect 177294 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 177914 646954
rect 177294 646634 177914 646718
rect 177294 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 177914 646634
rect 177294 610954 177914 646398
rect 177294 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 177914 610954
rect 177294 610634 177914 610718
rect 177294 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 177914 610634
rect 177294 574954 177914 610398
rect 177294 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 177914 574954
rect 177294 574634 177914 574718
rect 177294 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 177914 574634
rect 177294 538954 177914 574398
rect 177294 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 177914 538954
rect 177294 538634 177914 538718
rect 177294 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 177914 538634
rect 177294 502954 177914 538398
rect 177294 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 177914 502954
rect 177294 502634 177914 502718
rect 177294 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 177914 502634
rect 177294 466954 177914 502398
rect 177294 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 177914 466954
rect 177294 466634 177914 466718
rect 177294 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 177914 466634
rect 177294 430954 177914 466398
rect 177294 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 177914 430954
rect 177294 430634 177914 430718
rect 177294 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 177914 430634
rect 177294 394954 177914 430398
rect 177294 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 177914 394954
rect 177294 394634 177914 394718
rect 177294 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 177914 394634
rect 177294 358954 177914 394398
rect 177294 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 177914 358954
rect 177294 358634 177914 358718
rect 177294 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 177914 358634
rect 177294 322954 177914 358398
rect 177294 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 177914 322954
rect 177294 322634 177914 322718
rect 177294 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 177914 322634
rect 177294 286954 177914 322398
rect 177294 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 177914 286954
rect 177294 286634 177914 286718
rect 177294 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 177914 286634
rect 177294 250954 177914 286398
rect 177294 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 177914 250954
rect 177294 250634 177914 250718
rect 177294 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 177914 250634
rect 177294 248684 177914 250398
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 248684 182414 254898
rect 186294 705798 186914 711590
rect 186294 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 186914 705798
rect 186294 705478 186914 705562
rect 186294 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 186914 705478
rect 186294 691954 186914 705242
rect 186294 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 186914 691954
rect 186294 691634 186914 691718
rect 186294 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 186914 691634
rect 186294 655954 186914 691398
rect 186294 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 186914 655954
rect 186294 655634 186914 655718
rect 186294 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 186914 655634
rect 186294 619954 186914 655398
rect 186294 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 186914 619954
rect 186294 619634 186914 619718
rect 186294 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 186914 619634
rect 186294 583954 186914 619398
rect 186294 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 186914 583954
rect 186294 583634 186914 583718
rect 186294 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 186914 583634
rect 186294 547954 186914 583398
rect 186294 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 186914 547954
rect 186294 547634 186914 547718
rect 186294 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 186914 547634
rect 186294 511954 186914 547398
rect 186294 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 186914 511954
rect 186294 511634 186914 511718
rect 186294 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 186914 511634
rect 186294 475954 186914 511398
rect 186294 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 186914 475954
rect 186294 475634 186914 475718
rect 186294 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 186914 475634
rect 186294 439954 186914 475398
rect 186294 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 186914 439954
rect 186294 439634 186914 439718
rect 186294 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 186914 439634
rect 186294 403954 186914 439398
rect 186294 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 186914 403954
rect 186294 403634 186914 403718
rect 186294 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 186914 403634
rect 186294 367954 186914 403398
rect 186294 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 186914 367954
rect 186294 367634 186914 367718
rect 186294 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 186914 367634
rect 186294 331954 186914 367398
rect 186294 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 186914 331954
rect 186294 331634 186914 331718
rect 186294 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 186914 331634
rect 186294 295954 186914 331398
rect 186294 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 186914 295954
rect 186294 295634 186914 295718
rect 186294 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 186914 295634
rect 186294 259954 186914 295398
rect 186294 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 186914 259954
rect 186294 259634 186914 259718
rect 186294 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 186914 259634
rect 186294 248684 186914 259398
rect 190794 706758 191414 711590
rect 190794 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 191414 706758
rect 190794 706438 191414 706522
rect 190794 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 191414 706438
rect 190794 696454 191414 706202
rect 190794 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 191414 696454
rect 190794 696134 191414 696218
rect 190794 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 191414 696134
rect 190794 660454 191414 695898
rect 190794 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 191414 660454
rect 190794 660134 191414 660218
rect 190794 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 191414 660134
rect 190794 624454 191414 659898
rect 190794 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 191414 624454
rect 190794 624134 191414 624218
rect 190794 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 191414 624134
rect 190794 588454 191414 623898
rect 190794 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 191414 588454
rect 190794 588134 191414 588218
rect 190794 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 191414 588134
rect 190794 552454 191414 587898
rect 190794 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 191414 552454
rect 190794 552134 191414 552218
rect 190794 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 191414 552134
rect 190794 516454 191414 551898
rect 190794 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 191414 516454
rect 190794 516134 191414 516218
rect 190794 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 191414 516134
rect 190794 480454 191414 515898
rect 190794 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 191414 480454
rect 190794 480134 191414 480218
rect 190794 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 191414 480134
rect 190794 444454 191414 479898
rect 190794 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 191414 444454
rect 190794 444134 191414 444218
rect 190794 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 191414 444134
rect 190794 408454 191414 443898
rect 190794 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 191414 408454
rect 190794 408134 191414 408218
rect 190794 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 191414 408134
rect 190794 372454 191414 407898
rect 190794 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 191414 372454
rect 190794 372134 191414 372218
rect 190794 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 191414 372134
rect 190794 336454 191414 371898
rect 190794 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 191414 336454
rect 190794 336134 191414 336218
rect 190794 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 191414 336134
rect 190794 300454 191414 335898
rect 190794 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 191414 300454
rect 190794 300134 191414 300218
rect 190794 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 191414 300134
rect 190794 264454 191414 299898
rect 190794 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 191414 264454
rect 190794 264134 191414 264218
rect 190794 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 191414 264134
rect 190794 248684 191414 263898
rect 195294 707718 195914 711590
rect 195294 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 195914 707718
rect 195294 707398 195914 707482
rect 195294 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 195914 707398
rect 195294 700954 195914 707162
rect 195294 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 195914 700954
rect 195294 700634 195914 700718
rect 195294 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 195914 700634
rect 195294 664954 195914 700398
rect 195294 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 195914 664954
rect 195294 664634 195914 664718
rect 195294 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 195914 664634
rect 195294 628954 195914 664398
rect 195294 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 195914 628954
rect 195294 628634 195914 628718
rect 195294 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 195914 628634
rect 195294 592954 195914 628398
rect 195294 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 195914 592954
rect 195294 592634 195914 592718
rect 195294 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 195914 592634
rect 195294 556954 195914 592398
rect 195294 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 195914 556954
rect 195294 556634 195914 556718
rect 195294 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 195914 556634
rect 195294 520954 195914 556398
rect 195294 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 195914 520954
rect 195294 520634 195914 520718
rect 195294 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 195914 520634
rect 195294 484954 195914 520398
rect 195294 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 195914 484954
rect 195294 484634 195914 484718
rect 195294 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 195914 484634
rect 195294 448954 195914 484398
rect 195294 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 195914 448954
rect 195294 448634 195914 448718
rect 195294 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 195914 448634
rect 195294 412954 195914 448398
rect 195294 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 195914 412954
rect 195294 412634 195914 412718
rect 195294 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 195914 412634
rect 195294 376954 195914 412398
rect 195294 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 195914 376954
rect 195294 376634 195914 376718
rect 195294 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 195914 376634
rect 195294 340954 195914 376398
rect 195294 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 195914 340954
rect 195294 340634 195914 340718
rect 195294 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 195914 340634
rect 195294 304954 195914 340398
rect 195294 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 195914 304954
rect 195294 304634 195914 304718
rect 195294 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 195914 304634
rect 195294 268954 195914 304398
rect 195294 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 195914 268954
rect 195294 268634 195914 268718
rect 195294 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 195914 268634
rect 195294 248684 195914 268398
rect 199794 708678 200414 711590
rect 199794 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 200414 708678
rect 199794 708358 200414 708442
rect 199794 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 200414 708358
rect 199794 669454 200414 708122
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199794 248684 200414 272898
rect 204294 709638 204914 711590
rect 204294 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 204914 709638
rect 204294 709318 204914 709402
rect 204294 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 204914 709318
rect 204294 673954 204914 709082
rect 204294 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 204914 673954
rect 204294 673634 204914 673718
rect 204294 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 204914 673634
rect 204294 637954 204914 673398
rect 204294 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 204914 637954
rect 204294 637634 204914 637718
rect 204294 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 204914 637634
rect 204294 601954 204914 637398
rect 204294 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 204914 601954
rect 204294 601634 204914 601718
rect 204294 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 204914 601634
rect 204294 565954 204914 601398
rect 204294 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 204914 565954
rect 204294 565634 204914 565718
rect 204294 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 204914 565634
rect 204294 529954 204914 565398
rect 204294 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 204914 529954
rect 204294 529634 204914 529718
rect 204294 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 204914 529634
rect 204294 493954 204914 529398
rect 204294 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 204914 493954
rect 204294 493634 204914 493718
rect 204294 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 204914 493634
rect 204294 457954 204914 493398
rect 204294 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 204914 457954
rect 204294 457634 204914 457718
rect 204294 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 204914 457634
rect 204294 421954 204914 457398
rect 204294 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 204914 421954
rect 204294 421634 204914 421718
rect 204294 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 204914 421634
rect 204294 385954 204914 421398
rect 204294 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 204914 385954
rect 204294 385634 204914 385718
rect 204294 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 204914 385634
rect 204294 349954 204914 385398
rect 204294 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 204914 349954
rect 204294 349634 204914 349718
rect 204294 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 204914 349634
rect 204294 313954 204914 349398
rect 204294 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 204914 313954
rect 204294 313634 204914 313718
rect 204294 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 204914 313634
rect 204294 277954 204914 313398
rect 204294 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 204914 277954
rect 204294 277634 204914 277718
rect 204294 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 204914 277634
rect 204294 248684 204914 277398
rect 208794 710598 209414 711590
rect 208794 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 209414 710598
rect 208794 710278 209414 710362
rect 208794 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 209414 710278
rect 208794 678454 209414 710042
rect 208794 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 209414 678454
rect 208794 678134 209414 678218
rect 208794 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 209414 678134
rect 208794 642454 209414 677898
rect 208794 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 209414 642454
rect 208794 642134 209414 642218
rect 208794 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 209414 642134
rect 208794 606454 209414 641898
rect 208794 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 209414 606454
rect 208794 606134 209414 606218
rect 208794 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 209414 606134
rect 208794 570454 209414 605898
rect 208794 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 209414 570454
rect 208794 570134 209414 570218
rect 208794 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 209414 570134
rect 208794 534454 209414 569898
rect 208794 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 209414 534454
rect 208794 534134 209414 534218
rect 208794 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 209414 534134
rect 208794 498454 209414 533898
rect 208794 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 209414 498454
rect 208794 498134 209414 498218
rect 208794 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 209414 498134
rect 208794 462454 209414 497898
rect 208794 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 209414 462454
rect 208794 462134 209414 462218
rect 208794 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 209414 462134
rect 208794 426454 209414 461898
rect 208794 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 209414 426454
rect 208794 426134 209414 426218
rect 208794 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 209414 426134
rect 208794 390454 209414 425898
rect 208794 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 209414 390454
rect 208794 390134 209414 390218
rect 208794 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 209414 390134
rect 208794 354454 209414 389898
rect 208794 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 209414 354454
rect 208794 354134 209414 354218
rect 208794 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 209414 354134
rect 208794 318454 209414 353898
rect 208794 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 209414 318454
rect 208794 318134 209414 318218
rect 208794 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 209414 318134
rect 208794 282454 209414 317898
rect 208794 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 209414 282454
rect 208794 282134 209414 282218
rect 208794 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 209414 282134
rect 208794 248684 209414 281898
rect 213294 711558 213914 711590
rect 213294 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 213914 711558
rect 213294 711238 213914 711322
rect 213294 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 213914 711238
rect 213294 682954 213914 711002
rect 213294 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 213914 682954
rect 213294 682634 213914 682718
rect 213294 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 213914 682634
rect 213294 646954 213914 682398
rect 213294 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 213914 646954
rect 213294 646634 213914 646718
rect 213294 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 213914 646634
rect 213294 610954 213914 646398
rect 213294 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 213914 610954
rect 213294 610634 213914 610718
rect 213294 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 213914 610634
rect 213294 574954 213914 610398
rect 213294 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 213914 574954
rect 213294 574634 213914 574718
rect 213294 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 213914 574634
rect 213294 538954 213914 574398
rect 213294 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 213914 538954
rect 213294 538634 213914 538718
rect 213294 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 213914 538634
rect 213294 502954 213914 538398
rect 213294 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 213914 502954
rect 213294 502634 213914 502718
rect 213294 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 213914 502634
rect 213294 466954 213914 502398
rect 213294 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 213914 466954
rect 213294 466634 213914 466718
rect 213294 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 213914 466634
rect 213294 430954 213914 466398
rect 213294 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 213914 430954
rect 213294 430634 213914 430718
rect 213294 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 213914 430634
rect 213294 394954 213914 430398
rect 213294 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 213914 394954
rect 213294 394634 213914 394718
rect 213294 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 213914 394634
rect 213294 358954 213914 394398
rect 213294 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 213914 358954
rect 213294 358634 213914 358718
rect 213294 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 213914 358634
rect 213294 322954 213914 358398
rect 213294 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 213914 322954
rect 213294 322634 213914 322718
rect 213294 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 213914 322634
rect 213294 286954 213914 322398
rect 213294 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 213914 286954
rect 213294 286634 213914 286718
rect 213294 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 213914 286634
rect 213294 250954 213914 286398
rect 213294 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 213914 250954
rect 213294 250634 213914 250718
rect 213294 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 213914 250634
rect 213294 248684 213914 250398
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 248684 218414 254898
rect 222294 705798 222914 711590
rect 222294 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 222914 705798
rect 222294 705478 222914 705562
rect 222294 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 222914 705478
rect 222294 691954 222914 705242
rect 222294 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 222914 691954
rect 222294 691634 222914 691718
rect 222294 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 222914 691634
rect 222294 655954 222914 691398
rect 222294 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 222914 655954
rect 222294 655634 222914 655718
rect 222294 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 222914 655634
rect 222294 619954 222914 655398
rect 222294 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 222914 619954
rect 222294 619634 222914 619718
rect 222294 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 222914 619634
rect 222294 583954 222914 619398
rect 222294 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 222914 583954
rect 222294 583634 222914 583718
rect 222294 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 222914 583634
rect 222294 547954 222914 583398
rect 222294 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 222914 547954
rect 222294 547634 222914 547718
rect 222294 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 222914 547634
rect 222294 511954 222914 547398
rect 222294 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 222914 511954
rect 222294 511634 222914 511718
rect 222294 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 222914 511634
rect 222294 475954 222914 511398
rect 222294 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 222914 475954
rect 222294 475634 222914 475718
rect 222294 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 222914 475634
rect 222294 439954 222914 475398
rect 222294 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 222914 439954
rect 222294 439634 222914 439718
rect 222294 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 222914 439634
rect 222294 403954 222914 439398
rect 222294 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 222914 403954
rect 222294 403634 222914 403718
rect 222294 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 222914 403634
rect 222294 367954 222914 403398
rect 222294 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 222914 367954
rect 222294 367634 222914 367718
rect 222294 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 222914 367634
rect 222294 331954 222914 367398
rect 222294 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 222914 331954
rect 222294 331634 222914 331718
rect 222294 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 222914 331634
rect 222294 295954 222914 331398
rect 222294 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 222914 295954
rect 222294 295634 222914 295718
rect 222294 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 222914 295634
rect 222294 259954 222914 295398
rect 222294 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 222914 259954
rect 222294 259634 222914 259718
rect 222294 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 222914 259634
rect 222294 248684 222914 259398
rect 226794 706758 227414 711590
rect 226794 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 227414 706758
rect 226794 706438 227414 706522
rect 226794 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 227414 706438
rect 226794 696454 227414 706202
rect 226794 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 227414 696454
rect 226794 696134 227414 696218
rect 226794 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 227414 696134
rect 226794 660454 227414 695898
rect 226794 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 227414 660454
rect 226794 660134 227414 660218
rect 226794 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 227414 660134
rect 226794 624454 227414 659898
rect 226794 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 227414 624454
rect 226794 624134 227414 624218
rect 226794 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 227414 624134
rect 226794 588454 227414 623898
rect 226794 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 227414 588454
rect 226794 588134 227414 588218
rect 226794 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 227414 588134
rect 226794 552454 227414 587898
rect 226794 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 227414 552454
rect 226794 552134 227414 552218
rect 226794 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 227414 552134
rect 226794 516454 227414 551898
rect 226794 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 227414 516454
rect 226794 516134 227414 516218
rect 226794 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 227414 516134
rect 226794 480454 227414 515898
rect 226794 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 227414 480454
rect 226794 480134 227414 480218
rect 226794 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 227414 480134
rect 226794 444454 227414 479898
rect 226794 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 227414 444454
rect 226794 444134 227414 444218
rect 226794 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 227414 444134
rect 226794 408454 227414 443898
rect 226794 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 227414 408454
rect 226794 408134 227414 408218
rect 226794 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 227414 408134
rect 226794 372454 227414 407898
rect 226794 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 227414 372454
rect 226794 372134 227414 372218
rect 226794 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 227414 372134
rect 226794 336454 227414 371898
rect 226794 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 227414 336454
rect 226794 336134 227414 336218
rect 226794 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 227414 336134
rect 226794 300454 227414 335898
rect 226794 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 227414 300454
rect 226794 300134 227414 300218
rect 226794 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 227414 300134
rect 226794 264454 227414 299898
rect 226794 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 227414 264454
rect 226794 264134 227414 264218
rect 226794 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 227414 264134
rect 226794 248684 227414 263898
rect 231294 707718 231914 711590
rect 231294 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 231914 707718
rect 231294 707398 231914 707482
rect 231294 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 231914 707398
rect 231294 700954 231914 707162
rect 231294 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 231914 700954
rect 231294 700634 231914 700718
rect 231294 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 231914 700634
rect 231294 664954 231914 700398
rect 231294 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 231914 664954
rect 231294 664634 231914 664718
rect 231294 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 231914 664634
rect 231294 628954 231914 664398
rect 231294 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 231914 628954
rect 231294 628634 231914 628718
rect 231294 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 231914 628634
rect 231294 592954 231914 628398
rect 231294 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 231914 592954
rect 231294 592634 231914 592718
rect 231294 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 231914 592634
rect 231294 556954 231914 592398
rect 231294 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 231914 556954
rect 231294 556634 231914 556718
rect 231294 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 231914 556634
rect 231294 520954 231914 556398
rect 231294 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 231914 520954
rect 231294 520634 231914 520718
rect 231294 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 231914 520634
rect 231294 484954 231914 520398
rect 231294 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 231914 484954
rect 231294 484634 231914 484718
rect 231294 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 231914 484634
rect 231294 448954 231914 484398
rect 231294 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 231914 448954
rect 231294 448634 231914 448718
rect 231294 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 231914 448634
rect 231294 412954 231914 448398
rect 231294 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 231914 412954
rect 231294 412634 231914 412718
rect 231294 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 231914 412634
rect 231294 376954 231914 412398
rect 231294 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 231914 376954
rect 231294 376634 231914 376718
rect 231294 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 231914 376634
rect 231294 340954 231914 376398
rect 231294 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 231914 340954
rect 231294 340634 231914 340718
rect 231294 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 231914 340634
rect 231294 304954 231914 340398
rect 231294 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 231914 304954
rect 231294 304634 231914 304718
rect 231294 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 231914 304634
rect 231294 268954 231914 304398
rect 231294 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 231914 268954
rect 231294 268634 231914 268718
rect 231294 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 231914 268634
rect 231294 248684 231914 268398
rect 235794 708678 236414 711590
rect 235794 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 236414 708678
rect 235794 708358 236414 708442
rect 235794 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 236414 708358
rect 235794 669454 236414 708122
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381454 236414 416898
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 273454 236414 308898
rect 235794 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 236414 273454
rect 235794 273134 236414 273218
rect 235794 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 236414 273134
rect 235794 248684 236414 272898
rect 240294 709638 240914 711590
rect 240294 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 240914 709638
rect 240294 709318 240914 709402
rect 240294 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 240914 709318
rect 240294 673954 240914 709082
rect 240294 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 240914 673954
rect 240294 673634 240914 673718
rect 240294 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 240914 673634
rect 240294 637954 240914 673398
rect 240294 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 240914 637954
rect 240294 637634 240914 637718
rect 240294 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 240914 637634
rect 240294 601954 240914 637398
rect 240294 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 240914 601954
rect 240294 601634 240914 601718
rect 240294 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 240914 601634
rect 240294 565954 240914 601398
rect 240294 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 240914 565954
rect 240294 565634 240914 565718
rect 240294 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 240914 565634
rect 240294 529954 240914 565398
rect 240294 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 240914 529954
rect 240294 529634 240914 529718
rect 240294 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 240914 529634
rect 240294 493954 240914 529398
rect 240294 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 240914 493954
rect 240294 493634 240914 493718
rect 240294 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 240914 493634
rect 240294 457954 240914 493398
rect 240294 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 240914 457954
rect 240294 457634 240914 457718
rect 240294 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 240914 457634
rect 240294 421954 240914 457398
rect 240294 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 240914 421954
rect 240294 421634 240914 421718
rect 240294 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 240914 421634
rect 240294 385954 240914 421398
rect 240294 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 240914 385954
rect 240294 385634 240914 385718
rect 240294 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 240914 385634
rect 240294 349954 240914 385398
rect 240294 349718 240326 349954
rect 240562 349718 240646 349954
rect 240882 349718 240914 349954
rect 240294 349634 240914 349718
rect 240294 349398 240326 349634
rect 240562 349398 240646 349634
rect 240882 349398 240914 349634
rect 240294 313954 240914 349398
rect 240294 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 240914 313954
rect 240294 313634 240914 313718
rect 240294 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 240914 313634
rect 240294 277954 240914 313398
rect 240294 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 240914 277954
rect 240294 277634 240914 277718
rect 240294 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 240914 277634
rect 240294 248684 240914 277398
rect 244794 710598 245414 711590
rect 244794 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 245414 710598
rect 244794 710278 245414 710362
rect 244794 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 245414 710278
rect 244794 678454 245414 710042
rect 244794 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 245414 678454
rect 244794 678134 245414 678218
rect 244794 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 245414 678134
rect 244794 642454 245414 677898
rect 244794 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 245414 642454
rect 244794 642134 245414 642218
rect 244794 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 245414 642134
rect 244794 606454 245414 641898
rect 244794 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 245414 606454
rect 244794 606134 245414 606218
rect 244794 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 245414 606134
rect 244794 570454 245414 605898
rect 244794 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 245414 570454
rect 244794 570134 245414 570218
rect 244794 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 245414 570134
rect 244794 534454 245414 569898
rect 244794 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 245414 534454
rect 244794 534134 245414 534218
rect 244794 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 245414 534134
rect 244794 498454 245414 533898
rect 244794 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 245414 498454
rect 244794 498134 245414 498218
rect 244794 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 245414 498134
rect 244794 462454 245414 497898
rect 244794 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 245414 462454
rect 244794 462134 245414 462218
rect 244794 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 245414 462134
rect 244794 426454 245414 461898
rect 244794 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 245414 426454
rect 244794 426134 245414 426218
rect 244794 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 245414 426134
rect 244794 390454 245414 425898
rect 244794 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 245414 390454
rect 244794 390134 245414 390218
rect 244794 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 245414 390134
rect 244794 354454 245414 389898
rect 244794 354218 244826 354454
rect 245062 354218 245146 354454
rect 245382 354218 245414 354454
rect 244794 354134 245414 354218
rect 244794 353898 244826 354134
rect 245062 353898 245146 354134
rect 245382 353898 245414 354134
rect 244794 318454 245414 353898
rect 244794 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 245414 318454
rect 244794 318134 245414 318218
rect 244794 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 245414 318134
rect 244794 282454 245414 317898
rect 244794 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 245414 282454
rect 244794 282134 245414 282218
rect 244794 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 245414 282134
rect 244794 248684 245414 281898
rect 249294 711558 249914 711590
rect 249294 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 249914 711558
rect 249294 711238 249914 711322
rect 249294 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 249914 711238
rect 249294 682954 249914 711002
rect 249294 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 249914 682954
rect 249294 682634 249914 682718
rect 249294 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 249914 682634
rect 249294 646954 249914 682398
rect 249294 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 249914 646954
rect 249294 646634 249914 646718
rect 249294 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 249914 646634
rect 249294 610954 249914 646398
rect 249294 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 249914 610954
rect 249294 610634 249914 610718
rect 249294 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 249914 610634
rect 249294 574954 249914 610398
rect 249294 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 249914 574954
rect 249294 574634 249914 574718
rect 249294 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 249914 574634
rect 249294 538954 249914 574398
rect 249294 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 249914 538954
rect 249294 538634 249914 538718
rect 249294 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 249914 538634
rect 249294 502954 249914 538398
rect 249294 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 249914 502954
rect 249294 502634 249914 502718
rect 249294 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 249914 502634
rect 249294 466954 249914 502398
rect 249294 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 249914 466954
rect 249294 466634 249914 466718
rect 249294 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 249914 466634
rect 249294 430954 249914 466398
rect 249294 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 249914 430954
rect 249294 430634 249914 430718
rect 249294 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 249914 430634
rect 249294 394954 249914 430398
rect 249294 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 249914 394954
rect 249294 394634 249914 394718
rect 249294 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 249914 394634
rect 249294 358954 249914 394398
rect 249294 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 249914 358954
rect 249294 358634 249914 358718
rect 249294 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 249914 358634
rect 249294 322954 249914 358398
rect 249294 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 249914 322954
rect 249294 322634 249914 322718
rect 249294 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 249914 322634
rect 249294 286954 249914 322398
rect 249294 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 249914 286954
rect 249294 286634 249914 286718
rect 249294 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 249914 286634
rect 249294 250954 249914 286398
rect 249294 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 249914 250954
rect 249294 250634 249914 250718
rect 249294 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 249914 250634
rect 249294 248684 249914 250398
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 291454 254414 326898
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 248684 254414 254898
rect 258294 705798 258914 711590
rect 258294 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 258914 705798
rect 258294 705478 258914 705562
rect 258294 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 258914 705478
rect 258294 691954 258914 705242
rect 258294 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 258914 691954
rect 258294 691634 258914 691718
rect 258294 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 258914 691634
rect 258294 655954 258914 691398
rect 258294 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 258914 655954
rect 258294 655634 258914 655718
rect 258294 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 258914 655634
rect 258294 619954 258914 655398
rect 258294 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 258914 619954
rect 258294 619634 258914 619718
rect 258294 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 258914 619634
rect 258294 583954 258914 619398
rect 258294 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 258914 583954
rect 258294 583634 258914 583718
rect 258294 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 258914 583634
rect 258294 547954 258914 583398
rect 258294 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 258914 547954
rect 258294 547634 258914 547718
rect 258294 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 258914 547634
rect 258294 511954 258914 547398
rect 258294 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 258914 511954
rect 258294 511634 258914 511718
rect 258294 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 258914 511634
rect 258294 475954 258914 511398
rect 258294 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 258914 475954
rect 258294 475634 258914 475718
rect 258294 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 258914 475634
rect 258294 439954 258914 475398
rect 258294 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 258914 439954
rect 258294 439634 258914 439718
rect 258294 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 258914 439634
rect 258294 403954 258914 439398
rect 258294 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 258914 403954
rect 258294 403634 258914 403718
rect 258294 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 258914 403634
rect 258294 367954 258914 403398
rect 258294 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 258914 367954
rect 258294 367634 258914 367718
rect 258294 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 258914 367634
rect 258294 331954 258914 367398
rect 258294 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 258914 331954
rect 258294 331634 258914 331718
rect 258294 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 258914 331634
rect 258294 295954 258914 331398
rect 258294 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 258914 295954
rect 258294 295634 258914 295718
rect 258294 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 258914 295634
rect 258294 259954 258914 295398
rect 258294 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 258914 259954
rect 258294 259634 258914 259718
rect 258294 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 258914 259634
rect 258294 248684 258914 259398
rect 262794 706758 263414 711590
rect 262794 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 263414 706758
rect 262794 706438 263414 706522
rect 262794 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 263414 706438
rect 262794 696454 263414 706202
rect 262794 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 263414 696454
rect 262794 696134 263414 696218
rect 262794 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 263414 696134
rect 262794 660454 263414 695898
rect 262794 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 263414 660454
rect 262794 660134 263414 660218
rect 262794 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 263414 660134
rect 262794 624454 263414 659898
rect 262794 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 263414 624454
rect 262794 624134 263414 624218
rect 262794 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 263414 624134
rect 262794 588454 263414 623898
rect 262794 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 263414 588454
rect 262794 588134 263414 588218
rect 262794 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 263414 588134
rect 262794 552454 263414 587898
rect 262794 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 263414 552454
rect 262794 552134 263414 552218
rect 262794 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 263414 552134
rect 262794 516454 263414 551898
rect 262794 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 263414 516454
rect 262794 516134 263414 516218
rect 262794 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 263414 516134
rect 262794 480454 263414 515898
rect 262794 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 263414 480454
rect 262794 480134 263414 480218
rect 262794 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 263414 480134
rect 262794 444454 263414 479898
rect 262794 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 263414 444454
rect 262794 444134 263414 444218
rect 262794 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 263414 444134
rect 262794 408454 263414 443898
rect 262794 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 263414 408454
rect 262794 408134 263414 408218
rect 262794 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 263414 408134
rect 262794 372454 263414 407898
rect 262794 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 263414 372454
rect 262794 372134 263414 372218
rect 262794 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 263414 372134
rect 262794 336454 263414 371898
rect 262794 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 263414 336454
rect 262794 336134 263414 336218
rect 262794 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 263414 336134
rect 262794 300454 263414 335898
rect 262794 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 263414 300454
rect 262794 300134 263414 300218
rect 262794 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 263414 300134
rect 262794 264454 263414 299898
rect 262794 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 263414 264454
rect 262794 264134 263414 264218
rect 262794 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 263414 264134
rect 262794 248684 263414 263898
rect 267294 707718 267914 711590
rect 267294 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 267914 707718
rect 267294 707398 267914 707482
rect 267294 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 267914 707398
rect 267294 700954 267914 707162
rect 267294 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 267914 700954
rect 267294 700634 267914 700718
rect 267294 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 267914 700634
rect 267294 664954 267914 700398
rect 267294 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 267914 664954
rect 267294 664634 267914 664718
rect 267294 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 267914 664634
rect 267294 628954 267914 664398
rect 267294 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 267914 628954
rect 267294 628634 267914 628718
rect 267294 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 267914 628634
rect 267294 592954 267914 628398
rect 267294 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 267914 592954
rect 267294 592634 267914 592718
rect 267294 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 267914 592634
rect 267294 556954 267914 592398
rect 267294 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 267914 556954
rect 267294 556634 267914 556718
rect 267294 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 267914 556634
rect 267294 520954 267914 556398
rect 267294 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 267914 520954
rect 267294 520634 267914 520718
rect 267294 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 267914 520634
rect 267294 484954 267914 520398
rect 267294 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 267914 484954
rect 267294 484634 267914 484718
rect 267294 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 267914 484634
rect 267294 448954 267914 484398
rect 267294 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 267914 448954
rect 267294 448634 267914 448718
rect 267294 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 267914 448634
rect 267294 412954 267914 448398
rect 267294 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 267914 412954
rect 267294 412634 267914 412718
rect 267294 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 267914 412634
rect 267294 376954 267914 412398
rect 267294 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 267914 376954
rect 267294 376634 267914 376718
rect 267294 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 267914 376634
rect 267294 340954 267914 376398
rect 267294 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 267914 340954
rect 267294 340634 267914 340718
rect 267294 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 267914 340634
rect 267294 304954 267914 340398
rect 267294 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 267914 304954
rect 267294 304634 267914 304718
rect 267294 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 267914 304634
rect 267294 268954 267914 304398
rect 267294 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 267914 268954
rect 267294 268634 267914 268718
rect 267294 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 267914 268634
rect 267294 248684 267914 268398
rect 271794 708678 272414 711590
rect 271794 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 272414 708678
rect 271794 708358 272414 708442
rect 271794 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 272414 708358
rect 271794 669454 272414 708122
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 345454 272414 380898
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 273454 272414 308898
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 248684 272414 272898
rect 276294 709638 276914 711590
rect 276294 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 276914 709638
rect 276294 709318 276914 709402
rect 276294 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 276914 709318
rect 276294 673954 276914 709082
rect 276294 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 276914 673954
rect 276294 673634 276914 673718
rect 276294 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 276914 673634
rect 276294 637954 276914 673398
rect 276294 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 276914 637954
rect 276294 637634 276914 637718
rect 276294 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 276914 637634
rect 276294 601954 276914 637398
rect 276294 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 276914 601954
rect 276294 601634 276914 601718
rect 276294 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 276914 601634
rect 276294 565954 276914 601398
rect 276294 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 276914 565954
rect 276294 565634 276914 565718
rect 276294 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 276914 565634
rect 276294 529954 276914 565398
rect 276294 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 276914 529954
rect 276294 529634 276914 529718
rect 276294 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 276914 529634
rect 276294 493954 276914 529398
rect 276294 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 276914 493954
rect 276294 493634 276914 493718
rect 276294 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 276914 493634
rect 276294 457954 276914 493398
rect 276294 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 276914 457954
rect 276294 457634 276914 457718
rect 276294 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 276914 457634
rect 276294 421954 276914 457398
rect 276294 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 276914 421954
rect 276294 421634 276914 421718
rect 276294 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 276914 421634
rect 276294 385954 276914 421398
rect 276294 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 276914 385954
rect 276294 385634 276914 385718
rect 276294 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 276914 385634
rect 276294 349954 276914 385398
rect 276294 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 276914 349954
rect 276294 349634 276914 349718
rect 276294 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 276914 349634
rect 276294 313954 276914 349398
rect 276294 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 276914 313954
rect 276294 313634 276914 313718
rect 276294 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 276914 313634
rect 276294 277954 276914 313398
rect 276294 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 276914 277954
rect 276294 277634 276914 277718
rect 276294 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 276914 277634
rect 276294 248684 276914 277398
rect 280794 710598 281414 711590
rect 280794 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 281414 710598
rect 280794 710278 281414 710362
rect 280794 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 281414 710278
rect 280794 678454 281414 710042
rect 280794 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 281414 678454
rect 280794 678134 281414 678218
rect 280794 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 281414 678134
rect 280794 642454 281414 677898
rect 280794 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 281414 642454
rect 280794 642134 281414 642218
rect 280794 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 281414 642134
rect 280794 606454 281414 641898
rect 280794 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 281414 606454
rect 280794 606134 281414 606218
rect 280794 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 281414 606134
rect 280794 570454 281414 605898
rect 280794 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 281414 570454
rect 280794 570134 281414 570218
rect 280794 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 281414 570134
rect 280794 534454 281414 569898
rect 280794 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 281414 534454
rect 280794 534134 281414 534218
rect 280794 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 281414 534134
rect 280794 498454 281414 533898
rect 280794 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 281414 498454
rect 280794 498134 281414 498218
rect 280794 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 281414 498134
rect 280794 462454 281414 497898
rect 280794 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 281414 462454
rect 280794 462134 281414 462218
rect 280794 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 281414 462134
rect 280794 426454 281414 461898
rect 280794 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 281414 426454
rect 280794 426134 281414 426218
rect 280794 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 281414 426134
rect 280794 390454 281414 425898
rect 280794 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 281414 390454
rect 280794 390134 281414 390218
rect 280794 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 281414 390134
rect 280794 354454 281414 389898
rect 280794 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 281414 354454
rect 280794 354134 281414 354218
rect 280794 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 281414 354134
rect 280794 318454 281414 353898
rect 280794 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 281414 318454
rect 280794 318134 281414 318218
rect 280794 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 281414 318134
rect 280794 282454 281414 317898
rect 280794 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 281414 282454
rect 280794 282134 281414 282218
rect 280794 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 281414 282134
rect 280794 248684 281414 281898
rect 285294 711558 285914 711590
rect 285294 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 285914 711558
rect 285294 711238 285914 711322
rect 285294 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 285914 711238
rect 285294 682954 285914 711002
rect 285294 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 285914 682954
rect 285294 682634 285914 682718
rect 285294 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 285914 682634
rect 285294 646954 285914 682398
rect 285294 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 285914 646954
rect 285294 646634 285914 646718
rect 285294 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 285914 646634
rect 285294 610954 285914 646398
rect 285294 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 285914 610954
rect 285294 610634 285914 610718
rect 285294 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 285914 610634
rect 285294 574954 285914 610398
rect 285294 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 285914 574954
rect 285294 574634 285914 574718
rect 285294 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 285914 574634
rect 285294 538954 285914 574398
rect 285294 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 285914 538954
rect 285294 538634 285914 538718
rect 285294 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 285914 538634
rect 285294 502954 285914 538398
rect 285294 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 285914 502954
rect 285294 502634 285914 502718
rect 285294 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 285914 502634
rect 285294 466954 285914 502398
rect 285294 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 285914 466954
rect 285294 466634 285914 466718
rect 285294 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 285914 466634
rect 285294 430954 285914 466398
rect 285294 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 285914 430954
rect 285294 430634 285914 430718
rect 285294 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 285914 430634
rect 285294 394954 285914 430398
rect 285294 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 285914 394954
rect 285294 394634 285914 394718
rect 285294 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 285914 394634
rect 285294 358954 285914 394398
rect 285294 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 285914 358954
rect 285294 358634 285914 358718
rect 285294 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 285914 358634
rect 285294 322954 285914 358398
rect 285294 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 285914 322954
rect 285294 322634 285914 322718
rect 285294 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 285914 322634
rect 285294 286954 285914 322398
rect 285294 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 285914 286954
rect 285294 286634 285914 286718
rect 285294 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 285914 286634
rect 285294 250954 285914 286398
rect 285294 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 285914 250954
rect 285294 250634 285914 250718
rect 285294 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 285914 250634
rect 285294 248684 285914 250398
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 248684 290414 254898
rect 294294 705798 294914 711590
rect 294294 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 294914 705798
rect 294294 705478 294914 705562
rect 294294 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 294914 705478
rect 294294 691954 294914 705242
rect 294294 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 294914 691954
rect 294294 691634 294914 691718
rect 294294 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 294914 691634
rect 294294 655954 294914 691398
rect 294294 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 294914 655954
rect 294294 655634 294914 655718
rect 294294 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 294914 655634
rect 294294 619954 294914 655398
rect 294294 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 294914 619954
rect 294294 619634 294914 619718
rect 294294 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 294914 619634
rect 294294 583954 294914 619398
rect 294294 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 294914 583954
rect 294294 583634 294914 583718
rect 294294 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 294914 583634
rect 294294 547954 294914 583398
rect 294294 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 294914 547954
rect 294294 547634 294914 547718
rect 294294 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 294914 547634
rect 294294 511954 294914 547398
rect 294294 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 294914 511954
rect 294294 511634 294914 511718
rect 294294 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 294914 511634
rect 294294 475954 294914 511398
rect 294294 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 294914 475954
rect 294294 475634 294914 475718
rect 294294 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 294914 475634
rect 294294 439954 294914 475398
rect 294294 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 294914 439954
rect 294294 439634 294914 439718
rect 294294 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 294914 439634
rect 294294 403954 294914 439398
rect 294294 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 294914 403954
rect 294294 403634 294914 403718
rect 294294 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 294914 403634
rect 294294 367954 294914 403398
rect 294294 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 294914 367954
rect 294294 367634 294914 367718
rect 294294 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 294914 367634
rect 294294 331954 294914 367398
rect 294294 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 294914 331954
rect 294294 331634 294914 331718
rect 294294 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 294914 331634
rect 294294 295954 294914 331398
rect 294294 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 294914 295954
rect 294294 295634 294914 295718
rect 294294 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 294914 295634
rect 294294 259954 294914 295398
rect 294294 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 294914 259954
rect 294294 259634 294914 259718
rect 294294 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 294914 259634
rect 294294 248684 294914 259398
rect 298794 706758 299414 711590
rect 298794 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 299414 706758
rect 298794 706438 299414 706522
rect 298794 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 299414 706438
rect 298794 696454 299414 706202
rect 298794 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 299414 696454
rect 298794 696134 299414 696218
rect 298794 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 299414 696134
rect 298794 660454 299414 695898
rect 298794 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 299414 660454
rect 298794 660134 299414 660218
rect 298794 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 299414 660134
rect 298794 624454 299414 659898
rect 298794 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 299414 624454
rect 298794 624134 299414 624218
rect 298794 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 299414 624134
rect 298794 588454 299414 623898
rect 298794 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 299414 588454
rect 298794 588134 299414 588218
rect 298794 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 299414 588134
rect 298794 552454 299414 587898
rect 298794 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 299414 552454
rect 298794 552134 299414 552218
rect 298794 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 299414 552134
rect 298794 516454 299414 551898
rect 298794 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 299414 516454
rect 298794 516134 299414 516218
rect 298794 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 299414 516134
rect 298794 480454 299414 515898
rect 298794 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 299414 480454
rect 298794 480134 299414 480218
rect 298794 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 299414 480134
rect 298794 444454 299414 479898
rect 298794 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 299414 444454
rect 298794 444134 299414 444218
rect 298794 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 299414 444134
rect 298794 408454 299414 443898
rect 298794 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 299414 408454
rect 298794 408134 299414 408218
rect 298794 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 299414 408134
rect 298794 372454 299414 407898
rect 298794 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 299414 372454
rect 298794 372134 299414 372218
rect 298794 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 299414 372134
rect 298794 336454 299414 371898
rect 298794 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 299414 336454
rect 298794 336134 299414 336218
rect 298794 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 299414 336134
rect 298794 300454 299414 335898
rect 298794 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 299414 300454
rect 298794 300134 299414 300218
rect 298794 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 299414 300134
rect 298794 264454 299414 299898
rect 298794 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 299414 264454
rect 298794 264134 299414 264218
rect 298794 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 299414 264134
rect 298794 248684 299414 263898
rect 303294 707718 303914 711590
rect 303294 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 303914 707718
rect 303294 707398 303914 707482
rect 303294 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 303914 707398
rect 303294 700954 303914 707162
rect 303294 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 303914 700954
rect 303294 700634 303914 700718
rect 303294 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 303914 700634
rect 303294 664954 303914 700398
rect 303294 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 303914 664954
rect 303294 664634 303914 664718
rect 303294 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 303914 664634
rect 303294 628954 303914 664398
rect 303294 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 303914 628954
rect 303294 628634 303914 628718
rect 303294 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 303914 628634
rect 303294 592954 303914 628398
rect 303294 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 303914 592954
rect 303294 592634 303914 592718
rect 303294 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 303914 592634
rect 303294 556954 303914 592398
rect 303294 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 303914 556954
rect 303294 556634 303914 556718
rect 303294 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 303914 556634
rect 303294 520954 303914 556398
rect 303294 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 303914 520954
rect 303294 520634 303914 520718
rect 303294 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 303914 520634
rect 303294 484954 303914 520398
rect 303294 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 303914 484954
rect 303294 484634 303914 484718
rect 303294 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 303914 484634
rect 303294 448954 303914 484398
rect 303294 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 303914 448954
rect 303294 448634 303914 448718
rect 303294 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 303914 448634
rect 303294 412954 303914 448398
rect 303294 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 303914 412954
rect 303294 412634 303914 412718
rect 303294 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 303914 412634
rect 303294 376954 303914 412398
rect 303294 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 303914 376954
rect 303294 376634 303914 376718
rect 303294 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 303914 376634
rect 303294 340954 303914 376398
rect 303294 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 303914 340954
rect 303294 340634 303914 340718
rect 303294 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 303914 340634
rect 303294 304954 303914 340398
rect 303294 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 303914 304954
rect 303294 304634 303914 304718
rect 303294 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 303914 304634
rect 303294 268954 303914 304398
rect 303294 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 303914 268954
rect 303294 268634 303914 268718
rect 303294 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 303914 268634
rect 303294 248684 303914 268398
rect 307794 708678 308414 711590
rect 307794 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 308414 708678
rect 307794 708358 308414 708442
rect 307794 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 308414 708358
rect 307794 669454 308414 708122
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 248684 308414 272898
rect 312294 709638 312914 711590
rect 312294 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 312914 709638
rect 312294 709318 312914 709402
rect 312294 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 312914 709318
rect 312294 673954 312914 709082
rect 312294 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 312914 673954
rect 312294 673634 312914 673718
rect 312294 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 312914 673634
rect 312294 637954 312914 673398
rect 312294 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 312914 637954
rect 312294 637634 312914 637718
rect 312294 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 312914 637634
rect 312294 601954 312914 637398
rect 312294 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 312914 601954
rect 312294 601634 312914 601718
rect 312294 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 312914 601634
rect 312294 565954 312914 601398
rect 312294 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 312914 565954
rect 312294 565634 312914 565718
rect 312294 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 312914 565634
rect 312294 529954 312914 565398
rect 312294 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 312914 529954
rect 312294 529634 312914 529718
rect 312294 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 312914 529634
rect 312294 493954 312914 529398
rect 312294 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 312914 493954
rect 312294 493634 312914 493718
rect 312294 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 312914 493634
rect 312294 457954 312914 493398
rect 312294 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 312914 457954
rect 312294 457634 312914 457718
rect 312294 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 312914 457634
rect 312294 421954 312914 457398
rect 312294 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 312914 421954
rect 312294 421634 312914 421718
rect 312294 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 312914 421634
rect 312294 385954 312914 421398
rect 312294 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 312914 385954
rect 312294 385634 312914 385718
rect 312294 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 312914 385634
rect 312294 349954 312914 385398
rect 312294 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 312914 349954
rect 312294 349634 312914 349718
rect 312294 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 312914 349634
rect 312294 313954 312914 349398
rect 312294 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 312914 313954
rect 312294 313634 312914 313718
rect 312294 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 312914 313634
rect 312294 277954 312914 313398
rect 312294 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 312914 277954
rect 312294 277634 312914 277718
rect 312294 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 312914 277634
rect 312294 248684 312914 277398
rect 316794 710598 317414 711590
rect 316794 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 317414 710598
rect 316794 710278 317414 710362
rect 316794 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 317414 710278
rect 316794 678454 317414 710042
rect 316794 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 317414 678454
rect 316794 678134 317414 678218
rect 316794 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 317414 678134
rect 316794 642454 317414 677898
rect 316794 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 317414 642454
rect 316794 642134 317414 642218
rect 316794 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 317414 642134
rect 316794 606454 317414 641898
rect 316794 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 317414 606454
rect 316794 606134 317414 606218
rect 316794 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 317414 606134
rect 316794 570454 317414 605898
rect 316794 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 317414 570454
rect 316794 570134 317414 570218
rect 316794 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 317414 570134
rect 316794 534454 317414 569898
rect 316794 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 317414 534454
rect 316794 534134 317414 534218
rect 316794 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 317414 534134
rect 316794 498454 317414 533898
rect 316794 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 317414 498454
rect 316794 498134 317414 498218
rect 316794 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 317414 498134
rect 316794 462454 317414 497898
rect 316794 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 317414 462454
rect 316794 462134 317414 462218
rect 316794 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 317414 462134
rect 316794 426454 317414 461898
rect 316794 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 317414 426454
rect 316794 426134 317414 426218
rect 316794 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 317414 426134
rect 316794 390454 317414 425898
rect 316794 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 317414 390454
rect 316794 390134 317414 390218
rect 316794 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 317414 390134
rect 316794 354454 317414 389898
rect 316794 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 317414 354454
rect 316794 354134 317414 354218
rect 316794 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 317414 354134
rect 316794 318454 317414 353898
rect 316794 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 317414 318454
rect 316794 318134 317414 318218
rect 316794 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 317414 318134
rect 316794 282454 317414 317898
rect 316794 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 317414 282454
rect 316794 282134 317414 282218
rect 316794 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 317414 282134
rect 316794 248684 317414 281898
rect 321294 711558 321914 711590
rect 321294 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 321914 711558
rect 321294 711238 321914 711322
rect 321294 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 321914 711238
rect 321294 682954 321914 711002
rect 321294 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 321914 682954
rect 321294 682634 321914 682718
rect 321294 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 321914 682634
rect 321294 646954 321914 682398
rect 321294 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 321914 646954
rect 321294 646634 321914 646718
rect 321294 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 321914 646634
rect 321294 610954 321914 646398
rect 321294 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 321914 610954
rect 321294 610634 321914 610718
rect 321294 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 321914 610634
rect 321294 574954 321914 610398
rect 321294 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 321914 574954
rect 321294 574634 321914 574718
rect 321294 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 321914 574634
rect 321294 538954 321914 574398
rect 321294 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 321914 538954
rect 321294 538634 321914 538718
rect 321294 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 321914 538634
rect 321294 502954 321914 538398
rect 321294 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 321914 502954
rect 321294 502634 321914 502718
rect 321294 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 321914 502634
rect 321294 466954 321914 502398
rect 321294 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 321914 466954
rect 321294 466634 321914 466718
rect 321294 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 321914 466634
rect 321294 430954 321914 466398
rect 321294 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 321914 430954
rect 321294 430634 321914 430718
rect 321294 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 321914 430634
rect 321294 394954 321914 430398
rect 321294 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 321914 394954
rect 321294 394634 321914 394718
rect 321294 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 321914 394634
rect 321294 358954 321914 394398
rect 321294 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 321914 358954
rect 321294 358634 321914 358718
rect 321294 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 321914 358634
rect 321294 322954 321914 358398
rect 321294 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 321914 322954
rect 321294 322634 321914 322718
rect 321294 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 321914 322634
rect 321294 286954 321914 322398
rect 321294 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 321914 286954
rect 321294 286634 321914 286718
rect 321294 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 321914 286634
rect 321294 250954 321914 286398
rect 321294 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 321914 250954
rect 321294 250634 321914 250718
rect 321294 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 321914 250634
rect 321294 248684 321914 250398
rect 325794 704838 326414 711590
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 248684 326414 254898
rect 330294 705798 330914 711590
rect 330294 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 330914 705798
rect 330294 705478 330914 705562
rect 330294 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 330914 705478
rect 330294 691954 330914 705242
rect 330294 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 330914 691954
rect 330294 691634 330914 691718
rect 330294 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 330914 691634
rect 330294 655954 330914 691398
rect 330294 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 330914 655954
rect 330294 655634 330914 655718
rect 330294 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 330914 655634
rect 330294 619954 330914 655398
rect 330294 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 330914 619954
rect 330294 619634 330914 619718
rect 330294 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 330914 619634
rect 330294 583954 330914 619398
rect 330294 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 330914 583954
rect 330294 583634 330914 583718
rect 330294 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 330914 583634
rect 330294 547954 330914 583398
rect 330294 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 330914 547954
rect 330294 547634 330914 547718
rect 330294 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 330914 547634
rect 330294 511954 330914 547398
rect 330294 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 330914 511954
rect 330294 511634 330914 511718
rect 330294 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 330914 511634
rect 330294 475954 330914 511398
rect 330294 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 330914 475954
rect 330294 475634 330914 475718
rect 330294 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 330914 475634
rect 330294 439954 330914 475398
rect 330294 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 330914 439954
rect 330294 439634 330914 439718
rect 330294 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 330914 439634
rect 330294 403954 330914 439398
rect 330294 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 330914 403954
rect 330294 403634 330914 403718
rect 330294 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 330914 403634
rect 330294 367954 330914 403398
rect 330294 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 330914 367954
rect 330294 367634 330914 367718
rect 330294 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 330914 367634
rect 330294 331954 330914 367398
rect 330294 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 330914 331954
rect 330294 331634 330914 331718
rect 330294 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 330914 331634
rect 330294 295954 330914 331398
rect 330294 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 330914 295954
rect 330294 295634 330914 295718
rect 330294 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 330914 295634
rect 330294 259954 330914 295398
rect 330294 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 330914 259954
rect 330294 259634 330914 259718
rect 330294 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 330914 259634
rect 330294 248684 330914 259398
rect 334794 706758 335414 711590
rect 334794 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 335414 706758
rect 334794 706438 335414 706522
rect 334794 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 335414 706438
rect 334794 696454 335414 706202
rect 334794 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 335414 696454
rect 334794 696134 335414 696218
rect 334794 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 335414 696134
rect 334794 660454 335414 695898
rect 334794 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 335414 660454
rect 334794 660134 335414 660218
rect 334794 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 335414 660134
rect 334794 624454 335414 659898
rect 334794 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 335414 624454
rect 334794 624134 335414 624218
rect 334794 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 335414 624134
rect 334794 588454 335414 623898
rect 334794 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 335414 588454
rect 334794 588134 335414 588218
rect 334794 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 335414 588134
rect 334794 552454 335414 587898
rect 334794 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 335414 552454
rect 334794 552134 335414 552218
rect 334794 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 335414 552134
rect 334794 516454 335414 551898
rect 334794 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 335414 516454
rect 334794 516134 335414 516218
rect 334794 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 335414 516134
rect 334794 480454 335414 515898
rect 334794 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 335414 480454
rect 334794 480134 335414 480218
rect 334794 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 335414 480134
rect 334794 444454 335414 479898
rect 334794 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 335414 444454
rect 334794 444134 335414 444218
rect 334794 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 335414 444134
rect 334794 408454 335414 443898
rect 334794 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 335414 408454
rect 334794 408134 335414 408218
rect 334794 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 335414 408134
rect 334794 372454 335414 407898
rect 334794 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 335414 372454
rect 334794 372134 335414 372218
rect 334794 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 335414 372134
rect 334794 336454 335414 371898
rect 334794 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 335414 336454
rect 334794 336134 335414 336218
rect 334794 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 335414 336134
rect 334794 300454 335414 335898
rect 334794 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 335414 300454
rect 334794 300134 335414 300218
rect 334794 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 335414 300134
rect 334794 264454 335414 299898
rect 334794 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 335414 264454
rect 334794 264134 335414 264218
rect 334794 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 335414 264134
rect 334794 248684 335414 263898
rect 339294 707718 339914 711590
rect 339294 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 339914 707718
rect 339294 707398 339914 707482
rect 339294 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 339914 707398
rect 339294 700954 339914 707162
rect 339294 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 339914 700954
rect 339294 700634 339914 700718
rect 339294 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 339914 700634
rect 339294 664954 339914 700398
rect 339294 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 339914 664954
rect 339294 664634 339914 664718
rect 339294 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 339914 664634
rect 339294 628954 339914 664398
rect 339294 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 339914 628954
rect 339294 628634 339914 628718
rect 339294 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 339914 628634
rect 339294 592954 339914 628398
rect 339294 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 339914 592954
rect 339294 592634 339914 592718
rect 339294 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 339914 592634
rect 339294 556954 339914 592398
rect 339294 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 339914 556954
rect 339294 556634 339914 556718
rect 339294 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 339914 556634
rect 339294 520954 339914 556398
rect 339294 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 339914 520954
rect 339294 520634 339914 520718
rect 339294 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 339914 520634
rect 339294 484954 339914 520398
rect 339294 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 339914 484954
rect 339294 484634 339914 484718
rect 339294 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 339914 484634
rect 339294 448954 339914 484398
rect 339294 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 339914 448954
rect 339294 448634 339914 448718
rect 339294 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 339914 448634
rect 339294 412954 339914 448398
rect 339294 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 339914 412954
rect 339294 412634 339914 412718
rect 339294 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 339914 412634
rect 339294 376954 339914 412398
rect 339294 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 339914 376954
rect 339294 376634 339914 376718
rect 339294 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 339914 376634
rect 339294 340954 339914 376398
rect 339294 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 339914 340954
rect 339294 340634 339914 340718
rect 339294 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 339914 340634
rect 339294 304954 339914 340398
rect 339294 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 339914 304954
rect 339294 304634 339914 304718
rect 339294 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 339914 304634
rect 339294 268954 339914 304398
rect 339294 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 339914 268954
rect 339294 268634 339914 268718
rect 339294 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 339914 268634
rect 339294 248684 339914 268398
rect 343794 708678 344414 711590
rect 343794 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 344414 708678
rect 343794 708358 344414 708442
rect 343794 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 344414 708358
rect 343794 669454 344414 708122
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 248684 344414 272898
rect 348294 709638 348914 711590
rect 348294 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 348914 709638
rect 348294 709318 348914 709402
rect 348294 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 348914 709318
rect 348294 673954 348914 709082
rect 348294 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 348914 673954
rect 348294 673634 348914 673718
rect 348294 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 348914 673634
rect 348294 637954 348914 673398
rect 348294 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 348914 637954
rect 348294 637634 348914 637718
rect 348294 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 348914 637634
rect 348294 601954 348914 637398
rect 348294 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 348914 601954
rect 348294 601634 348914 601718
rect 348294 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 348914 601634
rect 348294 565954 348914 601398
rect 348294 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 348914 565954
rect 348294 565634 348914 565718
rect 348294 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 348914 565634
rect 348294 529954 348914 565398
rect 348294 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 348914 529954
rect 348294 529634 348914 529718
rect 348294 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 348914 529634
rect 348294 493954 348914 529398
rect 348294 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 348914 493954
rect 348294 493634 348914 493718
rect 348294 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 348914 493634
rect 348294 457954 348914 493398
rect 348294 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 348914 457954
rect 348294 457634 348914 457718
rect 348294 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 348914 457634
rect 348294 421954 348914 457398
rect 348294 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 348914 421954
rect 348294 421634 348914 421718
rect 348294 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 348914 421634
rect 348294 385954 348914 421398
rect 348294 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 348914 385954
rect 348294 385634 348914 385718
rect 348294 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 348914 385634
rect 348294 349954 348914 385398
rect 348294 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 348914 349954
rect 348294 349634 348914 349718
rect 348294 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 348914 349634
rect 348294 313954 348914 349398
rect 348294 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 348914 313954
rect 348294 313634 348914 313718
rect 348294 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 348914 313634
rect 348294 277954 348914 313398
rect 348294 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 348914 277954
rect 348294 277634 348914 277718
rect 348294 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 348914 277634
rect 348294 248684 348914 277398
rect 352794 710598 353414 711590
rect 352794 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 353414 710598
rect 352794 710278 353414 710362
rect 352794 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 353414 710278
rect 352794 678454 353414 710042
rect 352794 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 353414 678454
rect 352794 678134 353414 678218
rect 352794 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 353414 678134
rect 352794 642454 353414 677898
rect 352794 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 353414 642454
rect 352794 642134 353414 642218
rect 352794 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 353414 642134
rect 352794 606454 353414 641898
rect 352794 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 353414 606454
rect 352794 606134 353414 606218
rect 352794 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 353414 606134
rect 352794 570454 353414 605898
rect 352794 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 353414 570454
rect 352794 570134 353414 570218
rect 352794 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 353414 570134
rect 352794 534454 353414 569898
rect 352794 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 353414 534454
rect 352794 534134 353414 534218
rect 352794 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 353414 534134
rect 352794 498454 353414 533898
rect 352794 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 353414 498454
rect 352794 498134 353414 498218
rect 352794 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 353414 498134
rect 352794 462454 353414 497898
rect 352794 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 353414 462454
rect 352794 462134 353414 462218
rect 352794 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 353414 462134
rect 352794 426454 353414 461898
rect 352794 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 353414 426454
rect 352794 426134 353414 426218
rect 352794 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 353414 426134
rect 352794 390454 353414 425898
rect 352794 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 353414 390454
rect 352794 390134 353414 390218
rect 352794 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 353414 390134
rect 352794 354454 353414 389898
rect 352794 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 353414 354454
rect 352794 354134 353414 354218
rect 352794 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 353414 354134
rect 352794 318454 353414 353898
rect 352794 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 353414 318454
rect 352794 318134 353414 318218
rect 352794 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 353414 318134
rect 352794 282454 353414 317898
rect 352794 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 353414 282454
rect 352794 282134 353414 282218
rect 352794 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 353414 282134
rect 352794 248684 353414 281898
rect 357294 711558 357914 711590
rect 357294 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 357914 711558
rect 357294 711238 357914 711322
rect 357294 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 357914 711238
rect 357294 682954 357914 711002
rect 357294 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 357914 682954
rect 357294 682634 357914 682718
rect 357294 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 357914 682634
rect 357294 646954 357914 682398
rect 357294 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 357914 646954
rect 357294 646634 357914 646718
rect 357294 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 357914 646634
rect 357294 610954 357914 646398
rect 357294 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 357914 610954
rect 357294 610634 357914 610718
rect 357294 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 357914 610634
rect 357294 574954 357914 610398
rect 357294 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 357914 574954
rect 357294 574634 357914 574718
rect 357294 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 357914 574634
rect 357294 538954 357914 574398
rect 357294 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 357914 538954
rect 357294 538634 357914 538718
rect 357294 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 357914 538634
rect 357294 502954 357914 538398
rect 357294 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 357914 502954
rect 357294 502634 357914 502718
rect 357294 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 357914 502634
rect 357294 466954 357914 502398
rect 357294 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 357914 466954
rect 357294 466634 357914 466718
rect 357294 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 357914 466634
rect 357294 430954 357914 466398
rect 357294 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 357914 430954
rect 357294 430634 357914 430718
rect 357294 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 357914 430634
rect 357294 394954 357914 430398
rect 357294 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 357914 394954
rect 357294 394634 357914 394718
rect 357294 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 357914 394634
rect 357294 358954 357914 394398
rect 357294 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 357914 358954
rect 357294 358634 357914 358718
rect 357294 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 357914 358634
rect 357294 322954 357914 358398
rect 357294 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 357914 322954
rect 357294 322634 357914 322718
rect 357294 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 357914 322634
rect 357294 286954 357914 322398
rect 357294 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 357914 286954
rect 357294 286634 357914 286718
rect 357294 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 357914 286634
rect 357294 250954 357914 286398
rect 357294 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 357914 250954
rect 357294 250634 357914 250718
rect 357294 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 357914 250634
rect 357294 248684 357914 250398
rect 361794 704838 362414 711590
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 248684 362414 254898
rect 366294 705798 366914 711590
rect 366294 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 366914 705798
rect 366294 705478 366914 705562
rect 366294 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 366914 705478
rect 366294 691954 366914 705242
rect 366294 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 366914 691954
rect 366294 691634 366914 691718
rect 366294 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 366914 691634
rect 366294 655954 366914 691398
rect 366294 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 366914 655954
rect 366294 655634 366914 655718
rect 366294 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 366914 655634
rect 366294 619954 366914 655398
rect 366294 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 366914 619954
rect 366294 619634 366914 619718
rect 366294 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 366914 619634
rect 366294 583954 366914 619398
rect 366294 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 366914 583954
rect 366294 583634 366914 583718
rect 366294 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 366914 583634
rect 366294 547954 366914 583398
rect 366294 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 366914 547954
rect 366294 547634 366914 547718
rect 366294 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 366914 547634
rect 366294 511954 366914 547398
rect 366294 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 366914 511954
rect 366294 511634 366914 511718
rect 366294 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 366914 511634
rect 366294 475954 366914 511398
rect 366294 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 366914 475954
rect 366294 475634 366914 475718
rect 366294 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 366914 475634
rect 366294 439954 366914 475398
rect 366294 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 366914 439954
rect 366294 439634 366914 439718
rect 366294 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 366914 439634
rect 366294 403954 366914 439398
rect 366294 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 366914 403954
rect 366294 403634 366914 403718
rect 366294 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 366914 403634
rect 366294 367954 366914 403398
rect 366294 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 366914 367954
rect 366294 367634 366914 367718
rect 366294 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 366914 367634
rect 366294 331954 366914 367398
rect 366294 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 366914 331954
rect 366294 331634 366914 331718
rect 366294 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 366914 331634
rect 366294 295954 366914 331398
rect 366294 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 366914 295954
rect 366294 295634 366914 295718
rect 366294 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 366914 295634
rect 366294 259954 366914 295398
rect 366294 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 366914 259954
rect 366294 259634 366914 259718
rect 366294 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 366914 259634
rect 366294 248684 366914 259398
rect 370794 706758 371414 711590
rect 370794 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 371414 706758
rect 370794 706438 371414 706522
rect 370794 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 371414 706438
rect 370794 696454 371414 706202
rect 370794 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 371414 696454
rect 370794 696134 371414 696218
rect 370794 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 371414 696134
rect 370794 660454 371414 695898
rect 370794 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 371414 660454
rect 370794 660134 371414 660218
rect 370794 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 371414 660134
rect 370794 624454 371414 659898
rect 370794 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 371414 624454
rect 370794 624134 371414 624218
rect 370794 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 371414 624134
rect 370794 588454 371414 623898
rect 370794 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 371414 588454
rect 370794 588134 371414 588218
rect 370794 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 371414 588134
rect 370794 552454 371414 587898
rect 370794 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 371414 552454
rect 370794 552134 371414 552218
rect 370794 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 371414 552134
rect 370794 516454 371414 551898
rect 370794 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 371414 516454
rect 370794 516134 371414 516218
rect 370794 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 371414 516134
rect 370794 480454 371414 515898
rect 370794 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 371414 480454
rect 370794 480134 371414 480218
rect 370794 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 371414 480134
rect 370794 444454 371414 479898
rect 370794 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 371414 444454
rect 370794 444134 371414 444218
rect 370794 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 371414 444134
rect 370794 408454 371414 443898
rect 370794 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 371414 408454
rect 370794 408134 371414 408218
rect 370794 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 371414 408134
rect 370794 372454 371414 407898
rect 370794 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 371414 372454
rect 370794 372134 371414 372218
rect 370794 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 371414 372134
rect 370794 336454 371414 371898
rect 370794 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 371414 336454
rect 370794 336134 371414 336218
rect 370794 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 371414 336134
rect 370794 300454 371414 335898
rect 370794 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 371414 300454
rect 370794 300134 371414 300218
rect 370794 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 371414 300134
rect 370794 264454 371414 299898
rect 370794 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 371414 264454
rect 370794 264134 371414 264218
rect 370794 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 371414 264134
rect 370794 248684 371414 263898
rect 375294 707718 375914 711590
rect 375294 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 375914 707718
rect 375294 707398 375914 707482
rect 375294 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 375914 707398
rect 375294 700954 375914 707162
rect 375294 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 375914 700954
rect 375294 700634 375914 700718
rect 375294 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 375914 700634
rect 375294 664954 375914 700398
rect 375294 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 375914 664954
rect 375294 664634 375914 664718
rect 375294 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 375914 664634
rect 375294 628954 375914 664398
rect 375294 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 375914 628954
rect 375294 628634 375914 628718
rect 375294 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 375914 628634
rect 375294 592954 375914 628398
rect 375294 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 375914 592954
rect 375294 592634 375914 592718
rect 375294 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 375914 592634
rect 375294 556954 375914 592398
rect 375294 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 375914 556954
rect 375294 556634 375914 556718
rect 375294 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 375914 556634
rect 375294 520954 375914 556398
rect 375294 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 375914 520954
rect 375294 520634 375914 520718
rect 375294 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 375914 520634
rect 375294 484954 375914 520398
rect 375294 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 375914 484954
rect 375294 484634 375914 484718
rect 375294 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 375914 484634
rect 375294 448954 375914 484398
rect 375294 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 375914 448954
rect 375294 448634 375914 448718
rect 375294 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 375914 448634
rect 375294 412954 375914 448398
rect 375294 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 375914 412954
rect 375294 412634 375914 412718
rect 375294 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 375914 412634
rect 375294 376954 375914 412398
rect 375294 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 375914 376954
rect 375294 376634 375914 376718
rect 375294 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 375914 376634
rect 375294 340954 375914 376398
rect 375294 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 375914 340954
rect 375294 340634 375914 340718
rect 375294 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 375914 340634
rect 375294 304954 375914 340398
rect 375294 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 375914 304954
rect 375294 304634 375914 304718
rect 375294 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 375914 304634
rect 375294 268954 375914 304398
rect 375294 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 375914 268954
rect 375294 268634 375914 268718
rect 375294 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 375914 268634
rect 375294 248684 375914 268398
rect 379794 708678 380414 711590
rect 379794 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 380414 708678
rect 379794 708358 380414 708442
rect 379794 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 380414 708358
rect 379794 669454 380414 708122
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 248684 380414 272898
rect 384294 709638 384914 711590
rect 384294 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 384914 709638
rect 384294 709318 384914 709402
rect 384294 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 384914 709318
rect 384294 673954 384914 709082
rect 384294 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 384914 673954
rect 384294 673634 384914 673718
rect 384294 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 384914 673634
rect 384294 637954 384914 673398
rect 384294 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 384914 637954
rect 384294 637634 384914 637718
rect 384294 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 384914 637634
rect 384294 601954 384914 637398
rect 384294 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 384914 601954
rect 384294 601634 384914 601718
rect 384294 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 384914 601634
rect 384294 565954 384914 601398
rect 384294 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 384914 565954
rect 384294 565634 384914 565718
rect 384294 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 384914 565634
rect 384294 529954 384914 565398
rect 384294 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 384914 529954
rect 384294 529634 384914 529718
rect 384294 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 384914 529634
rect 384294 493954 384914 529398
rect 384294 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 384914 493954
rect 384294 493634 384914 493718
rect 384294 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 384914 493634
rect 384294 457954 384914 493398
rect 384294 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 384914 457954
rect 384294 457634 384914 457718
rect 384294 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 384914 457634
rect 384294 421954 384914 457398
rect 384294 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 384914 421954
rect 384294 421634 384914 421718
rect 384294 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 384914 421634
rect 384294 385954 384914 421398
rect 384294 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 384914 385954
rect 384294 385634 384914 385718
rect 384294 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 384914 385634
rect 384294 349954 384914 385398
rect 384294 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 384914 349954
rect 384294 349634 384914 349718
rect 384294 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 384914 349634
rect 384294 313954 384914 349398
rect 384294 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 384914 313954
rect 384294 313634 384914 313718
rect 384294 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 384914 313634
rect 384294 277954 384914 313398
rect 384294 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 384914 277954
rect 384294 277634 384914 277718
rect 384294 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 384914 277634
rect 384294 248684 384914 277398
rect 388794 710598 389414 711590
rect 388794 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 389414 710598
rect 388794 710278 389414 710362
rect 388794 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 389414 710278
rect 388794 678454 389414 710042
rect 388794 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 389414 678454
rect 388794 678134 389414 678218
rect 388794 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 389414 678134
rect 388794 642454 389414 677898
rect 388794 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 389414 642454
rect 388794 642134 389414 642218
rect 388794 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 389414 642134
rect 388794 606454 389414 641898
rect 388794 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 389414 606454
rect 388794 606134 389414 606218
rect 388794 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 389414 606134
rect 388794 570454 389414 605898
rect 388794 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 389414 570454
rect 388794 570134 389414 570218
rect 388794 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 389414 570134
rect 388794 534454 389414 569898
rect 388794 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 389414 534454
rect 388794 534134 389414 534218
rect 388794 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 389414 534134
rect 388794 498454 389414 533898
rect 388794 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 389414 498454
rect 388794 498134 389414 498218
rect 388794 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 389414 498134
rect 388794 462454 389414 497898
rect 388794 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 389414 462454
rect 388794 462134 389414 462218
rect 388794 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 389414 462134
rect 388794 426454 389414 461898
rect 388794 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 389414 426454
rect 388794 426134 389414 426218
rect 388794 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 389414 426134
rect 388794 390454 389414 425898
rect 388794 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 389414 390454
rect 388794 390134 389414 390218
rect 388794 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 389414 390134
rect 388794 354454 389414 389898
rect 388794 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 389414 354454
rect 388794 354134 389414 354218
rect 388794 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 389414 354134
rect 388794 318454 389414 353898
rect 388794 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 389414 318454
rect 388794 318134 389414 318218
rect 388794 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 389414 318134
rect 388794 282454 389414 317898
rect 388794 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 389414 282454
rect 388794 282134 389414 282218
rect 388794 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 389414 282134
rect 388794 248684 389414 281898
rect 393294 711558 393914 711590
rect 393294 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 393914 711558
rect 393294 711238 393914 711322
rect 393294 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 393914 711238
rect 393294 682954 393914 711002
rect 393294 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 393914 682954
rect 393294 682634 393914 682718
rect 393294 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 393914 682634
rect 393294 646954 393914 682398
rect 393294 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 393914 646954
rect 393294 646634 393914 646718
rect 393294 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 393914 646634
rect 393294 610954 393914 646398
rect 393294 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 393914 610954
rect 393294 610634 393914 610718
rect 393294 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 393914 610634
rect 393294 574954 393914 610398
rect 393294 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 393914 574954
rect 393294 574634 393914 574718
rect 393294 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 393914 574634
rect 393294 538954 393914 574398
rect 393294 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 393914 538954
rect 393294 538634 393914 538718
rect 393294 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 393914 538634
rect 393294 502954 393914 538398
rect 393294 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 393914 502954
rect 393294 502634 393914 502718
rect 393294 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 393914 502634
rect 393294 466954 393914 502398
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 396579 470660 396645 470661
rect 396579 470596 396580 470660
rect 396644 470596 396645 470660
rect 396579 470595 396645 470596
rect 393294 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 393914 466954
rect 393294 466634 393914 466718
rect 393294 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 393914 466634
rect 393294 430954 393914 466398
rect 393294 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 393914 430954
rect 393294 430634 393914 430718
rect 393294 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 393914 430634
rect 393294 394954 393914 430398
rect 393294 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 393914 394954
rect 393294 394634 393914 394718
rect 393294 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 393914 394634
rect 393294 358954 393914 394398
rect 393294 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 393914 358954
rect 393294 358634 393914 358718
rect 393294 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 393914 358634
rect 393294 322954 393914 358398
rect 393294 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 393914 322954
rect 393294 322634 393914 322718
rect 393294 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 393914 322634
rect 393294 286954 393914 322398
rect 393294 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 393914 286954
rect 393294 286634 393914 286718
rect 393294 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 393914 286634
rect 393294 250954 393914 286398
rect 393294 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 393914 250954
rect 393294 250634 393914 250718
rect 393294 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 393914 250634
rect 393294 248684 393914 250398
rect 65300 246303 70100 246486
rect 65300 246067 65342 246303
rect 65578 246067 65662 246303
rect 65898 246067 65982 246303
rect 66218 246067 66302 246303
rect 66538 246067 66622 246303
rect 66858 246067 66942 246303
rect 67178 246067 67262 246303
rect 67498 246067 67582 246303
rect 67818 246067 67902 246303
rect 68138 246067 68222 246303
rect 68458 246067 68542 246303
rect 68778 246067 68862 246303
rect 69098 246067 69182 246303
rect 69418 246067 69502 246303
rect 69738 246067 69822 246303
rect 70058 246067 70100 246303
rect 65300 245884 70100 246067
rect 65300 241953 71300 241984
rect 65300 241717 65462 241953
rect 65698 241717 65782 241953
rect 66018 241717 66102 241953
rect 66338 241717 66422 241953
rect 66658 241717 66742 241953
rect 66978 241717 67062 241953
rect 67298 241717 67382 241953
rect 67618 241717 67702 241953
rect 67938 241717 68022 241953
rect 68258 241717 68342 241953
rect 68578 241717 68662 241953
rect 68898 241717 68982 241953
rect 69218 241717 69302 241953
rect 69538 241717 69622 241953
rect 69858 241717 69942 241953
rect 70178 241717 70262 241953
rect 70498 241717 70582 241953
rect 70818 241717 70902 241953
rect 71138 241717 71300 241953
rect 65300 241633 71300 241717
rect 65300 241397 65462 241633
rect 65698 241397 65782 241633
rect 66018 241397 66102 241633
rect 66338 241397 66422 241633
rect 66658 241397 66742 241633
rect 66978 241397 67062 241633
rect 67298 241397 67382 241633
rect 67618 241397 67702 241633
rect 67938 241397 68022 241633
rect 68258 241397 68342 241633
rect 68578 241397 68662 241633
rect 68898 241397 68982 241633
rect 69218 241397 69302 241633
rect 69538 241397 69622 241633
rect 69858 241397 69942 241633
rect 70178 241397 70262 241633
rect 70498 241397 70582 241633
rect 70818 241397 70902 241633
rect 71138 241397 71300 241633
rect 65300 241366 71300 241397
rect 42294 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 42914 223954
rect 42294 223634 42914 223718
rect 42294 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 42914 223634
rect 42294 187954 42914 223398
rect 42294 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 42914 187954
rect 42294 187634 42914 187718
rect 42294 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 42914 187634
rect 42294 151954 42914 187398
rect 42294 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 42914 151954
rect 42294 151634 42914 151718
rect 42294 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 42914 151634
rect 42294 115954 42914 151398
rect 42294 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 42914 115954
rect 42294 115634 42914 115718
rect 42294 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 42914 115634
rect 42294 79954 42914 115398
rect 42294 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 42914 79954
rect 42294 79634 42914 79718
rect 42294 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 42914 79634
rect 42294 43954 42914 79398
rect 42294 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 42914 43954
rect 42294 43634 42914 43718
rect 42294 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 42914 43634
rect 42294 7954 42914 43398
rect 42294 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 42914 7954
rect 42294 7634 42914 7718
rect 42294 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 42914 7634
rect 42294 -1306 42914 7398
rect 42294 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 42914 -1306
rect 42294 -1626 42914 -1542
rect 42294 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 42914 -1626
rect 42294 -7654 42914 -1862
rect 46794 228453 47414 228484
rect 46794 228217 46826 228453
rect 47062 228217 47146 228453
rect 47382 228217 47414 228453
rect 46794 228133 47414 228217
rect 46794 227897 46826 228133
rect 47062 227897 47146 228133
rect 47382 227897 47414 228133
rect 46794 192454 47414 227897
rect 46794 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 47414 192454
rect 46794 192134 47414 192218
rect 46794 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 47414 192134
rect 46794 156454 47414 191898
rect 46794 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 47414 156454
rect 46794 156134 47414 156218
rect 46794 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 47414 156134
rect 46794 120454 47414 155898
rect 46794 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 47414 120454
rect 46794 120134 47414 120218
rect 46794 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 47414 120134
rect 46794 84454 47414 119898
rect 46794 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 47414 84454
rect 46794 84134 47414 84218
rect 46794 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 47414 84134
rect 46794 48454 47414 83898
rect 46794 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 47414 48454
rect 46794 48134 47414 48218
rect 46794 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 47414 48134
rect 46794 12454 47414 47898
rect 46794 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 47414 12454
rect 46794 12134 47414 12218
rect 46794 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 47414 12134
rect 46794 -2266 47414 11898
rect 46794 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 47414 -2266
rect 46794 -2586 47414 -2502
rect 46794 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 47414 -2586
rect 46794 -7654 47414 -2822
rect 51294 196954 51914 228484
rect 51294 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 51914 196954
rect 51294 196634 51914 196718
rect 51294 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 51914 196634
rect 51294 160954 51914 196398
rect 51294 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 51914 160954
rect 51294 160634 51914 160718
rect 51294 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 51914 160634
rect 51294 124954 51914 160398
rect 51294 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 51914 124954
rect 51294 124634 51914 124718
rect 51294 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 51914 124634
rect 51294 88954 51914 124398
rect 51294 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 51914 88954
rect 51294 88634 51914 88718
rect 51294 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 51914 88634
rect 51294 52954 51914 88398
rect 51294 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 51914 52954
rect 51294 52634 51914 52718
rect 51294 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 51914 52634
rect 51294 16954 51914 52398
rect 51294 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 51914 16954
rect 51294 16634 51914 16718
rect 51294 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 51914 16634
rect 51294 -3226 51914 16398
rect 51294 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 51914 -3226
rect 51294 -3546 51914 -3462
rect 51294 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 51914 -3546
rect 51294 -7654 51914 -3782
rect 55794 201454 56414 228484
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -4186 56414 20898
rect 55794 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 56414 -4186
rect 55794 -4506 56414 -4422
rect 55794 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 56414 -4506
rect 55794 -7654 56414 -4742
rect 60294 205954 60914 228484
rect 60294 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 60914 205954
rect 60294 205634 60914 205718
rect 60294 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 60914 205634
rect 60294 169954 60914 205398
rect 60294 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 60914 169954
rect 60294 169634 60914 169718
rect 60294 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 60914 169634
rect 60294 133954 60914 169398
rect 60294 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 60914 133954
rect 60294 133634 60914 133718
rect 60294 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 60914 133634
rect 60294 97954 60914 133398
rect 60294 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 60914 97954
rect 60294 97634 60914 97718
rect 60294 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 60914 97634
rect 60294 61954 60914 97398
rect 60294 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 60914 61954
rect 60294 61634 60914 61718
rect 60294 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 60914 61634
rect 60294 25954 60914 61398
rect 60294 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 60914 25954
rect 60294 25634 60914 25718
rect 60294 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 60914 25634
rect 60294 -5146 60914 25398
rect 60294 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 60914 -5146
rect 60294 -5466 60914 -5382
rect 60294 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 60914 -5466
rect 60294 -7654 60914 -5702
rect 64794 210454 65414 228484
rect 64794 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 65414 210454
rect 64794 210134 65414 210218
rect 64794 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 65414 210134
rect 64794 174454 65414 209898
rect 64794 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 65414 174454
rect 64794 174134 65414 174218
rect 64794 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 65414 174134
rect 64794 138454 65414 173898
rect 64794 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 65414 138454
rect 64794 138134 65414 138218
rect 64794 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 65414 138134
rect 64794 102454 65414 137898
rect 64794 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 65414 102454
rect 64794 102134 65414 102218
rect 64794 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 65414 102134
rect 64794 66454 65414 101898
rect 64794 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 65414 66454
rect 64794 66134 65414 66218
rect 64794 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 65414 66134
rect 64794 30454 65414 65898
rect 64794 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 65414 30454
rect 64794 30134 65414 30218
rect 64794 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 65414 30134
rect 64794 -6106 65414 29898
rect 64794 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 65414 -6106
rect 64794 -6426 65414 -6342
rect 64794 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 65414 -6426
rect 64794 -7654 65414 -6662
rect 69294 214954 69914 228484
rect 69294 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 69914 214954
rect 69294 214634 69914 214718
rect 69294 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 69914 214634
rect 69294 178954 69914 214398
rect 69294 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 69914 178954
rect 69294 178634 69914 178718
rect 69294 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 69914 178634
rect 69294 142954 69914 178398
rect 69294 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 69914 142954
rect 69294 142634 69914 142718
rect 69294 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 69914 142634
rect 69294 106954 69914 142398
rect 69294 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 69914 106954
rect 69294 106634 69914 106718
rect 69294 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 69914 106634
rect 69294 70954 69914 106398
rect 69294 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 69914 70954
rect 69294 70634 69914 70718
rect 69294 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 69914 70634
rect 69294 34954 69914 70398
rect 69294 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 69914 34954
rect 69294 34634 69914 34718
rect 69294 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 69914 34634
rect 69294 -7066 69914 34398
rect 69294 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 69914 -7066
rect 69294 -7386 69914 -7302
rect 69294 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 69914 -7386
rect 69294 -7654 69914 -7622
rect 73794 219454 74414 228484
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 78294 223954 78914 228484
rect 78294 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 78914 223954
rect 78294 223634 78914 223718
rect 78294 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 78914 223634
rect 78294 187954 78914 223398
rect 78294 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 78914 187954
rect 78294 187634 78914 187718
rect 78294 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 78914 187634
rect 78294 151954 78914 187398
rect 78294 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 78914 151954
rect 78294 151634 78914 151718
rect 78294 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 78914 151634
rect 78294 115954 78914 151398
rect 78294 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 78914 115954
rect 78294 115634 78914 115718
rect 78294 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 78914 115634
rect 78294 79954 78914 115398
rect 78294 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 78914 79954
rect 78294 79634 78914 79718
rect 78294 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 78914 79634
rect 78294 43954 78914 79398
rect 78294 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 78914 43954
rect 78294 43634 78914 43718
rect 78294 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 78914 43634
rect 78294 7954 78914 43398
rect 78294 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 78914 7954
rect 78294 7634 78914 7718
rect 78294 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 78914 7634
rect 78294 -1306 78914 7398
rect 78294 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 78914 -1306
rect 78294 -1626 78914 -1542
rect 78294 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 78914 -1626
rect 78294 -7654 78914 -1862
rect 82794 228453 83414 228484
rect 82794 228217 82826 228453
rect 83062 228217 83146 228453
rect 83382 228217 83414 228453
rect 82794 228133 83414 228217
rect 82794 227897 82826 228133
rect 83062 227897 83146 228133
rect 83382 227897 83414 228133
rect 82794 192454 83414 227897
rect 82794 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 83414 192454
rect 82794 192134 83414 192218
rect 82794 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 83414 192134
rect 82794 156454 83414 191898
rect 82794 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 83414 156454
rect 82794 156134 83414 156218
rect 82794 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 83414 156134
rect 82794 120454 83414 155898
rect 82794 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 83414 120454
rect 82794 120134 83414 120218
rect 82794 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 83414 120134
rect 82794 84454 83414 119898
rect 82794 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 83414 84454
rect 82794 84134 83414 84218
rect 82794 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 83414 84134
rect 82794 48454 83414 83898
rect 82794 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 83414 48454
rect 82794 48134 83414 48218
rect 82794 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 83414 48134
rect 82794 12454 83414 47898
rect 82794 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 83414 12454
rect 82794 12134 83414 12218
rect 82794 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 83414 12134
rect 82794 -2266 83414 11898
rect 82794 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 83414 -2266
rect 82794 -2586 83414 -2502
rect 82794 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 83414 -2586
rect 82794 -7654 83414 -2822
rect 87294 196954 87914 228484
rect 87294 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 87914 196954
rect 87294 196634 87914 196718
rect 87294 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 87914 196634
rect 87294 160954 87914 196398
rect 87294 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 87914 160954
rect 87294 160634 87914 160718
rect 87294 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 87914 160634
rect 87294 124954 87914 160398
rect 87294 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 87914 124954
rect 87294 124634 87914 124718
rect 87294 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 87914 124634
rect 87294 88954 87914 124398
rect 87294 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 87914 88954
rect 87294 88634 87914 88718
rect 87294 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 87914 88634
rect 87294 52954 87914 88398
rect 87294 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 87914 52954
rect 87294 52634 87914 52718
rect 87294 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 87914 52634
rect 87294 16954 87914 52398
rect 87294 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 87914 16954
rect 87294 16634 87914 16718
rect 87294 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 87914 16634
rect 87294 -3226 87914 16398
rect 87294 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 87914 -3226
rect 87294 -3546 87914 -3462
rect 87294 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 87914 -3546
rect 87294 -7654 87914 -3782
rect 91794 201454 92414 228484
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 129454 92414 164898
rect 91794 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 92414 129454
rect 91794 129134 92414 129218
rect 91794 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 92414 129134
rect 91794 93454 92414 128898
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 91794 57454 92414 92898
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -4186 92414 20898
rect 91794 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 92414 -4186
rect 91794 -4506 92414 -4422
rect 91794 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 92414 -4506
rect 91794 -7654 92414 -4742
rect 96294 205954 96914 228484
rect 96294 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 96914 205954
rect 96294 205634 96914 205718
rect 96294 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 96914 205634
rect 96294 169954 96914 205398
rect 96294 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 96914 169954
rect 96294 169634 96914 169718
rect 96294 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 96914 169634
rect 96294 133954 96914 169398
rect 96294 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 96914 133954
rect 96294 133634 96914 133718
rect 96294 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 96914 133634
rect 96294 97954 96914 133398
rect 96294 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 96914 97954
rect 96294 97634 96914 97718
rect 96294 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 96914 97634
rect 96294 61954 96914 97398
rect 96294 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 96914 61954
rect 96294 61634 96914 61718
rect 96294 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 96914 61634
rect 96294 25954 96914 61398
rect 96294 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 96914 25954
rect 96294 25634 96914 25718
rect 96294 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 96914 25634
rect 96294 -5146 96914 25398
rect 96294 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 96914 -5146
rect 96294 -5466 96914 -5382
rect 96294 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 96914 -5466
rect 96294 -7654 96914 -5702
rect 100794 210454 101414 228484
rect 100794 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 101414 210454
rect 100794 210134 101414 210218
rect 100794 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 101414 210134
rect 100794 174454 101414 209898
rect 100794 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 101414 174454
rect 100794 174134 101414 174218
rect 100794 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 101414 174134
rect 100794 138454 101414 173898
rect 100794 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 101414 138454
rect 100794 138134 101414 138218
rect 100794 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 101414 138134
rect 100794 102454 101414 137898
rect 100794 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 101414 102454
rect 100794 102134 101414 102218
rect 100794 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 101414 102134
rect 100794 66454 101414 101898
rect 100794 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 101414 66454
rect 100794 66134 101414 66218
rect 100794 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 101414 66134
rect 100794 30454 101414 65898
rect 100794 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 101414 30454
rect 100794 30134 101414 30218
rect 100794 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 101414 30134
rect 100794 -6106 101414 29898
rect 100794 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 101414 -6106
rect 100794 -6426 101414 -6342
rect 100794 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 101414 -6426
rect 100794 -7654 101414 -6662
rect 105294 214954 105914 228484
rect 105294 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 105914 214954
rect 105294 214634 105914 214718
rect 105294 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 105914 214634
rect 105294 178954 105914 214398
rect 105294 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 105914 178954
rect 105294 178634 105914 178718
rect 105294 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 105914 178634
rect 105294 142954 105914 178398
rect 105294 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 105914 142954
rect 105294 142634 105914 142718
rect 105294 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 105914 142634
rect 105294 106954 105914 142398
rect 105294 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 105914 106954
rect 105294 106634 105914 106718
rect 105294 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 105914 106634
rect 105294 70954 105914 106398
rect 105294 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 105914 70954
rect 105294 70634 105914 70718
rect 105294 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 105914 70634
rect 105294 34954 105914 70398
rect 105294 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 105914 34954
rect 105294 34634 105914 34718
rect 105294 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 105914 34634
rect 105294 -7066 105914 34398
rect 105294 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 105914 -7066
rect 105294 -7386 105914 -7302
rect 105294 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 105914 -7386
rect 105294 -7654 105914 -7622
rect 109794 219454 110414 228484
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 114294 223954 114914 228484
rect 114294 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 114914 223954
rect 114294 223634 114914 223718
rect 114294 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 114914 223634
rect 114294 187954 114914 223398
rect 114294 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 114914 187954
rect 114294 187634 114914 187718
rect 114294 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 114914 187634
rect 114294 151954 114914 187398
rect 114294 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 114914 151954
rect 114294 151634 114914 151718
rect 114294 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 114914 151634
rect 114294 137000 114914 151398
rect 118794 228453 119414 228484
rect 118794 228217 118826 228453
rect 119062 228217 119146 228453
rect 119382 228217 119414 228453
rect 118794 228133 119414 228217
rect 118794 227897 118826 228133
rect 119062 227897 119146 228133
rect 119382 227897 119414 228133
rect 118794 192454 119414 227897
rect 118794 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 119414 192454
rect 118794 192134 119414 192218
rect 118794 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 119414 192134
rect 118794 156454 119414 191898
rect 118794 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 119414 156454
rect 118794 156134 119414 156218
rect 118794 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 119414 156134
rect 118794 137000 119414 155898
rect 123294 196954 123914 228484
rect 123294 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 123914 196954
rect 123294 196634 123914 196718
rect 123294 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 123914 196634
rect 123294 160954 123914 196398
rect 123294 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 123914 160954
rect 123294 160634 123914 160718
rect 123294 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 123914 160634
rect 123294 137000 123914 160398
rect 127794 201454 128414 228484
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 127794 165454 128414 200898
rect 127794 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 128414 165454
rect 127794 165134 128414 165218
rect 127794 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 128414 165134
rect 127794 137000 128414 164898
rect 132294 205954 132914 228484
rect 172794 210454 173414 228484
rect 172794 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 173414 210454
rect 172794 210134 173414 210218
rect 172794 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 173414 210134
rect 132294 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205718 132914 205954
rect 132294 205634 132914 205718
rect 132294 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205398 132914 205634
rect 135914 205861 165514 205986
rect 135914 205625 136036 205861
rect 136272 205625 136356 205861
rect 136592 205625 136676 205861
rect 136912 205625 136996 205861
rect 137232 205625 137316 205861
rect 137552 205625 137636 205861
rect 137872 205625 137956 205861
rect 138192 205625 138276 205861
rect 138512 205625 138596 205861
rect 138832 205625 138916 205861
rect 139152 205625 139236 205861
rect 139472 205625 139556 205861
rect 139792 205625 139876 205861
rect 140112 205625 140196 205861
rect 140432 205625 140516 205861
rect 140752 205625 140836 205861
rect 141072 205625 141156 205861
rect 141392 205625 141476 205861
rect 141712 205625 141796 205861
rect 142032 205625 142116 205861
rect 142352 205625 142436 205861
rect 142672 205625 142756 205861
rect 142992 205625 143076 205861
rect 143312 205625 143396 205861
rect 143632 205625 143716 205861
rect 143952 205625 144036 205861
rect 144272 205625 144356 205861
rect 144592 205625 144676 205861
rect 144912 205625 144996 205861
rect 145232 205625 145316 205861
rect 145552 205625 145636 205861
rect 145872 205625 145956 205861
rect 146192 205625 146276 205861
rect 146512 205625 146596 205861
rect 146832 205625 146916 205861
rect 147152 205625 147236 205861
rect 147472 205625 147556 205861
rect 147792 205625 147876 205861
rect 148112 205625 148196 205861
rect 148432 205625 148516 205861
rect 148752 205625 148836 205861
rect 149072 205625 149156 205861
rect 149392 205625 149476 205861
rect 149712 205625 149796 205861
rect 150032 205625 150116 205861
rect 150352 205625 150436 205861
rect 150672 205625 150756 205861
rect 150992 205625 151076 205861
rect 151312 205625 151396 205861
rect 151632 205625 151716 205861
rect 151952 205625 152036 205861
rect 152272 205625 152356 205861
rect 152592 205625 152676 205861
rect 152912 205625 152996 205861
rect 153232 205625 153316 205861
rect 153552 205625 153636 205861
rect 153872 205625 153956 205861
rect 154192 205625 154276 205861
rect 154512 205625 154596 205861
rect 154832 205625 154916 205861
rect 155152 205625 155236 205861
rect 155472 205625 155556 205861
rect 155792 205625 155876 205861
rect 156112 205625 156196 205861
rect 156432 205625 156516 205861
rect 156752 205625 156836 205861
rect 157072 205625 157156 205861
rect 157392 205625 157476 205861
rect 157712 205625 157796 205861
rect 158032 205625 158116 205861
rect 158352 205625 158436 205861
rect 158672 205625 158756 205861
rect 158992 205625 159076 205861
rect 159312 205625 159396 205861
rect 159632 205625 159716 205861
rect 159952 205625 160036 205861
rect 160272 205625 160356 205861
rect 160592 205625 160676 205861
rect 160912 205625 160996 205861
rect 161232 205625 161316 205861
rect 161552 205625 161636 205861
rect 161872 205625 161956 205861
rect 162192 205625 162276 205861
rect 162512 205625 162596 205861
rect 162832 205625 162916 205861
rect 163152 205625 163236 205861
rect 163472 205625 163556 205861
rect 163792 205625 163876 205861
rect 164112 205625 164196 205861
rect 164432 205625 164516 205861
rect 164752 205625 164836 205861
rect 165072 205625 165156 205861
rect 165392 205625 165514 205861
rect 135914 205500 165514 205625
rect 132294 169954 132914 205398
rect 137314 201411 165514 201486
rect 137314 201175 137376 201411
rect 137612 201175 137696 201411
rect 137932 201175 138016 201411
rect 138252 201175 138336 201411
rect 138572 201175 138656 201411
rect 138892 201175 138976 201411
rect 139212 201175 139296 201411
rect 139532 201175 139616 201411
rect 139852 201175 139936 201411
rect 140172 201175 140256 201411
rect 140492 201175 140576 201411
rect 140812 201175 140896 201411
rect 141132 201175 141216 201411
rect 141452 201175 141536 201411
rect 141772 201175 141856 201411
rect 142092 201175 142176 201411
rect 142412 201175 142496 201411
rect 142732 201175 142816 201411
rect 143052 201175 143136 201411
rect 143372 201175 143456 201411
rect 143692 201175 143776 201411
rect 144012 201175 144096 201411
rect 144332 201175 144416 201411
rect 144652 201175 144736 201411
rect 144972 201175 145056 201411
rect 145292 201175 145376 201411
rect 145612 201175 145696 201411
rect 145932 201175 146016 201411
rect 146252 201175 146336 201411
rect 146572 201175 146656 201411
rect 146892 201175 146976 201411
rect 147212 201175 147296 201411
rect 147532 201175 147616 201411
rect 147852 201175 147936 201411
rect 148172 201175 148256 201411
rect 148492 201175 148576 201411
rect 148812 201175 148896 201411
rect 149132 201175 149216 201411
rect 149452 201175 149536 201411
rect 149772 201175 149856 201411
rect 150092 201175 150176 201411
rect 150412 201175 150496 201411
rect 150732 201175 150816 201411
rect 151052 201175 151136 201411
rect 151372 201175 151456 201411
rect 151692 201175 151776 201411
rect 152012 201175 152096 201411
rect 152332 201175 152416 201411
rect 152652 201175 152736 201411
rect 152972 201175 153056 201411
rect 153292 201175 153376 201411
rect 153612 201175 153696 201411
rect 153932 201175 154016 201411
rect 154252 201175 154336 201411
rect 154572 201175 154656 201411
rect 154892 201175 154976 201411
rect 155212 201175 155296 201411
rect 155532 201175 155616 201411
rect 155852 201175 155936 201411
rect 156172 201175 156256 201411
rect 156492 201175 156576 201411
rect 156812 201175 156896 201411
rect 157132 201175 157216 201411
rect 157452 201175 157536 201411
rect 157772 201175 157856 201411
rect 158092 201175 158176 201411
rect 158412 201175 158496 201411
rect 158732 201175 158816 201411
rect 159052 201175 159136 201411
rect 159372 201175 159456 201411
rect 159692 201175 159776 201411
rect 160012 201175 160096 201411
rect 160332 201175 160416 201411
rect 160652 201175 160736 201411
rect 160972 201175 161056 201411
rect 161292 201175 161376 201411
rect 161612 201175 161696 201411
rect 161932 201175 162016 201411
rect 162252 201175 162336 201411
rect 162572 201175 162656 201411
rect 162892 201175 162976 201411
rect 163212 201175 163296 201411
rect 163532 201175 163616 201411
rect 163852 201175 163936 201411
rect 164172 201175 164256 201411
rect 164492 201175 164576 201411
rect 164812 201175 164896 201411
rect 165132 201175 165216 201411
rect 165452 201175 165514 201411
rect 137314 201100 165514 201175
rect 143395 193356 143461 193357
rect 143395 193292 143396 193356
rect 143460 193292 143461 193356
rect 143395 193291 143461 193292
rect 155171 193356 155237 193357
rect 155171 193292 155172 193356
rect 155236 193292 155237 193356
rect 155171 193291 155237 193292
rect 141187 184380 141253 184381
rect 141187 184316 141188 184380
rect 141252 184316 141253 184380
rect 141187 184315 141253 184316
rect 140819 184244 140885 184245
rect 140819 184180 140820 184244
rect 140884 184180 140885 184244
rect 140819 184179 140885 184180
rect 140822 178669 140882 184179
rect 141190 178805 141250 184315
rect 142843 184108 142909 184109
rect 142843 184044 142844 184108
rect 142908 184044 142909 184108
rect 142843 184043 142909 184044
rect 142291 179076 142357 179077
rect 142291 179012 142292 179076
rect 142356 179012 142357 179076
rect 142291 179011 142357 179012
rect 141187 178804 141253 178805
rect 141187 178740 141188 178804
rect 141252 178740 141253 178804
rect 141187 178739 141253 178740
rect 140819 178668 140885 178669
rect 140819 178604 140820 178668
rect 140884 178604 140885 178668
rect 140819 178603 140885 178604
rect 142294 176670 142354 179011
rect 142846 178941 142906 184043
rect 143398 181253 143458 193291
rect 143579 191632 143645 191633
rect 143579 191568 143580 191632
rect 143644 191568 143645 191632
rect 143579 191567 143645 191568
rect 143395 181252 143461 181253
rect 143395 181188 143396 181252
rect 143460 181188 143461 181252
rect 143395 181187 143461 181188
rect 143395 180980 143461 180981
rect 143395 180916 143396 180980
rect 143460 180916 143461 180980
rect 143395 180915 143461 180916
rect 142843 178940 142909 178941
rect 142843 178876 142844 178940
rect 142908 178876 142909 178940
rect 142843 178875 142909 178876
rect 141926 176610 142354 176670
rect 137014 174454 141514 174486
rect 137014 174218 137066 174454
rect 137302 174218 137386 174454
rect 137622 174218 137706 174454
rect 137942 174218 138026 174454
rect 138262 174218 138346 174454
rect 138582 174218 138666 174454
rect 138902 174218 138986 174454
rect 139222 174218 139306 174454
rect 139542 174218 139626 174454
rect 139862 174218 139946 174454
rect 140182 174218 140266 174454
rect 140502 174218 140586 174454
rect 140822 174218 140906 174454
rect 141142 174218 141226 174454
rect 141462 174218 141514 174454
rect 137014 174134 141514 174218
rect 137014 173898 137066 174134
rect 137302 173898 137386 174134
rect 137622 173898 137706 174134
rect 137942 173898 138026 174134
rect 138262 173898 138346 174134
rect 138582 173898 138666 174134
rect 138902 173898 138986 174134
rect 139222 173898 139306 174134
rect 139542 173898 139626 174134
rect 139862 173898 139946 174134
rect 140182 173898 140266 174134
rect 140502 173898 140586 174134
rect 140822 173898 140906 174134
rect 141142 173898 141226 174134
rect 141462 173898 141514 174134
rect 137014 173866 141514 173898
rect 132294 169718 132326 169954
rect 132562 169718 132646 169954
rect 132882 169718 132914 169954
rect 132294 169634 132914 169718
rect 132294 169398 132326 169634
rect 132562 169398 132646 169634
rect 132882 169398 132914 169634
rect 132294 137000 132914 169398
rect 141926 138005 141986 176610
rect 141923 138004 141989 138005
rect 141923 137940 141924 138004
rect 141988 137940 141989 138004
rect 141923 137939 141989 137940
rect 143398 137461 143458 180915
rect 143582 137733 143642 191567
rect 144499 191044 144565 191045
rect 144499 190980 144500 191044
rect 144564 190980 144565 191044
rect 144499 190979 144565 190980
rect 144502 189277 144562 190979
rect 145787 189820 145853 189821
rect 145787 189756 145788 189820
rect 145852 189756 145853 189820
rect 145787 189755 145853 189756
rect 144499 189276 144565 189277
rect 144499 189212 144500 189276
rect 144564 189212 144565 189276
rect 144499 189211 144565 189212
rect 145790 179430 145850 189755
rect 155174 189005 155234 193291
rect 155171 189004 155237 189005
rect 155171 188940 155172 189004
rect 155236 188940 155237 189004
rect 155171 188939 155237 188940
rect 147259 182068 147325 182069
rect 147259 182004 147260 182068
rect 147324 182004 147325 182068
rect 147259 182003 147325 182004
rect 145790 179370 146218 179430
rect 143579 137732 143645 137733
rect 143579 137668 143580 137732
rect 143644 137668 143645 137732
rect 143579 137667 143645 137668
rect 146158 137597 146218 179370
rect 147262 174589 147322 182003
rect 147259 174588 147325 174589
rect 147259 174524 147260 174588
rect 147324 174524 147325 174588
rect 147259 174523 147325 174524
rect 172794 174454 173414 209898
rect 172794 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 173414 174454
rect 172794 174134 173414 174218
rect 172794 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 173414 174134
rect 172794 138454 173414 173898
rect 172794 138218 172826 138454
rect 173062 138218 173146 138454
rect 173382 138218 173414 138454
rect 172794 138134 173414 138218
rect 172794 137898 172826 138134
rect 173062 137898 173146 138134
rect 173382 137898 173414 138134
rect 146155 137596 146221 137597
rect 146155 137532 146156 137596
rect 146220 137532 146221 137596
rect 146155 137531 146221 137532
rect 143395 137460 143461 137461
rect 143395 137396 143396 137460
rect 143460 137396 143461 137460
rect 143395 137395 143461 137396
rect 172794 137000 173414 137898
rect 177294 214954 177914 228484
rect 177294 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 177914 214954
rect 177294 214634 177914 214718
rect 177294 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 177914 214634
rect 177294 178954 177914 214398
rect 177294 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 177914 178954
rect 177294 178634 177914 178718
rect 177294 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 177914 178634
rect 177294 142954 177914 178398
rect 177294 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 177914 142954
rect 177294 142634 177914 142718
rect 177294 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 177914 142634
rect 177294 137000 177914 142398
rect 181794 219454 182414 228484
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 135568 115954 135888 115986
rect 135568 115718 135610 115954
rect 135846 115718 135888 115954
rect 135568 115634 135888 115718
rect 135568 115398 135610 115634
rect 135846 115398 135888 115634
rect 135568 115366 135888 115398
rect 166288 115954 166608 115986
rect 166288 115718 166330 115954
rect 166566 115718 166608 115954
rect 166288 115634 166608 115718
rect 166288 115398 166330 115634
rect 166566 115398 166608 115634
rect 166288 115366 166608 115398
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 120208 111454 120528 111486
rect 120208 111218 120250 111454
rect 120486 111218 120528 111454
rect 120208 111134 120528 111218
rect 120208 110898 120250 111134
rect 120486 110898 120528 111134
rect 120208 110866 120528 110898
rect 150928 111454 151248 111486
rect 150928 111218 150970 111454
rect 151206 111218 151248 111454
rect 150928 111134 151248 111218
rect 150928 110898 150970 111134
rect 151206 110898 151248 111134
rect 150928 110866 151248 110898
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 135568 79954 135888 79986
rect 135568 79718 135610 79954
rect 135846 79718 135888 79954
rect 135568 79634 135888 79718
rect 135568 79398 135610 79634
rect 135846 79398 135888 79634
rect 135568 79366 135888 79398
rect 166288 79954 166608 79986
rect 166288 79718 166330 79954
rect 166566 79718 166608 79954
rect 166288 79634 166608 79718
rect 166288 79398 166330 79634
rect 166566 79398 166608 79634
rect 166288 79366 166608 79398
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 168606 75790 169402 75850
rect 168419 75444 168485 75445
rect 168419 75380 168420 75444
rect 168484 75380 168485 75444
rect 168419 75379 168485 75380
rect 167683 75308 167749 75309
rect 167683 75244 167684 75308
rect 167748 75244 167749 75308
rect 167683 75243 167749 75244
rect 109794 75134 110414 75218
rect 167686 75170 167746 75243
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 167502 75110 167746 75170
rect 109794 39454 110414 74898
rect 162899 74900 162965 74901
rect 162899 74836 162900 74900
rect 162964 74836 162965 74900
rect 162899 74835 162965 74836
rect 128491 73132 128557 73133
rect 128491 73068 128492 73132
rect 128556 73068 128557 73132
rect 128491 73067 128557 73068
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 114294 43954 114914 73000
rect 114294 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 114914 43954
rect 114294 43634 114914 43718
rect 114294 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 114914 43634
rect 114294 7954 114914 43398
rect 114294 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 114914 7954
rect 114294 7634 114914 7718
rect 114294 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 114914 7634
rect 114294 -1306 114914 7398
rect 114294 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 114914 -1306
rect 114294 -1626 114914 -1542
rect 114294 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 114914 -1626
rect 114294 -7654 114914 -1862
rect 118794 48454 119414 73000
rect 121683 72044 121749 72045
rect 121683 71980 121684 72044
rect 121748 71980 121749 72044
rect 121683 71979 121749 71980
rect 122787 72044 122853 72045
rect 122787 71980 122788 72044
rect 122852 71980 122853 72044
rect 122787 71979 122853 71980
rect 121499 71908 121565 71909
rect 121499 71844 121500 71908
rect 121564 71844 121565 71908
rect 121499 71843 121565 71844
rect 118794 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 119414 48454
rect 118794 48134 119414 48218
rect 118794 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 119414 48134
rect 118794 12454 119414 47898
rect 118794 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 119414 12454
rect 118794 12134 119414 12218
rect 118794 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 119414 12134
rect 118794 -2266 119414 11898
rect 121502 3365 121562 71843
rect 121686 3501 121746 71979
rect 122790 71770 122850 71979
rect 122971 71908 123037 71909
rect 122971 71844 122972 71908
rect 123036 71844 123037 71908
rect 122971 71843 123037 71844
rect 122606 71710 122850 71770
rect 122606 3637 122666 71710
rect 122974 6221 123034 71843
rect 123294 52954 123914 73000
rect 126099 72316 126165 72317
rect 126099 72252 126100 72316
rect 126164 72252 126165 72316
rect 126099 72251 126165 72252
rect 124627 72180 124693 72181
rect 124627 72116 124628 72180
rect 124692 72116 124693 72180
rect 124627 72115 124693 72116
rect 125547 72180 125613 72181
rect 125547 72116 125548 72180
rect 125612 72116 125613 72180
rect 125547 72115 125613 72116
rect 124259 72044 124325 72045
rect 124259 71980 124260 72044
rect 124324 71980 124325 72044
rect 124259 71979 124325 71980
rect 123294 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 123914 52954
rect 123294 52634 123914 52718
rect 123294 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 123914 52634
rect 123294 16954 123914 52398
rect 123294 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 123914 16954
rect 123294 16634 123914 16718
rect 123294 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 123914 16634
rect 122971 6220 123037 6221
rect 122971 6156 122972 6220
rect 123036 6156 123037 6220
rect 122971 6155 123037 6156
rect 122603 3636 122669 3637
rect 122603 3572 122604 3636
rect 122668 3572 122669 3636
rect 122603 3571 122669 3572
rect 121683 3500 121749 3501
rect 121683 3436 121684 3500
rect 121748 3436 121749 3500
rect 121683 3435 121749 3436
rect 121499 3364 121565 3365
rect 121499 3300 121500 3364
rect 121564 3300 121565 3364
rect 121499 3299 121565 3300
rect 118794 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 119414 -2266
rect 118794 -2586 119414 -2502
rect 118794 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 119414 -2586
rect 118794 -7654 119414 -2822
rect 123294 -3226 123914 16398
rect 124262 4861 124322 71979
rect 124443 71908 124509 71909
rect 124443 71844 124444 71908
rect 124508 71844 124509 71908
rect 124443 71843 124509 71844
rect 124446 9077 124506 71843
rect 124443 9076 124509 9077
rect 124443 9012 124444 9076
rect 124508 9012 124509 9076
rect 124443 9011 124509 9012
rect 124630 8941 124690 72115
rect 124627 8940 124693 8941
rect 124627 8876 124628 8940
rect 124692 8876 124693 8940
rect 124627 8875 124693 8876
rect 124259 4860 124325 4861
rect 124259 4796 124260 4860
rect 124324 4796 124325 4860
rect 124259 4795 124325 4796
rect 125550 3773 125610 72115
rect 125731 72044 125797 72045
rect 125731 71980 125732 72044
rect 125796 71980 125797 72044
rect 125731 71979 125797 71980
rect 125734 6357 125794 71979
rect 125915 71908 125981 71909
rect 125915 71844 125916 71908
rect 125980 71844 125981 71908
rect 125915 71843 125981 71844
rect 125918 6493 125978 71843
rect 126102 9213 126162 72251
rect 127203 72044 127269 72045
rect 127203 71980 127204 72044
rect 127268 71980 127269 72044
rect 127203 71979 127269 71980
rect 127019 71908 127085 71909
rect 127019 71844 127020 71908
rect 127084 71844 127085 71908
rect 127019 71843 127085 71844
rect 126099 9212 126165 9213
rect 126099 9148 126100 9212
rect 126164 9148 126165 9212
rect 126099 9147 126165 9148
rect 127022 7581 127082 71843
rect 127206 10301 127266 71979
rect 127794 57454 128414 73000
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127203 10300 127269 10301
rect 127203 10236 127204 10300
rect 127268 10236 127269 10300
rect 127203 10235 127269 10236
rect 127019 7580 127085 7581
rect 127019 7516 127020 7580
rect 127084 7516 127085 7580
rect 127019 7515 127085 7516
rect 125915 6492 125981 6493
rect 125915 6428 125916 6492
rect 125980 6428 125981 6492
rect 125915 6427 125981 6428
rect 125731 6356 125797 6357
rect 125731 6292 125732 6356
rect 125796 6292 125797 6356
rect 125731 6291 125797 6292
rect 125547 3772 125613 3773
rect 125547 3708 125548 3772
rect 125612 3708 125613 3772
rect 125547 3707 125613 3708
rect 123294 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 123914 -3226
rect 123294 -3546 123914 -3462
rect 123294 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 123914 -3546
rect 123294 -7654 123914 -3782
rect 127794 -4186 128414 20898
rect 128494 6930 128554 73067
rect 129043 72180 129109 72181
rect 129043 72116 129044 72180
rect 129108 72116 129109 72180
rect 129043 72115 129109 72116
rect 129963 72180 130029 72181
rect 129963 72116 129964 72180
rect 130028 72116 130029 72180
rect 129963 72115 130029 72116
rect 128859 72044 128925 72045
rect 128859 71980 128860 72044
rect 128924 71980 128925 72044
rect 128859 71979 128925 71980
rect 128675 71908 128741 71909
rect 128675 71844 128676 71908
rect 128740 71844 128741 71908
rect 128675 71843 128741 71844
rect 128678 7853 128738 71843
rect 128675 7852 128741 7853
rect 128675 7788 128676 7852
rect 128740 7788 128741 7852
rect 128675 7787 128741 7788
rect 128862 7717 128922 71979
rect 129046 10437 129106 72115
rect 129779 71908 129845 71909
rect 129779 71844 129780 71908
rect 129844 71844 129845 71908
rect 129779 71843 129845 71844
rect 129043 10436 129109 10437
rect 129043 10372 129044 10436
rect 129108 10372 129109 10436
rect 129043 10371 129109 10372
rect 128859 7716 128925 7717
rect 128859 7652 128860 7716
rect 128924 7652 128925 7716
rect 128859 7651 128925 7652
rect 128494 6870 128738 6930
rect 128678 4997 128738 6870
rect 129782 6629 129842 71843
rect 129966 9349 130026 72115
rect 130147 72044 130213 72045
rect 130147 71980 130148 72044
rect 130212 71980 130213 72044
rect 130147 71979 130213 71980
rect 131251 72044 131317 72045
rect 131251 71980 131252 72044
rect 131316 71980 131317 72044
rect 131251 71979 131317 71980
rect 131803 72044 131869 72045
rect 131803 71980 131804 72044
rect 131868 71980 131869 72044
rect 131803 71979 131869 71980
rect 130150 9485 130210 71979
rect 131067 71908 131133 71909
rect 131067 71844 131068 71908
rect 131132 71844 131133 71908
rect 131067 71843 131133 71844
rect 130147 9484 130213 9485
rect 130147 9420 130148 9484
rect 130212 9420 130213 9484
rect 130147 9419 130213 9420
rect 129963 9348 130029 9349
rect 129963 9284 129964 9348
rect 130028 9284 130029 9348
rect 129963 9283 130029 9284
rect 129779 6628 129845 6629
rect 129779 6564 129780 6628
rect 129844 6564 129845 6628
rect 129779 6563 129845 6564
rect 128675 4996 128741 4997
rect 128675 4932 128676 4996
rect 128740 4932 128741 4996
rect 128675 4931 128741 4932
rect 131070 3637 131130 71843
rect 131067 3636 131133 3637
rect 131067 3572 131068 3636
rect 131132 3572 131133 3636
rect 131067 3571 131133 3572
rect 131254 3501 131314 71979
rect 131806 3637 131866 71979
rect 131987 71908 132053 71909
rect 131987 71844 131988 71908
rect 132052 71844 132053 71908
rect 131987 71843 132053 71844
rect 131803 3636 131869 3637
rect 131803 3572 131804 3636
rect 131868 3572 131869 3636
rect 131803 3571 131869 3572
rect 131990 3501 132050 71843
rect 132294 61954 132914 73000
rect 133275 72180 133341 72181
rect 133275 72116 133276 72180
rect 133340 72116 133341 72180
rect 133275 72115 133341 72116
rect 134747 72180 134813 72181
rect 134747 72116 134748 72180
rect 134812 72116 134813 72180
rect 134747 72115 134813 72116
rect 136035 72180 136101 72181
rect 136035 72116 136036 72180
rect 136100 72116 136101 72180
rect 136035 72115 136101 72116
rect 132294 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 132914 61954
rect 132294 61634 132914 61718
rect 132294 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 132914 61634
rect 132294 25954 132914 61398
rect 132294 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 132914 25954
rect 132294 25634 132914 25718
rect 132294 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 132914 25634
rect 131251 3500 131317 3501
rect 131251 3436 131252 3500
rect 131316 3436 131317 3500
rect 131251 3435 131317 3436
rect 131987 3500 132053 3501
rect 131987 3436 131988 3500
rect 132052 3436 132053 3500
rect 131987 3435 132053 3436
rect 127794 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 128414 -4186
rect 127794 -4506 128414 -4422
rect 127794 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 128414 -4506
rect 127794 -7654 128414 -4742
rect 132294 -5146 132914 25398
rect 133278 4997 133338 72115
rect 133459 72044 133525 72045
rect 133459 71980 133460 72044
rect 133524 71980 133525 72044
rect 133459 71979 133525 71980
rect 133275 4996 133341 4997
rect 133275 4932 133276 4996
rect 133340 4932 133341 4996
rect 133275 4931 133341 4932
rect 133462 4861 133522 71979
rect 133643 71908 133709 71909
rect 133643 71844 133644 71908
rect 133708 71844 133709 71908
rect 133643 71843 133709 71844
rect 133459 4860 133525 4861
rect 133459 4796 133460 4860
rect 133524 4796 133525 4860
rect 133459 4795 133525 4796
rect 133646 3365 133706 71843
rect 134750 32741 134810 72115
rect 134931 72044 134997 72045
rect 134931 71980 134932 72044
rect 134996 71980 134997 72044
rect 134931 71979 134997 71980
rect 134747 32740 134813 32741
rect 134747 32676 134748 32740
rect 134812 32676 134813 32740
rect 134747 32675 134813 32676
rect 134934 25669 134994 71979
rect 135115 71908 135181 71909
rect 135115 71844 135116 71908
rect 135180 71844 135181 71908
rect 135115 71843 135181 71844
rect 135851 71908 135917 71909
rect 135851 71844 135852 71908
rect 135916 71844 135917 71908
rect 135851 71843 135917 71844
rect 134931 25668 134997 25669
rect 134931 25604 134932 25668
rect 134996 25604 134997 25668
rect 134931 25603 134997 25604
rect 135118 8125 135178 71843
rect 135854 32605 135914 71843
rect 135851 32604 135917 32605
rect 135851 32540 135852 32604
rect 135916 32540 135917 32604
rect 135851 32539 135917 32540
rect 136038 32469 136098 72115
rect 136219 72044 136285 72045
rect 136219 71980 136220 72044
rect 136284 71980 136285 72044
rect 136219 71979 136285 71980
rect 136035 32468 136101 32469
rect 136035 32404 136036 32468
rect 136100 32404 136101 32468
rect 136035 32403 136101 32404
rect 136222 27165 136282 71979
rect 136403 71908 136469 71909
rect 136403 71844 136404 71908
rect 136468 71844 136469 71908
rect 136403 71843 136469 71844
rect 136219 27164 136285 27165
rect 136219 27100 136220 27164
rect 136284 27100 136285 27164
rect 136219 27099 136285 27100
rect 135115 8124 135181 8125
rect 135115 8060 135116 8124
rect 135180 8060 135181 8124
rect 135115 8059 135181 8060
rect 136406 4725 136466 71843
rect 136794 66454 137414 73000
rect 138979 72180 139045 72181
rect 138979 72116 138980 72180
rect 139044 72116 139045 72180
rect 138979 72115 139045 72116
rect 140083 72180 140149 72181
rect 140083 72116 140084 72180
rect 140148 72116 140149 72180
rect 140083 72115 140149 72116
rect 137691 72044 137757 72045
rect 137691 71980 137692 72044
rect 137756 71980 137757 72044
rect 137691 71979 137757 71980
rect 138795 72044 138861 72045
rect 138795 71980 138796 72044
rect 138860 71980 138861 72044
rect 138795 71979 138861 71980
rect 136794 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 137414 66454
rect 136794 66134 137414 66218
rect 136794 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 137414 66134
rect 136794 30454 137414 65898
rect 137694 34101 137754 71979
rect 137875 71908 137941 71909
rect 137875 71844 137876 71908
rect 137940 71844 137941 71908
rect 137875 71843 137941 71844
rect 138611 71908 138677 71909
rect 138611 71844 138612 71908
rect 138676 71844 138677 71908
rect 138611 71843 138677 71844
rect 137691 34100 137757 34101
rect 137691 34036 137692 34100
rect 137756 34036 137757 34100
rect 137691 34035 137757 34036
rect 136794 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 137414 30454
rect 136794 30134 137414 30218
rect 136794 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 137414 30134
rect 136403 4724 136469 4725
rect 136403 4660 136404 4724
rect 136468 4660 136469 4724
rect 136403 4659 136469 4660
rect 133643 3364 133709 3365
rect 133643 3300 133644 3364
rect 133708 3300 133709 3364
rect 133643 3299 133709 3300
rect 132294 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 132914 -5146
rect 132294 -5466 132914 -5382
rect 132294 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 132914 -5466
rect 132294 -7654 132914 -5702
rect 136794 -6106 137414 29898
rect 137878 12205 137938 71843
rect 138614 20229 138674 71843
rect 138611 20228 138677 20229
rect 138611 20164 138612 20228
rect 138676 20164 138677 20228
rect 138611 20163 138677 20164
rect 138798 12885 138858 71979
rect 138795 12884 138861 12885
rect 138795 12820 138796 12884
rect 138860 12820 138861 12884
rect 138795 12819 138861 12820
rect 137875 12204 137941 12205
rect 137875 12140 137876 12204
rect 137940 12140 137941 12204
rect 137875 12139 137941 12140
rect 138982 6765 139042 72115
rect 139163 71908 139229 71909
rect 139163 71844 139164 71908
rect 139228 71844 139229 71908
rect 139163 71843 139229 71844
rect 139166 6901 139226 71843
rect 140086 33965 140146 72115
rect 140267 72044 140333 72045
rect 140267 71980 140268 72044
rect 140332 71980 140333 72044
rect 140267 71979 140333 71980
rect 140819 72044 140885 72045
rect 140819 71980 140820 72044
rect 140884 71980 140885 72044
rect 140819 71979 140885 71980
rect 140083 33964 140149 33965
rect 140083 33900 140084 33964
rect 140148 33900 140149 33964
rect 140083 33899 140149 33900
rect 140270 20093 140330 71979
rect 140451 71908 140517 71909
rect 140451 71844 140452 71908
rect 140516 71844 140517 71908
rect 140451 71843 140517 71844
rect 140635 71908 140701 71909
rect 140635 71844 140636 71908
rect 140700 71844 140701 71908
rect 140635 71843 140701 71844
rect 140267 20092 140333 20093
rect 140267 20028 140268 20092
rect 140332 20028 140333 20092
rect 140267 20027 140333 20028
rect 140454 13701 140514 71843
rect 140451 13700 140517 13701
rect 140451 13636 140452 13700
rect 140516 13636 140517 13700
rect 140451 13635 140517 13636
rect 139163 6900 139229 6901
rect 139163 6836 139164 6900
rect 139228 6836 139229 6900
rect 139163 6835 139229 6836
rect 138979 6764 139045 6765
rect 138979 6700 138980 6764
rect 139044 6700 139045 6764
rect 138979 6699 139045 6700
rect 140638 6629 140698 71843
rect 140822 33829 140882 71979
rect 141003 71908 141069 71909
rect 141003 71844 141004 71908
rect 141068 71844 141069 71908
rect 141003 71843 141069 71844
rect 140819 33828 140885 33829
rect 140819 33764 140820 33828
rect 140884 33764 140885 33828
rect 140819 33763 140885 33764
rect 141006 15197 141066 71843
rect 141294 70954 141914 73000
rect 142843 72316 142909 72317
rect 142843 72252 142844 72316
rect 142908 72252 142909 72316
rect 142843 72251 142909 72252
rect 141294 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 141914 70954
rect 141294 70634 141914 70718
rect 141294 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 141914 70634
rect 141294 34954 141914 70398
rect 141294 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 141914 34954
rect 141294 34634 141914 34718
rect 141294 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 141914 34634
rect 141003 15196 141069 15197
rect 141003 15132 141004 15196
rect 141068 15132 141069 15196
rect 141003 15131 141069 15132
rect 140635 6628 140701 6629
rect 140635 6564 140636 6628
rect 140700 6564 140701 6628
rect 140635 6563 140701 6564
rect 136794 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 137414 -6106
rect 136794 -6426 137414 -6342
rect 136794 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 137414 -6426
rect 136794 -7654 137414 -6662
rect 141294 -7066 141914 34398
rect 142846 27029 142906 72251
rect 143027 72180 143093 72181
rect 143027 72116 143028 72180
rect 143092 72116 143093 72180
rect 143027 72115 143093 72116
rect 144131 72180 144197 72181
rect 144131 72116 144132 72180
rect 144196 72116 144197 72180
rect 144131 72115 144197 72116
rect 145235 72180 145301 72181
rect 145235 72116 145236 72180
rect 145300 72116 145301 72180
rect 145235 72115 145301 72116
rect 142843 27028 142909 27029
rect 142843 26964 142844 27028
rect 142908 26964 142909 27028
rect 142843 26963 142909 26964
rect 143030 13565 143090 72115
rect 143211 72044 143277 72045
rect 143211 71980 143212 72044
rect 143276 71980 143277 72044
rect 143211 71979 143277 71980
rect 143027 13564 143093 13565
rect 143027 13500 143028 13564
rect 143092 13500 143093 13564
rect 143027 13499 143093 13500
rect 143214 7853 143274 71979
rect 143395 71908 143461 71909
rect 143395 71844 143396 71908
rect 143460 71844 143461 71908
rect 143395 71843 143461 71844
rect 143398 7989 143458 71843
rect 144134 35325 144194 72115
rect 144499 72044 144565 72045
rect 144499 71980 144500 72044
rect 144564 71980 144565 72044
rect 144499 71979 144565 71980
rect 144315 71908 144381 71909
rect 144315 71844 144316 71908
rect 144380 71844 144381 71908
rect 144315 71843 144381 71844
rect 144131 35324 144197 35325
rect 144131 35260 144132 35324
rect 144196 35260 144197 35324
rect 144131 35259 144197 35260
rect 144318 16285 144378 71843
rect 144315 16284 144381 16285
rect 144315 16220 144316 16284
rect 144380 16220 144381 16284
rect 144315 16219 144381 16220
rect 144502 15061 144562 71979
rect 144683 71908 144749 71909
rect 144683 71844 144684 71908
rect 144748 71844 144749 71908
rect 144683 71843 144749 71844
rect 144499 15060 144565 15061
rect 144499 14996 144500 15060
rect 144564 14996 144565 15060
rect 144499 14995 144565 14996
rect 144686 9213 144746 71843
rect 145238 29613 145298 72115
rect 145419 72044 145485 72045
rect 145419 71980 145420 72044
rect 145484 71980 145485 72044
rect 145419 71979 145485 71980
rect 145235 29612 145301 29613
rect 145235 29548 145236 29612
rect 145300 29548 145301 29612
rect 145235 29547 145301 29548
rect 145422 17645 145482 71979
rect 145603 71908 145669 71909
rect 145603 71844 145604 71908
rect 145668 71844 145669 71908
rect 145603 71843 145669 71844
rect 145419 17644 145485 17645
rect 145419 17580 145420 17644
rect 145484 17580 145485 17644
rect 145419 17579 145485 17580
rect 145606 14925 145666 71843
rect 145794 39454 146414 73000
rect 149467 72996 149533 72997
rect 149467 72932 149468 72996
rect 149532 72932 149533 72996
rect 149467 72931 149533 72932
rect 148731 72860 148797 72861
rect 148731 72796 148732 72860
rect 148796 72796 148797 72860
rect 148731 72795 148797 72796
rect 148363 72588 148429 72589
rect 148363 72524 148364 72588
rect 148428 72524 148429 72588
rect 148363 72523 148429 72524
rect 146891 72180 146957 72181
rect 146891 72116 146892 72180
rect 146956 72116 146957 72180
rect 146891 72115 146957 72116
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145603 14924 145669 14925
rect 145603 14860 145604 14924
rect 145668 14860 145669 14924
rect 145603 14859 145669 14860
rect 144683 9212 144749 9213
rect 144683 9148 144684 9212
rect 144748 9148 144749 9212
rect 144683 9147 144749 9148
rect 143395 7988 143461 7989
rect 143395 7924 143396 7988
rect 143460 7924 143461 7988
rect 143395 7923 143461 7924
rect 143211 7852 143277 7853
rect 143211 7788 143212 7852
rect 143276 7788 143277 7852
rect 143211 7787 143277 7788
rect 141294 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 141914 -7066
rect 141294 -7386 141914 -7302
rect 141294 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 141914 -7386
rect 141294 -7654 141914 -7622
rect 145794 3454 146414 38898
rect 146894 35189 146954 72115
rect 147075 72044 147141 72045
rect 147075 71980 147076 72044
rect 147140 71980 147141 72044
rect 147075 71979 147141 71980
rect 146891 35188 146957 35189
rect 146891 35124 146892 35188
rect 146956 35124 146957 35188
rect 146891 35123 146957 35124
rect 147078 14789 147138 71979
rect 147259 71908 147325 71909
rect 147259 71844 147260 71908
rect 147324 71844 147325 71908
rect 147259 71843 147325 71844
rect 147443 71908 147509 71909
rect 147443 71844 147444 71908
rect 147508 71844 147509 71908
rect 147443 71843 147509 71844
rect 147075 14788 147141 14789
rect 147075 14724 147076 14788
rect 147140 14724 147141 14788
rect 147075 14723 147141 14724
rect 147262 10437 147322 71843
rect 147259 10436 147325 10437
rect 147259 10372 147260 10436
rect 147324 10372 147325 10436
rect 147259 10371 147325 10372
rect 147446 10301 147506 71843
rect 148366 21589 148426 72523
rect 148547 72452 148613 72453
rect 148547 72388 148548 72452
rect 148612 72388 148613 72452
rect 148547 72387 148613 72388
rect 148363 21588 148429 21589
rect 148363 21524 148364 21588
rect 148428 21524 148429 21588
rect 148363 21523 148429 21524
rect 148550 16149 148610 72387
rect 148547 16148 148613 16149
rect 148547 16084 148548 16148
rect 148612 16084 148613 16148
rect 148547 16083 148613 16084
rect 148734 11933 148794 72795
rect 148915 72724 148981 72725
rect 148915 72660 148916 72724
rect 148980 72660 148981 72724
rect 148915 72659 148981 72660
rect 148918 12069 148978 72659
rect 149470 26893 149530 72931
rect 149835 72860 149901 72861
rect 149835 72796 149836 72860
rect 149900 72796 149901 72860
rect 149835 72795 149901 72796
rect 149651 72588 149717 72589
rect 149651 72524 149652 72588
rect 149716 72524 149717 72588
rect 149651 72523 149717 72524
rect 149467 26892 149533 26893
rect 149467 26828 149468 26892
rect 149532 26828 149533 26892
rect 149467 26827 149533 26828
rect 149654 13429 149714 72523
rect 149651 13428 149717 13429
rect 149651 13364 149652 13428
rect 149716 13364 149717 13428
rect 149651 13363 149717 13364
rect 149838 13293 149898 72795
rect 150019 72724 150085 72725
rect 150019 72660 150020 72724
rect 150084 72660 150085 72724
rect 150019 72659 150085 72660
rect 149835 13292 149901 13293
rect 149835 13228 149836 13292
rect 149900 13228 149901 13292
rect 149835 13227 149901 13228
rect 148915 12068 148981 12069
rect 148915 12004 148916 12068
rect 148980 12004 148981 12068
rect 148915 12003 148981 12004
rect 148731 11932 148797 11933
rect 148731 11868 148732 11932
rect 148796 11868 148797 11932
rect 148731 11867 148797 11868
rect 150022 11797 150082 72659
rect 150294 43954 150914 73000
rect 153883 72996 153949 72997
rect 153883 72932 153884 72996
rect 153948 72932 153949 72996
rect 153883 72931 153949 72932
rect 151491 72860 151557 72861
rect 151491 72796 151492 72860
rect 151556 72796 151557 72860
rect 151491 72795 151557 72796
rect 152779 72860 152845 72861
rect 152779 72796 152780 72860
rect 152844 72796 152845 72860
rect 152779 72795 152845 72796
rect 151307 72452 151373 72453
rect 151307 72388 151308 72452
rect 151372 72388 151373 72452
rect 151307 72387 151373 72388
rect 150294 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 150914 43954
rect 150294 43634 150914 43718
rect 150294 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 150914 43634
rect 150019 11796 150085 11797
rect 150019 11732 150020 11796
rect 150084 11732 150085 11796
rect 150019 11731 150085 11732
rect 147443 10300 147509 10301
rect 147443 10236 147444 10300
rect 147508 10236 147509 10300
rect 147443 10235 147509 10236
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 150294 7954 150914 43398
rect 151310 24445 151370 72387
rect 151307 24444 151373 24445
rect 151307 24380 151308 24444
rect 151372 24380 151373 24444
rect 151307 24379 151373 24380
rect 151494 14653 151554 72795
rect 151675 72724 151741 72725
rect 151675 72660 151676 72724
rect 151740 72660 151741 72724
rect 151675 72659 151741 72660
rect 151491 14652 151557 14653
rect 151491 14588 151492 14652
rect 151556 14588 151557 14652
rect 151491 14587 151557 14588
rect 150294 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 150914 7954
rect 150294 7634 150914 7718
rect 150294 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 150914 7634
rect 150294 -1306 150914 7398
rect 151678 6493 151738 72659
rect 152411 72588 152477 72589
rect 152411 72524 152412 72588
rect 152476 72524 152477 72588
rect 152411 72523 152477 72524
rect 152414 16013 152474 72523
rect 152595 72452 152661 72453
rect 152595 72388 152596 72452
rect 152660 72388 152661 72452
rect 152595 72387 152661 72388
rect 152411 16012 152477 16013
rect 152411 15948 152412 16012
rect 152476 15948 152477 16012
rect 152411 15947 152477 15948
rect 152598 14517 152658 72387
rect 152595 14516 152661 14517
rect 152595 14452 152596 14516
rect 152660 14452 152661 14516
rect 152595 14451 152661 14452
rect 152782 11661 152842 72795
rect 152963 72724 153029 72725
rect 152963 72660 152964 72724
rect 153028 72660 153029 72724
rect 152963 72659 153029 72660
rect 152779 11660 152845 11661
rect 152779 11596 152780 11660
rect 152844 11596 152845 11660
rect 152779 11595 152845 11596
rect 151675 6492 151741 6493
rect 151675 6428 151676 6492
rect 151740 6428 151741 6492
rect 151675 6427 151741 6428
rect 152966 5541 153026 72659
rect 153886 17509 153946 72931
rect 154435 72860 154501 72861
rect 154435 72796 154436 72860
rect 154500 72796 154501 72860
rect 154435 72795 154501 72796
rect 154251 72724 154317 72725
rect 154251 72660 154252 72724
rect 154316 72660 154317 72724
rect 154251 72659 154317 72660
rect 154067 72588 154133 72589
rect 154067 72524 154068 72588
rect 154132 72524 154133 72588
rect 154067 72523 154133 72524
rect 153883 17508 153949 17509
rect 153883 17444 153884 17508
rect 153948 17444 153949 17508
rect 153883 17443 153949 17444
rect 154070 17373 154130 72523
rect 154067 17372 154133 17373
rect 154067 17308 154068 17372
rect 154132 17308 154133 17372
rect 154067 17307 154133 17308
rect 154254 15877 154314 72659
rect 154251 15876 154317 15877
rect 154251 15812 154252 15876
rect 154316 15812 154317 15876
rect 154251 15811 154317 15812
rect 154438 13157 154498 72795
rect 154794 48454 155414 73000
rect 155539 72860 155605 72861
rect 155539 72796 155540 72860
rect 155604 72796 155605 72860
rect 155539 72795 155605 72796
rect 157195 72860 157261 72861
rect 157195 72796 157196 72860
rect 157260 72796 157261 72860
rect 157195 72795 157261 72796
rect 158299 72860 158365 72861
rect 158299 72796 158300 72860
rect 158364 72796 158365 72860
rect 158299 72795 158365 72796
rect 158851 72860 158917 72861
rect 158851 72796 158852 72860
rect 158916 72796 158917 72860
rect 158851 72795 158917 72796
rect 154794 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 155414 48454
rect 154794 48134 155414 48218
rect 154794 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 155414 48134
rect 154435 13156 154501 13157
rect 154435 13092 154436 13156
rect 154500 13092 154501 13156
rect 154435 13091 154501 13092
rect 154794 12454 155414 47898
rect 155542 21453 155602 72795
rect 155723 72724 155789 72725
rect 155723 72660 155724 72724
rect 155788 72660 155789 72724
rect 155723 72659 155789 72660
rect 156827 72724 156893 72725
rect 156827 72660 156828 72724
rect 156892 72660 156893 72724
rect 156827 72659 156893 72660
rect 157011 72724 157077 72725
rect 157011 72660 157012 72724
rect 157076 72660 157077 72724
rect 157011 72659 157077 72660
rect 155539 21452 155605 21453
rect 155539 21388 155540 21452
rect 155604 21388 155605 21452
rect 155539 21387 155605 21388
rect 155726 17237 155786 72659
rect 156643 72588 156709 72589
rect 156643 72524 156644 72588
rect 156708 72524 156709 72588
rect 156643 72523 156709 72524
rect 156646 25533 156706 72523
rect 156643 25532 156709 25533
rect 156643 25468 156644 25532
rect 156708 25468 156709 25532
rect 156643 25467 156709 25468
rect 156830 22813 156890 72659
rect 156827 22812 156893 22813
rect 156827 22748 156828 22812
rect 156892 22748 156893 22812
rect 156827 22747 156893 22748
rect 157014 18733 157074 72659
rect 157198 18869 157258 72795
rect 158115 72588 158181 72589
rect 158115 72524 158116 72588
rect 158180 72524 158181 72588
rect 158115 72523 158181 72524
rect 158118 31109 158178 72523
rect 158115 31108 158181 31109
rect 158115 31044 158116 31108
rect 158180 31044 158181 31108
rect 158115 31043 158181 31044
rect 158302 21317 158362 72795
rect 158483 72724 158549 72725
rect 158483 72660 158484 72724
rect 158548 72660 158549 72724
rect 158483 72659 158549 72660
rect 158299 21316 158365 21317
rect 158299 21252 158300 21316
rect 158364 21252 158365 21316
rect 158299 21251 158365 21252
rect 158486 19957 158546 72659
rect 158667 72452 158733 72453
rect 158667 72388 158668 72452
rect 158732 72388 158733 72452
rect 158667 72387 158733 72388
rect 158670 65517 158730 72387
rect 158667 65516 158733 65517
rect 158667 65452 158668 65516
rect 158732 65452 158733 65516
rect 158667 65451 158733 65452
rect 158854 30973 158914 72795
rect 159035 72724 159101 72725
rect 159035 72660 159036 72724
rect 159100 72660 159101 72724
rect 159035 72659 159101 72660
rect 158851 30972 158917 30973
rect 158851 30908 158852 30972
rect 158916 30908 158917 30972
rect 158851 30907 158917 30908
rect 158483 19956 158549 19957
rect 158483 19892 158484 19956
rect 158548 19892 158549 19956
rect 158483 19891 158549 19892
rect 157195 18868 157261 18869
rect 157195 18804 157196 18868
rect 157260 18804 157261 18868
rect 157195 18803 157261 18804
rect 157011 18732 157077 18733
rect 157011 18668 157012 18732
rect 157076 18668 157077 18732
rect 157011 18667 157077 18668
rect 155723 17236 155789 17237
rect 155723 17172 155724 17236
rect 155788 17172 155789 17236
rect 155723 17171 155789 17172
rect 154794 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 155414 12454
rect 154794 12134 155414 12218
rect 154794 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 155414 12134
rect 152963 5540 153029 5541
rect 152963 5476 152964 5540
rect 153028 5476 153029 5540
rect 152963 5475 153029 5476
rect 150294 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 150914 -1306
rect 150294 -1626 150914 -1542
rect 150294 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 150914 -1626
rect 150294 -7654 150914 -1862
rect 154794 -2266 155414 11898
rect 159038 4045 159098 72659
rect 159294 52954 159914 73000
rect 162163 72996 162229 72997
rect 162163 72932 162164 72996
rect 162228 72932 162229 72996
rect 162163 72931 162229 72932
rect 160691 72860 160757 72861
rect 160691 72796 160692 72860
rect 160756 72796 160757 72860
rect 160691 72795 160757 72796
rect 159294 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 159914 52954
rect 159294 52634 159914 52718
rect 159294 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 159914 52634
rect 159294 16954 159914 52398
rect 160694 22677 160754 72795
rect 160875 72724 160941 72725
rect 160875 72660 160876 72724
rect 160940 72660 160941 72724
rect 160875 72659 160941 72660
rect 160691 22676 160757 22677
rect 160691 22612 160692 22676
rect 160756 22612 160757 22676
rect 160691 22611 160757 22612
rect 159294 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 159914 16954
rect 159294 16634 159914 16718
rect 159294 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 159914 16634
rect 159035 4044 159101 4045
rect 159035 3980 159036 4044
rect 159100 3980 159101 4044
rect 159035 3979 159101 3980
rect 154794 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 155414 -2266
rect 154794 -2586 155414 -2502
rect 154794 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 155414 -2586
rect 154794 -7654 155414 -2822
rect 159294 -3226 159914 16398
rect 160878 13021 160938 72659
rect 161059 72588 161125 72589
rect 161059 72524 161060 72588
rect 161124 72524 161125 72588
rect 161059 72523 161125 72524
rect 160875 13020 160941 13021
rect 160875 12956 160876 13020
rect 160940 12956 160941 13020
rect 160875 12955 160941 12956
rect 161062 5269 161122 72523
rect 161243 72452 161309 72453
rect 161243 72388 161244 72452
rect 161308 72388 161309 72452
rect 161243 72387 161309 72388
rect 161246 5405 161306 72387
rect 162166 24309 162226 72931
rect 162531 72860 162597 72861
rect 162531 72796 162532 72860
rect 162596 72796 162597 72860
rect 162531 72795 162597 72796
rect 162347 72588 162413 72589
rect 162347 72524 162348 72588
rect 162412 72524 162413 72588
rect 162347 72523 162413 72524
rect 162163 24308 162229 24309
rect 162163 24244 162164 24308
rect 162228 24244 162229 24308
rect 162163 24243 162229 24244
rect 162350 18597 162410 72523
rect 162347 18596 162413 18597
rect 162347 18532 162348 18596
rect 162412 18532 162413 18596
rect 162347 18531 162413 18532
rect 162534 6221 162594 72795
rect 162715 72724 162781 72725
rect 162715 72660 162716 72724
rect 162780 72660 162781 72724
rect 162715 72659 162781 72660
rect 162718 6357 162778 72659
rect 162902 72453 162962 74835
rect 167502 74765 167562 75110
rect 168422 75037 168482 75379
rect 168606 75309 168666 75790
rect 168603 75308 168669 75309
rect 168603 75244 168604 75308
rect 168668 75244 168669 75308
rect 168603 75243 168669 75244
rect 168603 75172 168669 75173
rect 168603 75108 168604 75172
rect 168668 75170 168669 75172
rect 168668 75110 169218 75170
rect 168668 75108 168669 75110
rect 168603 75107 168669 75108
rect 168419 75036 168485 75037
rect 168419 74972 168420 75036
rect 168484 74972 168485 75036
rect 168419 74971 168485 74972
rect 169158 74901 169218 75110
rect 169155 74900 169221 74901
rect 169155 74836 169156 74900
rect 169220 74836 169221 74900
rect 169155 74835 169221 74836
rect 169342 74765 169402 75790
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 167499 74764 167565 74765
rect 167499 74700 167500 74764
rect 167564 74700 167565 74764
rect 167499 74699 167565 74700
rect 169339 74764 169405 74765
rect 169339 74700 169340 74764
rect 169404 74700 169405 74764
rect 169339 74699 169405 74700
rect 167499 73132 167565 73133
rect 167499 73068 167500 73132
rect 167564 73068 167565 73132
rect 167499 73067 167565 73068
rect 163267 72860 163333 72861
rect 163267 72796 163268 72860
rect 163332 72796 163333 72860
rect 163267 72795 163333 72796
rect 162899 72452 162965 72453
rect 162899 72388 162900 72452
rect 162964 72388 162965 72452
rect 162899 72387 162965 72388
rect 163270 31245 163330 72795
rect 163451 72724 163517 72725
rect 163451 72660 163452 72724
rect 163516 72660 163517 72724
rect 163451 72659 163517 72660
rect 163267 31244 163333 31245
rect 163267 31180 163268 31244
rect 163332 31180 163333 31244
rect 163267 31179 163333 31180
rect 163454 24173 163514 72659
rect 163635 72452 163701 72453
rect 163635 72388 163636 72452
rect 163700 72388 163701 72452
rect 163635 72387 163701 72388
rect 163451 24172 163517 24173
rect 163451 24108 163452 24172
rect 163516 24108 163517 24172
rect 163451 24107 163517 24108
rect 162715 6356 162781 6357
rect 162715 6292 162716 6356
rect 162780 6292 162781 6356
rect 162715 6291 162781 6292
rect 162531 6220 162597 6221
rect 162531 6156 162532 6220
rect 162596 6156 162597 6220
rect 162531 6155 162597 6156
rect 161243 5404 161309 5405
rect 161243 5340 161244 5404
rect 161308 5340 161309 5404
rect 161243 5339 161309 5340
rect 161059 5268 161125 5269
rect 161059 5204 161060 5268
rect 161124 5204 161125 5268
rect 161059 5203 161125 5204
rect 163638 5133 163698 72387
rect 163794 57454 164414 73000
rect 165291 72860 165357 72861
rect 165291 72796 165292 72860
rect 165356 72796 165357 72860
rect 165291 72795 165357 72796
rect 165107 72724 165173 72725
rect 165107 72660 165108 72724
rect 165172 72660 165173 72724
rect 165107 72659 165173 72660
rect 164923 72588 164989 72589
rect 164923 72524 164924 72588
rect 164988 72524 164989 72588
rect 164923 72523 164989 72524
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163635 5132 163701 5133
rect 163635 5068 163636 5132
rect 163700 5068 163701 5132
rect 163635 5067 163701 5068
rect 159294 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 159914 -3226
rect 159294 -3546 159914 -3462
rect 159294 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 159914 -3546
rect 159294 -7654 159914 -3782
rect 163794 -4186 164414 20898
rect 164926 7581 164986 72523
rect 165110 7717 165170 72659
rect 165107 7716 165173 7717
rect 165107 7652 165108 7716
rect 165172 7652 165173 7716
rect 165107 7651 165173 7652
rect 164923 7580 164989 7581
rect 164923 7516 164924 7580
rect 164988 7516 164989 7580
rect 164923 7515 164989 7516
rect 165294 4861 165354 72795
rect 166211 72724 166277 72725
rect 166211 72660 166212 72724
rect 166276 72660 166277 72724
rect 166211 72659 166277 72660
rect 166763 72724 166829 72725
rect 166763 72660 166764 72724
rect 166828 72660 166829 72724
rect 166763 72659 166829 72660
rect 166947 72724 167013 72725
rect 166947 72660 166948 72724
rect 167012 72660 167013 72724
rect 166947 72659 167013 72660
rect 165475 72452 165541 72453
rect 165475 72388 165476 72452
rect 165540 72388 165541 72452
rect 165475 72387 165541 72388
rect 165478 4997 165538 72387
rect 166214 31789 166274 72659
rect 166579 72588 166645 72589
rect 166579 72524 166580 72588
rect 166644 72524 166645 72588
rect 166579 72523 166645 72524
rect 166395 72452 166461 72453
rect 166395 72388 166396 72452
rect 166460 72388 166461 72452
rect 166395 72387 166461 72388
rect 166211 31788 166277 31789
rect 166211 31724 166212 31788
rect 166276 31724 166277 31788
rect 166211 31723 166277 31724
rect 166398 8941 166458 72387
rect 166582 9077 166642 72523
rect 166579 9076 166645 9077
rect 166579 9012 166580 9076
rect 166644 9012 166645 9076
rect 166579 9011 166645 9012
rect 166395 8940 166461 8941
rect 166395 8876 166396 8940
rect 166460 8876 166461 8940
rect 166395 8875 166461 8876
rect 165475 4996 165541 4997
rect 165475 4932 165476 4996
rect 165540 4932 165541 4996
rect 165475 4931 165541 4932
rect 165291 4860 165357 4861
rect 165291 4796 165292 4860
rect 165356 4796 165357 4860
rect 165291 4795 165357 4796
rect 166766 3365 166826 72659
rect 166950 71909 167010 72659
rect 166947 71908 167013 71909
rect 166947 71844 166948 71908
rect 167012 71844 167013 71908
rect 166947 71843 167013 71844
rect 167502 3773 167562 73067
rect 167683 72996 167749 72997
rect 167683 72932 167684 72996
rect 167748 72932 167749 72996
rect 167683 72931 167749 72932
rect 167499 3772 167565 3773
rect 167499 3708 167500 3772
rect 167564 3708 167565 3772
rect 167499 3707 167565 3708
rect 167686 3637 167746 72931
rect 167867 72860 167933 72861
rect 167867 72796 167868 72860
rect 167932 72796 167933 72860
rect 167867 72795 167933 72796
rect 167683 3636 167749 3637
rect 167683 3572 167684 3636
rect 167748 3572 167749 3636
rect 167683 3571 167749 3572
rect 167870 3501 167930 72795
rect 168294 61954 168914 73000
rect 168294 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 168914 61954
rect 168294 61634 168914 61718
rect 168294 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 168914 61634
rect 168294 25954 168914 61398
rect 168294 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 168914 25954
rect 168294 25634 168914 25718
rect 168294 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 168914 25634
rect 167867 3500 167933 3501
rect 167867 3436 167868 3500
rect 167932 3436 167933 3500
rect 167867 3435 167933 3436
rect 166763 3364 166829 3365
rect 166763 3300 166764 3364
rect 166828 3300 166829 3364
rect 166763 3299 166829 3300
rect 163794 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 164414 -4186
rect 163794 -4506 164414 -4422
rect 163794 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 164414 -4506
rect 163794 -7654 164414 -4742
rect 168294 -5146 168914 25398
rect 168294 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 168914 -5146
rect 168294 -5466 168914 -5382
rect 168294 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 168914 -5466
rect 168294 -7654 168914 -5702
rect 172794 66454 173414 73000
rect 172794 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 173414 66454
rect 172794 66134 173414 66218
rect 172794 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 173414 66134
rect 172794 30454 173414 65898
rect 172794 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 173414 30454
rect 172794 30134 173414 30218
rect 172794 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 173414 30134
rect 172794 -6106 173414 29898
rect 172794 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 173414 -6106
rect 172794 -6426 173414 -6342
rect 172794 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 173414 -6426
rect 172794 -7654 173414 -6662
rect 177294 70954 177914 73000
rect 177294 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 177914 70954
rect 177294 70634 177914 70718
rect 177294 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 177914 70634
rect 177294 34954 177914 70398
rect 177294 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 177914 34954
rect 177294 34634 177914 34718
rect 177294 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 177914 34634
rect 177294 -7066 177914 34398
rect 177294 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 177914 -7066
rect 177294 -7386 177914 -7302
rect 177294 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 177914 -7386
rect 177294 -7654 177914 -7622
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 186294 223954 186914 228484
rect 186294 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 186914 223954
rect 186294 223634 186914 223718
rect 186294 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 186914 223634
rect 186294 187954 186914 223398
rect 186294 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 186914 187954
rect 186294 187634 186914 187718
rect 186294 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 186914 187634
rect 186294 151954 186914 187398
rect 186294 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 186914 151954
rect 186294 151634 186914 151718
rect 186294 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 186914 151634
rect 186294 115954 186914 151398
rect 186294 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 186914 115954
rect 186294 115634 186914 115718
rect 186294 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 186914 115634
rect 186294 79954 186914 115398
rect 186294 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 186914 79954
rect 186294 79634 186914 79718
rect 186294 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 186914 79634
rect 186294 43954 186914 79398
rect 186294 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 186914 43954
rect 186294 43634 186914 43718
rect 186294 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 186914 43634
rect 186294 7954 186914 43398
rect 186294 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 186914 7954
rect 186294 7634 186914 7718
rect 186294 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 186914 7634
rect 186294 -1306 186914 7398
rect 186294 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 186914 -1306
rect 186294 -1626 186914 -1542
rect 186294 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 186914 -1626
rect 186294 -7654 186914 -1862
rect 190794 228453 191414 228484
rect 190794 228217 190826 228453
rect 191062 228217 191146 228453
rect 191382 228217 191414 228453
rect 190794 228133 191414 228217
rect 190794 227897 190826 228133
rect 191062 227897 191146 228133
rect 191382 227897 191414 228133
rect 190794 192454 191414 227897
rect 190794 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 191414 192454
rect 190794 192134 191414 192218
rect 190794 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 191414 192134
rect 190794 156454 191414 191898
rect 190794 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 191414 156454
rect 190794 156134 191414 156218
rect 190794 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 191414 156134
rect 190794 120454 191414 155898
rect 190794 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 191414 120454
rect 190794 120134 191414 120218
rect 190794 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 191414 120134
rect 190794 84454 191414 119898
rect 190794 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 191414 84454
rect 190794 84134 191414 84218
rect 190794 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 191414 84134
rect 190794 48454 191414 83898
rect 190794 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 191414 48454
rect 190794 48134 191414 48218
rect 190794 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 191414 48134
rect 190794 12454 191414 47898
rect 190794 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 191414 12454
rect 190794 12134 191414 12218
rect 190794 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 191414 12134
rect 190794 -2266 191414 11898
rect 190794 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 191414 -2266
rect 190794 -2586 191414 -2502
rect 190794 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 191414 -2586
rect 190794 -7654 191414 -2822
rect 195294 196954 195914 228484
rect 195294 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 195914 196954
rect 195294 196634 195914 196718
rect 195294 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 195914 196634
rect 195294 160954 195914 196398
rect 195294 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 195914 160954
rect 195294 160634 195914 160718
rect 195294 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 195914 160634
rect 195294 124954 195914 160398
rect 195294 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 195914 124954
rect 195294 124634 195914 124718
rect 195294 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 195914 124634
rect 195294 88954 195914 124398
rect 195294 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 195914 88954
rect 195294 88634 195914 88718
rect 195294 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 195914 88634
rect 195294 52954 195914 88398
rect 195294 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 195914 52954
rect 195294 52634 195914 52718
rect 195294 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 195914 52634
rect 195294 16954 195914 52398
rect 195294 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 195914 16954
rect 195294 16634 195914 16718
rect 195294 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 195914 16634
rect 195294 -3226 195914 16398
rect 195294 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 195914 -3226
rect 195294 -3546 195914 -3462
rect 195294 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 195914 -3546
rect 195294 -7654 195914 -3782
rect 199794 201454 200414 228484
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -4186 200414 20898
rect 199794 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 200414 -4186
rect 199794 -4506 200414 -4422
rect 199794 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 200414 -4506
rect 199794 -7654 200414 -4742
rect 204294 205954 204914 228484
rect 204294 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 204914 205954
rect 204294 205634 204914 205718
rect 204294 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 204914 205634
rect 204294 169954 204914 205398
rect 204294 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 204914 169954
rect 204294 169634 204914 169718
rect 204294 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 204914 169634
rect 204294 133954 204914 169398
rect 204294 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 204914 133954
rect 204294 133634 204914 133718
rect 204294 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 204914 133634
rect 204294 97954 204914 133398
rect 204294 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 204914 97954
rect 204294 97634 204914 97718
rect 204294 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 204914 97634
rect 204294 61954 204914 97398
rect 204294 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 204914 61954
rect 204294 61634 204914 61718
rect 204294 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 204914 61634
rect 204294 25954 204914 61398
rect 204294 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 204914 25954
rect 204294 25634 204914 25718
rect 204294 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 204914 25634
rect 204294 -5146 204914 25398
rect 204294 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 204914 -5146
rect 204294 -5466 204914 -5382
rect 204294 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 204914 -5466
rect 204294 -7654 204914 -5702
rect 208794 210454 209414 228484
rect 208794 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 209414 210454
rect 208794 210134 209414 210218
rect 208794 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 209414 210134
rect 208794 174454 209414 209898
rect 208794 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 209414 174454
rect 208794 174134 209414 174218
rect 208794 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 209414 174134
rect 208794 138454 209414 173898
rect 208794 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 209414 138454
rect 208794 138134 209414 138218
rect 208794 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 209414 138134
rect 208794 102454 209414 137898
rect 208794 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 209414 102454
rect 208794 102134 209414 102218
rect 208794 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 209414 102134
rect 208794 66454 209414 101898
rect 208794 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 209414 66454
rect 208794 66134 209414 66218
rect 208794 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 209414 66134
rect 208794 30454 209414 65898
rect 208794 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 209414 30454
rect 208794 30134 209414 30218
rect 208794 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 209414 30134
rect 208794 -6106 209414 29898
rect 208794 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 209414 -6106
rect 208794 -6426 209414 -6342
rect 208794 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 209414 -6426
rect 208794 -7654 209414 -6662
rect 213294 214954 213914 228484
rect 213294 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 213914 214954
rect 213294 214634 213914 214718
rect 213294 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 213914 214634
rect 213294 178954 213914 214398
rect 213294 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 213914 178954
rect 213294 178634 213914 178718
rect 213294 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 213914 178634
rect 213294 142954 213914 178398
rect 213294 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 213914 142954
rect 213294 142634 213914 142718
rect 213294 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 213914 142634
rect 213294 106954 213914 142398
rect 213294 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 213914 106954
rect 213294 106634 213914 106718
rect 213294 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 213914 106634
rect 213294 70954 213914 106398
rect 213294 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 213914 70954
rect 213294 70634 213914 70718
rect 213294 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 213914 70634
rect 213294 34954 213914 70398
rect 213294 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 213914 34954
rect 213294 34634 213914 34718
rect 213294 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 213914 34634
rect 213294 -7066 213914 34398
rect 213294 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 213914 -7066
rect 213294 -7386 213914 -7302
rect 213294 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 213914 -7386
rect 213294 -7654 213914 -7622
rect 217794 219454 218414 228484
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 147454 218414 182898
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 222294 223954 222914 228484
rect 222294 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 222914 223954
rect 222294 223634 222914 223718
rect 222294 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 222914 223634
rect 222294 187954 222914 223398
rect 222294 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 222914 187954
rect 222294 187634 222914 187718
rect 222294 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 222914 187634
rect 222294 151954 222914 187398
rect 222294 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 222914 151954
rect 222294 151634 222914 151718
rect 222294 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 222914 151634
rect 222294 115954 222914 151398
rect 222294 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 222914 115954
rect 222294 115634 222914 115718
rect 222294 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 222914 115634
rect 222294 79954 222914 115398
rect 222294 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 222914 79954
rect 222294 79634 222914 79718
rect 222294 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 222914 79634
rect 222294 43954 222914 79398
rect 222294 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 222914 43954
rect 222294 43634 222914 43718
rect 222294 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 222914 43634
rect 222294 7954 222914 43398
rect 222294 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 222914 7954
rect 222294 7634 222914 7718
rect 222294 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 222914 7634
rect 222294 -1306 222914 7398
rect 222294 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 222914 -1306
rect 222294 -1626 222914 -1542
rect 222294 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 222914 -1626
rect 222294 -7654 222914 -1862
rect 226794 228453 227414 228484
rect 226794 228217 226826 228453
rect 227062 228217 227146 228453
rect 227382 228217 227414 228453
rect 226794 228133 227414 228217
rect 226794 227897 226826 228133
rect 227062 227897 227146 228133
rect 227382 227897 227414 228133
rect 226794 192454 227414 227897
rect 226794 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 227414 192454
rect 226794 192134 227414 192218
rect 226794 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 227414 192134
rect 226794 156454 227414 191898
rect 226794 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 227414 156454
rect 226794 156134 227414 156218
rect 226794 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 227414 156134
rect 226794 120454 227414 155898
rect 226794 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 227414 120454
rect 226794 120134 227414 120218
rect 226794 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 227414 120134
rect 226794 84454 227414 119898
rect 226794 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 227414 84454
rect 226794 84134 227414 84218
rect 226794 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 227414 84134
rect 226794 48454 227414 83898
rect 226794 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 227414 48454
rect 226794 48134 227414 48218
rect 226794 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 227414 48134
rect 226794 12454 227414 47898
rect 226794 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 227414 12454
rect 226794 12134 227414 12218
rect 226794 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 227414 12134
rect 226794 -2266 227414 11898
rect 226794 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 227414 -2266
rect 226794 -2586 227414 -2502
rect 226794 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 227414 -2586
rect 226794 -7654 227414 -2822
rect 231294 196954 231914 228484
rect 231294 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 231914 196954
rect 231294 196634 231914 196718
rect 231294 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 231914 196634
rect 231294 160954 231914 196398
rect 231294 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 231914 160954
rect 231294 160634 231914 160718
rect 231294 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 231914 160634
rect 231294 124954 231914 160398
rect 231294 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 231914 124954
rect 231294 124634 231914 124718
rect 231294 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 231914 124634
rect 231294 88954 231914 124398
rect 231294 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 231914 88954
rect 231294 88634 231914 88718
rect 231294 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 231914 88634
rect 231294 52954 231914 88398
rect 231294 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 231914 52954
rect 231294 52634 231914 52718
rect 231294 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 231914 52634
rect 231294 16954 231914 52398
rect 231294 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 231914 16954
rect 231294 16634 231914 16718
rect 231294 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 231914 16634
rect 231294 -3226 231914 16398
rect 231294 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 231914 -3226
rect 231294 -3546 231914 -3462
rect 231294 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 231914 -3546
rect 231294 -7654 231914 -3782
rect 235794 201454 236414 228484
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 165454 236414 200898
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 235794 129454 236414 164898
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -4186 236414 20898
rect 235794 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 236414 -4186
rect 235794 -4506 236414 -4422
rect 235794 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 236414 -4506
rect 235794 -7654 236414 -4742
rect 240294 205954 240914 228484
rect 240294 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 240914 205954
rect 240294 205634 240914 205718
rect 240294 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 240914 205634
rect 240294 169954 240914 205398
rect 240294 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 240914 169954
rect 240294 169634 240914 169718
rect 240294 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 240914 169634
rect 240294 133954 240914 169398
rect 240294 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 240914 133954
rect 240294 133634 240914 133718
rect 240294 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 240914 133634
rect 240294 97954 240914 133398
rect 240294 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 240914 97954
rect 240294 97634 240914 97718
rect 240294 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 240914 97634
rect 240294 61954 240914 97398
rect 240294 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 240914 61954
rect 240294 61634 240914 61718
rect 240294 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 240914 61634
rect 240294 25954 240914 61398
rect 240294 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 240914 25954
rect 240294 25634 240914 25718
rect 240294 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 240914 25634
rect 240294 -5146 240914 25398
rect 240294 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 240914 -5146
rect 240294 -5466 240914 -5382
rect 240294 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 240914 -5466
rect 240294 -7654 240914 -5702
rect 244794 210454 245414 228484
rect 244794 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 245414 210454
rect 244794 210134 245414 210218
rect 244794 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 245414 210134
rect 244794 174454 245414 209898
rect 244794 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 245414 174454
rect 244794 174134 245414 174218
rect 244794 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 245414 174134
rect 244794 138454 245414 173898
rect 244794 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 245414 138454
rect 244794 138134 245414 138218
rect 244794 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 245414 138134
rect 244794 102454 245414 137898
rect 244794 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 245414 102454
rect 244794 102134 245414 102218
rect 244794 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 245414 102134
rect 244794 66454 245414 101898
rect 244794 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 245414 66454
rect 244794 66134 245414 66218
rect 244794 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 245414 66134
rect 244794 30454 245414 65898
rect 244794 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 245414 30454
rect 244794 30134 245414 30218
rect 244794 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 245414 30134
rect 244794 -6106 245414 29898
rect 244794 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 245414 -6106
rect 244794 -6426 245414 -6342
rect 244794 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 245414 -6426
rect 244794 -7654 245414 -6662
rect 249294 214954 249914 228484
rect 249294 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 249914 214954
rect 249294 214634 249914 214718
rect 249294 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 249914 214634
rect 249294 178954 249914 214398
rect 249294 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 249914 178954
rect 249294 178634 249914 178718
rect 249294 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 249914 178634
rect 249294 142954 249914 178398
rect 249294 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 249914 142954
rect 249294 142634 249914 142718
rect 249294 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 249914 142634
rect 249294 106954 249914 142398
rect 249294 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 249914 106954
rect 249294 106634 249914 106718
rect 249294 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 249914 106634
rect 249294 70954 249914 106398
rect 249294 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 249914 70954
rect 249294 70634 249914 70718
rect 249294 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 249914 70634
rect 249294 34954 249914 70398
rect 249294 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 249914 34954
rect 249294 34634 249914 34718
rect 249294 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 249914 34634
rect 249294 -7066 249914 34398
rect 249294 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 249914 -7066
rect 249294 -7386 249914 -7302
rect 249294 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 249914 -7386
rect 249294 -7654 249914 -7622
rect 253794 219454 254414 228484
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 258294 223954 258914 228484
rect 258294 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 258914 223954
rect 258294 223634 258914 223718
rect 258294 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 258914 223634
rect 258294 187954 258914 223398
rect 258294 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 258914 187954
rect 258294 187634 258914 187718
rect 258294 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 258914 187634
rect 258294 151954 258914 187398
rect 258294 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 258914 151954
rect 258294 151634 258914 151718
rect 258294 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 258914 151634
rect 258294 115954 258914 151398
rect 258294 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 258914 115954
rect 258294 115634 258914 115718
rect 258294 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 258914 115634
rect 258294 79954 258914 115398
rect 258294 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 258914 79954
rect 258294 79634 258914 79718
rect 258294 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 258914 79634
rect 258294 43954 258914 79398
rect 258294 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 258914 43954
rect 258294 43634 258914 43718
rect 258294 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 258914 43634
rect 258294 7954 258914 43398
rect 258294 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 258914 7954
rect 258294 7634 258914 7718
rect 258294 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 258914 7634
rect 258294 -1306 258914 7398
rect 258294 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 258914 -1306
rect 258294 -1626 258914 -1542
rect 258294 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 258914 -1626
rect 258294 -7654 258914 -1862
rect 262794 228453 263414 228484
rect 262794 228217 262826 228453
rect 263062 228217 263146 228453
rect 263382 228217 263414 228453
rect 262794 228133 263414 228217
rect 262794 227897 262826 228133
rect 263062 227897 263146 228133
rect 263382 227897 263414 228133
rect 262794 192454 263414 227897
rect 262794 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 263414 192454
rect 262794 192134 263414 192218
rect 262794 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 263414 192134
rect 262794 156454 263414 191898
rect 262794 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 263414 156454
rect 262794 156134 263414 156218
rect 262794 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 263414 156134
rect 262794 120454 263414 155898
rect 262794 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 263414 120454
rect 262794 120134 263414 120218
rect 262794 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 263414 120134
rect 262794 84454 263414 119898
rect 262794 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 263414 84454
rect 262794 84134 263414 84218
rect 262794 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 263414 84134
rect 262794 48454 263414 83898
rect 262794 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 263414 48454
rect 262794 48134 263414 48218
rect 262794 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 263414 48134
rect 262794 12454 263414 47898
rect 262794 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 263414 12454
rect 262794 12134 263414 12218
rect 262794 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 263414 12134
rect 262794 -2266 263414 11898
rect 262794 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 263414 -2266
rect 262794 -2586 263414 -2502
rect 262794 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 263414 -2586
rect 262794 -7654 263414 -2822
rect 267294 196954 267914 228484
rect 267294 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 267914 196954
rect 267294 196634 267914 196718
rect 267294 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 267914 196634
rect 267294 160954 267914 196398
rect 267294 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 267914 160954
rect 267294 160634 267914 160718
rect 267294 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 267914 160634
rect 267294 124954 267914 160398
rect 267294 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 267914 124954
rect 267294 124634 267914 124718
rect 267294 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 267914 124634
rect 267294 88954 267914 124398
rect 267294 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 267914 88954
rect 267294 88634 267914 88718
rect 267294 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 267914 88634
rect 267294 52954 267914 88398
rect 267294 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 267914 52954
rect 267294 52634 267914 52718
rect 267294 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 267914 52634
rect 267294 16954 267914 52398
rect 267294 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 267914 16954
rect 267294 16634 267914 16718
rect 267294 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 267914 16634
rect 267294 -3226 267914 16398
rect 267294 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 267914 -3226
rect 267294 -3546 267914 -3462
rect 267294 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 267914 -3546
rect 267294 -7654 267914 -3782
rect 271794 201454 272414 228484
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -4186 272414 20898
rect 271794 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 272414 -4186
rect 271794 -4506 272414 -4422
rect 271794 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 272414 -4506
rect 271794 -7654 272414 -4742
rect 276294 205954 276914 228484
rect 276294 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 276914 205954
rect 276294 205634 276914 205718
rect 276294 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 276914 205634
rect 276294 169954 276914 205398
rect 276294 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 276914 169954
rect 276294 169634 276914 169718
rect 276294 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 276914 169634
rect 276294 133954 276914 169398
rect 276294 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 276914 133954
rect 276294 133634 276914 133718
rect 276294 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 276914 133634
rect 276294 97954 276914 133398
rect 276294 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 276914 97954
rect 276294 97634 276914 97718
rect 276294 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 276914 97634
rect 276294 61954 276914 97398
rect 276294 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 276914 61954
rect 276294 61634 276914 61718
rect 276294 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 276914 61634
rect 276294 25954 276914 61398
rect 276294 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 276914 25954
rect 276294 25634 276914 25718
rect 276294 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 276914 25634
rect 276294 -5146 276914 25398
rect 276294 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 276914 -5146
rect 276294 -5466 276914 -5382
rect 276294 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 276914 -5466
rect 276294 -7654 276914 -5702
rect 280794 210454 281414 228484
rect 280794 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 281414 210454
rect 280794 210134 281414 210218
rect 280794 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 281414 210134
rect 280794 174454 281414 209898
rect 280794 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 281414 174454
rect 280794 174134 281414 174218
rect 280794 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 281414 174134
rect 280794 138454 281414 173898
rect 280794 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 281414 138454
rect 280794 138134 281414 138218
rect 280794 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 281414 138134
rect 280794 102454 281414 137898
rect 280794 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 281414 102454
rect 280794 102134 281414 102218
rect 280794 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 281414 102134
rect 280794 66454 281414 101898
rect 280794 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 281414 66454
rect 280794 66134 281414 66218
rect 280794 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 281414 66134
rect 280794 30454 281414 65898
rect 280794 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 281414 30454
rect 280794 30134 281414 30218
rect 280794 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 281414 30134
rect 280794 -6106 281414 29898
rect 280794 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 281414 -6106
rect 280794 -6426 281414 -6342
rect 280794 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 281414 -6426
rect 280794 -7654 281414 -6662
rect 285294 214954 285914 228484
rect 285294 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 285914 214954
rect 285294 214634 285914 214718
rect 285294 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 285914 214634
rect 285294 178954 285914 214398
rect 285294 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 285914 178954
rect 285294 178634 285914 178718
rect 285294 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 285914 178634
rect 285294 142954 285914 178398
rect 285294 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 285914 142954
rect 285294 142634 285914 142718
rect 285294 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 285914 142634
rect 285294 106954 285914 142398
rect 285294 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 285914 106954
rect 285294 106634 285914 106718
rect 285294 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 285914 106634
rect 285294 70954 285914 106398
rect 285294 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 285914 70954
rect 285294 70634 285914 70718
rect 285294 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 285914 70634
rect 285294 34954 285914 70398
rect 285294 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 285914 34954
rect 285294 34634 285914 34718
rect 285294 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 285914 34634
rect 285294 -7066 285914 34398
rect 285294 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 285914 -7066
rect 285294 -7386 285914 -7302
rect 285294 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 285914 -7386
rect 285294 -7654 285914 -7622
rect 289794 219454 290414 228484
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 294294 223954 294914 228484
rect 294294 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 294914 223954
rect 294294 223634 294914 223718
rect 294294 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 294914 223634
rect 294294 187954 294914 223398
rect 294294 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 294914 187954
rect 294294 187634 294914 187718
rect 294294 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 294914 187634
rect 294294 151954 294914 187398
rect 294294 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 294914 151954
rect 294294 151634 294914 151718
rect 294294 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 294914 151634
rect 294294 115954 294914 151398
rect 294294 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 294914 115954
rect 294294 115634 294914 115718
rect 294294 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 294914 115634
rect 294294 79954 294914 115398
rect 294294 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 294914 79954
rect 294294 79634 294914 79718
rect 294294 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 294914 79634
rect 294294 43954 294914 79398
rect 294294 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 294914 43954
rect 294294 43634 294914 43718
rect 294294 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 294914 43634
rect 294294 7954 294914 43398
rect 294294 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 294914 7954
rect 294294 7634 294914 7718
rect 294294 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 294914 7634
rect 294294 -1306 294914 7398
rect 294294 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 294914 -1306
rect 294294 -1626 294914 -1542
rect 294294 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 294914 -1626
rect 294294 -7654 294914 -1862
rect 298794 228453 299414 228484
rect 298794 228217 298826 228453
rect 299062 228217 299146 228453
rect 299382 228217 299414 228453
rect 298794 228133 299414 228217
rect 298794 227897 298826 228133
rect 299062 227897 299146 228133
rect 299382 227897 299414 228133
rect 298794 192454 299414 227897
rect 298794 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 299414 192454
rect 298794 192134 299414 192218
rect 298794 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 299414 192134
rect 298794 156454 299414 191898
rect 298794 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 299414 156454
rect 298794 156134 299414 156218
rect 298794 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 299414 156134
rect 298794 120454 299414 155898
rect 298794 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 299414 120454
rect 298794 120134 299414 120218
rect 298794 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 299414 120134
rect 298794 84454 299414 119898
rect 298794 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 299414 84454
rect 298794 84134 299414 84218
rect 298794 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 299414 84134
rect 298794 48454 299414 83898
rect 298794 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 299414 48454
rect 298794 48134 299414 48218
rect 298794 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 299414 48134
rect 298794 12454 299414 47898
rect 298794 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 299414 12454
rect 298794 12134 299414 12218
rect 298794 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 299414 12134
rect 298794 -2266 299414 11898
rect 298794 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 299414 -2266
rect 298794 -2586 299414 -2502
rect 298794 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 299414 -2586
rect 298794 -7654 299414 -2822
rect 303294 196954 303914 228484
rect 303294 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 303914 196954
rect 303294 196634 303914 196718
rect 303294 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 303914 196634
rect 303294 160954 303914 196398
rect 303294 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 303914 160954
rect 303294 160634 303914 160718
rect 303294 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 303914 160634
rect 303294 124954 303914 160398
rect 303294 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 303914 124954
rect 303294 124634 303914 124718
rect 303294 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 303914 124634
rect 303294 88954 303914 124398
rect 303294 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 303914 88954
rect 303294 88634 303914 88718
rect 303294 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 303914 88634
rect 303294 52954 303914 88398
rect 303294 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 303914 52954
rect 303294 52634 303914 52718
rect 303294 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 303914 52634
rect 303294 16954 303914 52398
rect 303294 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 303914 16954
rect 303294 16634 303914 16718
rect 303294 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 303914 16634
rect 303294 -3226 303914 16398
rect 303294 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 303914 -3226
rect 303294 -3546 303914 -3462
rect 303294 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 303914 -3546
rect 303294 -7654 303914 -3782
rect 307794 201454 308414 228484
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -4186 308414 20898
rect 307794 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 308414 -4186
rect 307794 -4506 308414 -4422
rect 307794 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 308414 -4506
rect 307794 -7654 308414 -4742
rect 312294 205954 312914 228484
rect 312294 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 312914 205954
rect 312294 205634 312914 205718
rect 312294 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 312914 205634
rect 312294 169954 312914 205398
rect 312294 169718 312326 169954
rect 312562 169718 312646 169954
rect 312882 169718 312914 169954
rect 312294 169634 312914 169718
rect 312294 169398 312326 169634
rect 312562 169398 312646 169634
rect 312882 169398 312914 169634
rect 312294 133954 312914 169398
rect 312294 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 312914 133954
rect 312294 133634 312914 133718
rect 312294 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 312914 133634
rect 312294 97954 312914 133398
rect 312294 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 312914 97954
rect 312294 97634 312914 97718
rect 312294 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 312914 97634
rect 312294 61954 312914 97398
rect 312294 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 312914 61954
rect 312294 61634 312914 61718
rect 312294 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 312914 61634
rect 312294 25954 312914 61398
rect 312294 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 312914 25954
rect 312294 25634 312914 25718
rect 312294 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 312914 25634
rect 312294 -5146 312914 25398
rect 312294 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 312914 -5146
rect 312294 -5466 312914 -5382
rect 312294 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 312914 -5466
rect 312294 -7654 312914 -5702
rect 316794 210454 317414 228484
rect 316794 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 317414 210454
rect 316794 210134 317414 210218
rect 316794 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 317414 210134
rect 316794 174454 317414 209898
rect 316794 174218 316826 174454
rect 317062 174218 317146 174454
rect 317382 174218 317414 174454
rect 316794 174134 317414 174218
rect 316794 173898 316826 174134
rect 317062 173898 317146 174134
rect 317382 173898 317414 174134
rect 316794 138454 317414 173898
rect 316794 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 317414 138454
rect 316794 138134 317414 138218
rect 316794 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 317414 138134
rect 316794 102454 317414 137898
rect 316794 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 317414 102454
rect 316794 102134 317414 102218
rect 316794 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 317414 102134
rect 316794 66454 317414 101898
rect 316794 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 317414 66454
rect 316794 66134 317414 66218
rect 316794 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 317414 66134
rect 316794 30454 317414 65898
rect 316794 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 317414 30454
rect 316794 30134 317414 30218
rect 316794 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 317414 30134
rect 316794 -6106 317414 29898
rect 316794 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 317414 -6106
rect 316794 -6426 317414 -6342
rect 316794 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 317414 -6426
rect 316794 -7654 317414 -6662
rect 321294 214954 321914 228484
rect 321294 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 321914 214954
rect 321294 214634 321914 214718
rect 321294 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 321914 214634
rect 321294 178954 321914 214398
rect 321294 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 321914 178954
rect 321294 178634 321914 178718
rect 321294 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 321914 178634
rect 321294 142954 321914 178398
rect 321294 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 321914 142954
rect 321294 142634 321914 142718
rect 321294 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 321914 142634
rect 321294 106954 321914 142398
rect 321294 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 321914 106954
rect 321294 106634 321914 106718
rect 321294 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 321914 106634
rect 321294 70954 321914 106398
rect 321294 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 321914 70954
rect 321294 70634 321914 70718
rect 321294 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 321914 70634
rect 321294 34954 321914 70398
rect 321294 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 321914 34954
rect 321294 34634 321914 34718
rect 321294 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 321914 34634
rect 321294 -7066 321914 34398
rect 321294 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 321914 -7066
rect 321294 -7386 321914 -7302
rect 321294 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 321914 -7386
rect 321294 -7654 321914 -7622
rect 325794 219454 326414 228484
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 330294 223954 330914 228484
rect 330294 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 330914 223954
rect 330294 223634 330914 223718
rect 330294 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 330914 223634
rect 330294 187954 330914 223398
rect 330294 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 330914 187954
rect 330294 187634 330914 187718
rect 330294 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 330914 187634
rect 330294 151954 330914 187398
rect 330294 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 330914 151954
rect 330294 151634 330914 151718
rect 330294 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 330914 151634
rect 330294 115954 330914 151398
rect 330294 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 330914 115954
rect 330294 115634 330914 115718
rect 330294 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 330914 115634
rect 330294 79954 330914 115398
rect 330294 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 330914 79954
rect 330294 79634 330914 79718
rect 330294 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 330914 79634
rect 330294 43954 330914 79398
rect 330294 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 330914 43954
rect 330294 43634 330914 43718
rect 330294 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 330914 43634
rect 330294 7954 330914 43398
rect 330294 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 330914 7954
rect 330294 7634 330914 7718
rect 330294 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 330914 7634
rect 330294 -1306 330914 7398
rect 330294 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 330914 -1306
rect 330294 -1626 330914 -1542
rect 330294 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 330914 -1626
rect 330294 -7654 330914 -1862
rect 334794 228453 335414 228484
rect 334794 228217 334826 228453
rect 335062 228217 335146 228453
rect 335382 228217 335414 228453
rect 334794 228133 335414 228217
rect 334794 227897 334826 228133
rect 335062 227897 335146 228133
rect 335382 227897 335414 228133
rect 334794 192454 335414 227897
rect 334794 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 335414 192454
rect 334794 192134 335414 192218
rect 334794 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 335414 192134
rect 334794 156454 335414 191898
rect 334794 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 335414 156454
rect 334794 156134 335414 156218
rect 334794 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 335414 156134
rect 334794 120454 335414 155898
rect 334794 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 335414 120454
rect 334794 120134 335414 120218
rect 334794 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 335414 120134
rect 334794 84454 335414 119898
rect 334794 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 335414 84454
rect 334794 84134 335414 84218
rect 334794 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 335414 84134
rect 334794 48454 335414 83898
rect 334794 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 335414 48454
rect 334794 48134 335414 48218
rect 334794 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 335414 48134
rect 334794 12454 335414 47898
rect 334794 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 335414 12454
rect 334794 12134 335414 12218
rect 334794 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 335414 12134
rect 334794 -2266 335414 11898
rect 334794 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 335414 -2266
rect 334794 -2586 335414 -2502
rect 334794 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 335414 -2586
rect 334794 -7654 335414 -2822
rect 339294 196954 339914 228484
rect 339294 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 339914 196954
rect 339294 196634 339914 196718
rect 339294 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 339914 196634
rect 339294 160954 339914 196398
rect 339294 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 339914 160954
rect 339294 160634 339914 160718
rect 339294 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 339914 160634
rect 339294 124954 339914 160398
rect 339294 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 339914 124954
rect 339294 124634 339914 124718
rect 339294 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 339914 124634
rect 339294 88954 339914 124398
rect 339294 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 339914 88954
rect 339294 88634 339914 88718
rect 339294 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 339914 88634
rect 339294 52954 339914 88398
rect 339294 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 339914 52954
rect 339294 52634 339914 52718
rect 339294 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 339914 52634
rect 339294 16954 339914 52398
rect 339294 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 339914 16954
rect 339294 16634 339914 16718
rect 339294 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 339914 16634
rect 339294 -3226 339914 16398
rect 339294 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 339914 -3226
rect 339294 -3546 339914 -3462
rect 339294 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 339914 -3546
rect 339294 -7654 339914 -3782
rect 343794 201454 344414 228484
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -4186 344414 20898
rect 343794 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 344414 -4186
rect 343794 -4506 344414 -4422
rect 343794 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 344414 -4506
rect 343794 -7654 344414 -4742
rect 348294 205954 348914 228484
rect 348294 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 348914 205954
rect 348294 205634 348914 205718
rect 348294 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 348914 205634
rect 348294 169954 348914 205398
rect 348294 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 348914 169954
rect 348294 169634 348914 169718
rect 348294 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 348914 169634
rect 348294 133954 348914 169398
rect 348294 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 348914 133954
rect 348294 133634 348914 133718
rect 348294 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 348914 133634
rect 348294 97954 348914 133398
rect 348294 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 348914 97954
rect 348294 97634 348914 97718
rect 348294 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 348914 97634
rect 348294 61954 348914 97398
rect 348294 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 348914 61954
rect 348294 61634 348914 61718
rect 348294 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 348914 61634
rect 348294 25954 348914 61398
rect 348294 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 348914 25954
rect 348294 25634 348914 25718
rect 348294 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 348914 25634
rect 348294 -5146 348914 25398
rect 348294 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 348914 -5146
rect 348294 -5466 348914 -5382
rect 348294 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 348914 -5466
rect 348294 -7654 348914 -5702
rect 352794 210454 353414 228484
rect 352794 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 353414 210454
rect 352794 210134 353414 210218
rect 352794 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 353414 210134
rect 352794 174454 353414 209898
rect 352794 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 353414 174454
rect 352794 174134 353414 174218
rect 352794 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 353414 174134
rect 352794 138454 353414 173898
rect 352794 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 353414 138454
rect 352794 138134 353414 138218
rect 352794 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 353414 138134
rect 352794 102454 353414 137898
rect 352794 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 353414 102454
rect 352794 102134 353414 102218
rect 352794 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 353414 102134
rect 352794 66454 353414 101898
rect 352794 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 353414 66454
rect 352794 66134 353414 66218
rect 352794 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 353414 66134
rect 352794 30454 353414 65898
rect 352794 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 353414 30454
rect 352794 30134 353414 30218
rect 352794 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 353414 30134
rect 352794 -6106 353414 29898
rect 352794 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 353414 -6106
rect 352794 -6426 353414 -6342
rect 352794 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 353414 -6426
rect 352794 -7654 353414 -6662
rect 357294 214954 357914 228484
rect 357294 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 357914 214954
rect 357294 214634 357914 214718
rect 357294 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 357914 214634
rect 357294 178954 357914 214398
rect 357294 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 357914 178954
rect 357294 178634 357914 178718
rect 357294 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 357914 178634
rect 357294 142954 357914 178398
rect 357294 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 357914 142954
rect 357294 142634 357914 142718
rect 357294 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 357914 142634
rect 357294 106954 357914 142398
rect 357294 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 357914 106954
rect 357294 106634 357914 106718
rect 357294 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 357914 106634
rect 357294 70954 357914 106398
rect 357294 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 357914 70954
rect 357294 70634 357914 70718
rect 357294 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 357914 70634
rect 357294 34954 357914 70398
rect 357294 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 357914 34954
rect 357294 34634 357914 34718
rect 357294 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 357914 34634
rect 357294 -7066 357914 34398
rect 357294 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 357914 -7066
rect 357294 -7386 357914 -7302
rect 357294 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 357914 -7386
rect 357294 -7654 357914 -7622
rect 361794 219454 362414 228484
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 366294 223954 366914 228484
rect 366294 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 366914 223954
rect 366294 223634 366914 223718
rect 366294 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 366914 223634
rect 366294 187954 366914 223398
rect 366294 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 366914 187954
rect 366294 187634 366914 187718
rect 366294 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 366914 187634
rect 366294 151954 366914 187398
rect 366294 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 366914 151954
rect 366294 151634 366914 151718
rect 366294 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 366914 151634
rect 366294 115954 366914 151398
rect 366294 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 366914 115954
rect 366294 115634 366914 115718
rect 366294 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 366914 115634
rect 366294 79954 366914 115398
rect 366294 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 366914 79954
rect 366294 79634 366914 79718
rect 366294 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 366914 79634
rect 366294 43954 366914 79398
rect 366294 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 366914 43954
rect 366294 43634 366914 43718
rect 366294 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 366914 43634
rect 366294 7954 366914 43398
rect 366294 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 366914 7954
rect 366294 7634 366914 7718
rect 366294 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 366914 7634
rect 366294 -1306 366914 7398
rect 366294 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 366914 -1306
rect 366294 -1626 366914 -1542
rect 366294 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 366914 -1626
rect 366294 -7654 366914 -1862
rect 370794 228453 371414 228484
rect 370794 228217 370826 228453
rect 371062 228217 371146 228453
rect 371382 228217 371414 228453
rect 370794 228133 371414 228217
rect 370794 227897 370826 228133
rect 371062 227897 371146 228133
rect 371382 227897 371414 228133
rect 370794 192454 371414 227897
rect 370794 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 371414 192454
rect 370794 192134 371414 192218
rect 370794 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 371414 192134
rect 370794 156454 371414 191898
rect 370794 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 371414 156454
rect 370794 156134 371414 156218
rect 370794 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 371414 156134
rect 370794 120454 371414 155898
rect 370794 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 371414 120454
rect 370794 120134 371414 120218
rect 370794 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 371414 120134
rect 370794 84454 371414 119898
rect 370794 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 371414 84454
rect 370794 84134 371414 84218
rect 370794 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 371414 84134
rect 370794 48454 371414 83898
rect 370794 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 371414 48454
rect 370794 48134 371414 48218
rect 370794 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 371414 48134
rect 370794 12454 371414 47898
rect 370794 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 371414 12454
rect 370794 12134 371414 12218
rect 370794 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 371414 12134
rect 370794 -2266 371414 11898
rect 370794 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 371414 -2266
rect 370794 -2586 371414 -2502
rect 370794 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 371414 -2586
rect 370794 -7654 371414 -2822
rect 375294 196954 375914 228484
rect 375294 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 375914 196954
rect 375294 196634 375914 196718
rect 375294 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 375914 196634
rect 375294 160954 375914 196398
rect 375294 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 375914 160954
rect 375294 160634 375914 160718
rect 375294 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 375914 160634
rect 375294 124954 375914 160398
rect 375294 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 375914 124954
rect 375294 124634 375914 124718
rect 375294 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 375914 124634
rect 375294 88954 375914 124398
rect 375294 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 375914 88954
rect 375294 88634 375914 88718
rect 375294 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 375914 88634
rect 375294 52954 375914 88398
rect 375294 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 375914 52954
rect 375294 52634 375914 52718
rect 375294 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 375914 52634
rect 375294 16954 375914 52398
rect 375294 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 375914 16954
rect 375294 16634 375914 16718
rect 375294 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 375914 16634
rect 375294 -3226 375914 16398
rect 375294 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 375914 -3226
rect 375294 -3546 375914 -3462
rect 375294 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 375914 -3546
rect 375294 -7654 375914 -3782
rect 379794 201454 380414 228484
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -4186 380414 20898
rect 379794 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 380414 -4186
rect 379794 -4506 380414 -4422
rect 379794 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 380414 -4506
rect 379794 -7654 380414 -4742
rect 384294 205954 384914 228484
rect 384294 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 384914 205954
rect 384294 205634 384914 205718
rect 384294 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 384914 205634
rect 384294 169954 384914 205398
rect 384294 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 384914 169954
rect 384294 169634 384914 169718
rect 384294 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 384914 169634
rect 384294 133954 384914 169398
rect 384294 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 384914 133954
rect 384294 133634 384914 133718
rect 384294 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 384914 133634
rect 384294 97954 384914 133398
rect 384294 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 384914 97954
rect 384294 97634 384914 97718
rect 384294 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 384914 97634
rect 384294 61954 384914 97398
rect 384294 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 384914 61954
rect 384294 61634 384914 61718
rect 384294 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 384914 61634
rect 384294 25954 384914 61398
rect 384294 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 384914 25954
rect 384294 25634 384914 25718
rect 384294 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 384914 25634
rect 384294 -5146 384914 25398
rect 384294 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 384914 -5146
rect 384294 -5466 384914 -5382
rect 384294 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 384914 -5466
rect 384294 -7654 384914 -5702
rect 388794 210454 389414 228484
rect 388794 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 389414 210454
rect 388794 210134 389414 210218
rect 388794 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 389414 210134
rect 388794 174454 389414 209898
rect 388794 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 389414 174454
rect 388794 174134 389414 174218
rect 388794 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 389414 174134
rect 388794 138454 389414 173898
rect 388794 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 389414 138454
rect 388794 138134 389414 138218
rect 388794 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 389414 138134
rect 388794 102454 389414 137898
rect 388794 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 389414 102454
rect 388794 102134 389414 102218
rect 388794 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 389414 102134
rect 388794 66454 389414 101898
rect 388794 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 389414 66454
rect 388794 66134 389414 66218
rect 388794 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 389414 66134
rect 388794 30454 389414 65898
rect 388794 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 389414 30454
rect 388794 30134 389414 30218
rect 388794 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 389414 30134
rect 388794 -6106 389414 29898
rect 388794 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 389414 -6106
rect 388794 -6426 389414 -6342
rect 388794 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 389414 -6426
rect 388794 -7654 389414 -6662
rect 393294 214954 393914 228484
rect 393294 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 393914 214954
rect 393294 214634 393914 214718
rect 393294 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 393914 214634
rect 393294 178954 393914 214398
rect 393294 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 393914 178954
rect 393294 178634 393914 178718
rect 393294 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 393914 178634
rect 393294 142954 393914 178398
rect 393294 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 393914 142954
rect 393294 142634 393914 142718
rect 393294 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 393914 142634
rect 393294 106954 393914 142398
rect 396582 137325 396642 470595
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 248684 398414 254898
rect 402294 705798 402914 711590
rect 402294 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 402914 705798
rect 402294 705478 402914 705562
rect 402294 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 402914 705478
rect 402294 691954 402914 705242
rect 402294 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 402914 691954
rect 402294 691634 402914 691718
rect 402294 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 402914 691634
rect 402294 655954 402914 691398
rect 402294 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 402914 655954
rect 402294 655634 402914 655718
rect 402294 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 402914 655634
rect 402294 619954 402914 655398
rect 402294 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 402914 619954
rect 402294 619634 402914 619718
rect 402294 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 402914 619634
rect 402294 583954 402914 619398
rect 402294 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 402914 583954
rect 402294 583634 402914 583718
rect 402294 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 402914 583634
rect 402294 547954 402914 583398
rect 402294 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 402914 547954
rect 402294 547634 402914 547718
rect 402294 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 402914 547634
rect 402294 511954 402914 547398
rect 402294 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 402914 511954
rect 402294 511634 402914 511718
rect 402294 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 402914 511634
rect 402294 475954 402914 511398
rect 402294 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 402914 475954
rect 402294 475634 402914 475718
rect 402294 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 402914 475634
rect 402294 439954 402914 475398
rect 402294 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 402914 439954
rect 402294 439634 402914 439718
rect 402294 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 402914 439634
rect 402294 403954 402914 439398
rect 402294 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 402914 403954
rect 402294 403634 402914 403718
rect 402294 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 402914 403634
rect 402294 367954 402914 403398
rect 402294 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 402914 367954
rect 402294 367634 402914 367718
rect 402294 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 402914 367634
rect 402294 331954 402914 367398
rect 402294 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 402914 331954
rect 402294 331634 402914 331718
rect 402294 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 402914 331634
rect 402294 295954 402914 331398
rect 402294 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 402914 295954
rect 402294 295634 402914 295718
rect 402294 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 402914 295634
rect 402294 259954 402914 295398
rect 402294 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 402914 259954
rect 402294 259634 402914 259718
rect 402294 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 402914 259634
rect 396763 240140 396829 240141
rect 396763 240076 396764 240140
rect 396828 240076 396829 240140
rect 396763 240075 396829 240076
rect 396766 232117 396826 240075
rect 396947 240004 397013 240005
rect 396947 239940 396948 240004
rect 397012 239940 397013 240004
rect 396947 239939 397013 239940
rect 396763 232116 396829 232117
rect 396763 232052 396764 232116
rect 396828 232052 396829 232116
rect 396763 232051 396829 232052
rect 396950 231165 397010 239939
rect 396947 231164 397013 231165
rect 396947 231100 396948 231164
rect 397012 231100 397013 231164
rect 396947 231099 397013 231100
rect 397794 219454 398414 228484
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 396579 137324 396645 137325
rect 396579 137260 396580 137324
rect 396644 137260 396645 137324
rect 396579 137259 396645 137260
rect 393294 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 393914 106954
rect 393294 106634 393914 106718
rect 393294 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 393914 106634
rect 393294 70954 393914 106398
rect 393294 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 393914 70954
rect 393294 70634 393914 70718
rect 393294 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 393914 70634
rect 393294 34954 393914 70398
rect 393294 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 393914 34954
rect 393294 34634 393914 34718
rect 393294 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 393914 34634
rect 393294 -7066 393914 34398
rect 393294 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 393914 -7066
rect 393294 -7386 393914 -7302
rect 393294 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 393914 -7386
rect 393294 -7654 393914 -7622
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 402294 223954 402914 259398
rect 402294 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 402914 223954
rect 402294 223634 402914 223718
rect 402294 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 402914 223634
rect 402294 187954 402914 223398
rect 402294 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 402914 187954
rect 402294 187634 402914 187718
rect 402294 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 402914 187634
rect 402294 151954 402914 187398
rect 402294 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 402914 151954
rect 402294 151634 402914 151718
rect 402294 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 402914 151634
rect 402294 115954 402914 151398
rect 402294 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 402914 115954
rect 402294 115634 402914 115718
rect 402294 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 402914 115634
rect 402294 79954 402914 115398
rect 402294 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 402914 79954
rect 402294 79634 402914 79718
rect 402294 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 402914 79634
rect 402294 43954 402914 79398
rect 402294 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 402914 43954
rect 402294 43634 402914 43718
rect 402294 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 402914 43634
rect 402294 7954 402914 43398
rect 402294 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 402914 7954
rect 402294 7634 402914 7718
rect 402294 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 402914 7634
rect 402294 -1306 402914 7398
rect 402294 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 402914 -1306
rect 402294 -1626 402914 -1542
rect 402294 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 402914 -1626
rect 402294 -7654 402914 -1862
rect 406794 706758 407414 711590
rect 406794 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 407414 706758
rect 406794 706438 407414 706522
rect 406794 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 407414 706438
rect 406794 696454 407414 706202
rect 406794 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 407414 696454
rect 406794 696134 407414 696218
rect 406794 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 407414 696134
rect 406794 660454 407414 695898
rect 406794 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 407414 660454
rect 406794 660134 407414 660218
rect 406794 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 407414 660134
rect 406794 624454 407414 659898
rect 406794 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 407414 624454
rect 406794 624134 407414 624218
rect 406794 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 407414 624134
rect 406794 588454 407414 623898
rect 406794 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 407414 588454
rect 406794 588134 407414 588218
rect 406794 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 407414 588134
rect 406794 552454 407414 587898
rect 406794 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 407414 552454
rect 406794 552134 407414 552218
rect 406794 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 407414 552134
rect 406794 516454 407414 551898
rect 406794 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 407414 516454
rect 406794 516134 407414 516218
rect 406794 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 407414 516134
rect 406794 480454 407414 515898
rect 406794 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 407414 480454
rect 406794 480134 407414 480218
rect 406794 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 407414 480134
rect 406794 444454 407414 479898
rect 406794 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 407414 444454
rect 406794 444134 407414 444218
rect 406794 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 407414 444134
rect 406794 408454 407414 443898
rect 406794 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 407414 408454
rect 406794 408134 407414 408218
rect 406794 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 407414 408134
rect 406794 372454 407414 407898
rect 406794 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 407414 372454
rect 406794 372134 407414 372218
rect 406794 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 407414 372134
rect 406794 336454 407414 371898
rect 406794 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 407414 336454
rect 406794 336134 407414 336218
rect 406794 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 407414 336134
rect 406794 300454 407414 335898
rect 406794 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 407414 300454
rect 406794 300134 407414 300218
rect 406794 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 407414 300134
rect 406794 264454 407414 299898
rect 406794 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 407414 264454
rect 406794 264134 407414 264218
rect 406794 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 407414 264134
rect 406794 228454 407414 263898
rect 406794 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 407414 228454
rect 406794 228134 407414 228218
rect 406794 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 407414 228134
rect 406794 192454 407414 227898
rect 406794 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 407414 192454
rect 406794 192134 407414 192218
rect 406794 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 407414 192134
rect 406794 156454 407414 191898
rect 406794 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 407414 156454
rect 406794 156134 407414 156218
rect 406794 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 407414 156134
rect 406794 120454 407414 155898
rect 406794 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 407414 120454
rect 406794 120134 407414 120218
rect 406794 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 407414 120134
rect 406794 84454 407414 119898
rect 406794 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 407414 84454
rect 406794 84134 407414 84218
rect 406794 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 407414 84134
rect 406794 48454 407414 83898
rect 406794 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 407414 48454
rect 406794 48134 407414 48218
rect 406794 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 407414 48134
rect 406794 12454 407414 47898
rect 406794 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 407414 12454
rect 406794 12134 407414 12218
rect 406794 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 407414 12134
rect 406794 -2266 407414 11898
rect 406794 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 407414 -2266
rect 406794 -2586 407414 -2502
rect 406794 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 407414 -2586
rect 406794 -7654 407414 -2822
rect 411294 707718 411914 711590
rect 411294 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 411914 707718
rect 411294 707398 411914 707482
rect 411294 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 411914 707398
rect 411294 700954 411914 707162
rect 411294 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 411914 700954
rect 411294 700634 411914 700718
rect 411294 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 411914 700634
rect 411294 664954 411914 700398
rect 411294 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 411914 664954
rect 411294 664634 411914 664718
rect 411294 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 411914 664634
rect 411294 628954 411914 664398
rect 411294 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 411914 628954
rect 411294 628634 411914 628718
rect 411294 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 411914 628634
rect 411294 592954 411914 628398
rect 411294 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 411914 592954
rect 411294 592634 411914 592718
rect 411294 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 411914 592634
rect 411294 556954 411914 592398
rect 411294 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 411914 556954
rect 411294 556634 411914 556718
rect 411294 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 411914 556634
rect 411294 520954 411914 556398
rect 411294 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 411914 520954
rect 411294 520634 411914 520718
rect 411294 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 411914 520634
rect 411294 484954 411914 520398
rect 411294 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 411914 484954
rect 411294 484634 411914 484718
rect 411294 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 411914 484634
rect 411294 448954 411914 484398
rect 411294 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 411914 448954
rect 411294 448634 411914 448718
rect 411294 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 411914 448634
rect 411294 412954 411914 448398
rect 411294 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 411914 412954
rect 411294 412634 411914 412718
rect 411294 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 411914 412634
rect 411294 376954 411914 412398
rect 411294 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 411914 376954
rect 411294 376634 411914 376718
rect 411294 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 411914 376634
rect 411294 340954 411914 376398
rect 411294 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 411914 340954
rect 411294 340634 411914 340718
rect 411294 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 411914 340634
rect 411294 304954 411914 340398
rect 411294 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 411914 304954
rect 411294 304634 411914 304718
rect 411294 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 411914 304634
rect 411294 268954 411914 304398
rect 411294 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 411914 268954
rect 411294 268634 411914 268718
rect 411294 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 411914 268634
rect 411294 232954 411914 268398
rect 411294 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 411914 232954
rect 411294 232634 411914 232718
rect 411294 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 411914 232634
rect 411294 196954 411914 232398
rect 411294 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 411914 196954
rect 411294 196634 411914 196718
rect 411294 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 411914 196634
rect 411294 160954 411914 196398
rect 411294 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 411914 160954
rect 411294 160634 411914 160718
rect 411294 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 411914 160634
rect 411294 124954 411914 160398
rect 411294 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 411914 124954
rect 411294 124634 411914 124718
rect 411294 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 411914 124634
rect 411294 88954 411914 124398
rect 411294 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 411914 88954
rect 411294 88634 411914 88718
rect 411294 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 411914 88634
rect 411294 52954 411914 88398
rect 411294 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 411914 52954
rect 411294 52634 411914 52718
rect 411294 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 411914 52634
rect 411294 16954 411914 52398
rect 411294 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 411914 16954
rect 411294 16634 411914 16718
rect 411294 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 411914 16634
rect 411294 -3226 411914 16398
rect 411294 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 411914 -3226
rect 411294 -3546 411914 -3462
rect 411294 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 411914 -3546
rect 411294 -7654 411914 -3782
rect 415794 708678 416414 711590
rect 415794 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 416414 708678
rect 415794 708358 416414 708442
rect 415794 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 416414 708358
rect 415794 669454 416414 708122
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -4186 416414 20898
rect 415794 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 416414 -4186
rect 415794 -4506 416414 -4422
rect 415794 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 416414 -4506
rect 415794 -7654 416414 -4742
rect 420294 709638 420914 711590
rect 420294 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 420914 709638
rect 420294 709318 420914 709402
rect 420294 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 420914 709318
rect 420294 673954 420914 709082
rect 420294 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 420914 673954
rect 420294 673634 420914 673718
rect 420294 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 420914 673634
rect 420294 637954 420914 673398
rect 420294 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 420914 637954
rect 420294 637634 420914 637718
rect 420294 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 420914 637634
rect 420294 601954 420914 637398
rect 420294 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 420914 601954
rect 420294 601634 420914 601718
rect 420294 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 420914 601634
rect 420294 565954 420914 601398
rect 420294 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 420914 565954
rect 420294 565634 420914 565718
rect 420294 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 420914 565634
rect 420294 529954 420914 565398
rect 420294 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 420914 529954
rect 420294 529634 420914 529718
rect 420294 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 420914 529634
rect 420294 493954 420914 529398
rect 420294 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 420914 493954
rect 420294 493634 420914 493718
rect 420294 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 420914 493634
rect 420294 457954 420914 493398
rect 420294 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 420914 457954
rect 420294 457634 420914 457718
rect 420294 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 420914 457634
rect 420294 421954 420914 457398
rect 420294 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 420914 421954
rect 420294 421634 420914 421718
rect 420294 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 420914 421634
rect 420294 385954 420914 421398
rect 420294 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 420914 385954
rect 420294 385634 420914 385718
rect 420294 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 420914 385634
rect 420294 349954 420914 385398
rect 420294 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 420914 349954
rect 420294 349634 420914 349718
rect 420294 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 420914 349634
rect 420294 313954 420914 349398
rect 420294 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 420914 313954
rect 420294 313634 420914 313718
rect 420294 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 420914 313634
rect 420294 277954 420914 313398
rect 420294 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 420914 277954
rect 420294 277634 420914 277718
rect 420294 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 420914 277634
rect 420294 241954 420914 277398
rect 420294 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 420914 241954
rect 420294 241634 420914 241718
rect 420294 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 420914 241634
rect 420294 205954 420914 241398
rect 420294 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 420914 205954
rect 420294 205634 420914 205718
rect 420294 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 420914 205634
rect 420294 169954 420914 205398
rect 420294 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 420914 169954
rect 420294 169634 420914 169718
rect 420294 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 420914 169634
rect 420294 133954 420914 169398
rect 420294 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 420914 133954
rect 420294 133634 420914 133718
rect 420294 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 420914 133634
rect 420294 97954 420914 133398
rect 420294 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 420914 97954
rect 420294 97634 420914 97718
rect 420294 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 420914 97634
rect 420294 61954 420914 97398
rect 420294 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 420914 61954
rect 420294 61634 420914 61718
rect 420294 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 420914 61634
rect 420294 25954 420914 61398
rect 420294 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 420914 25954
rect 420294 25634 420914 25718
rect 420294 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 420914 25634
rect 420294 -5146 420914 25398
rect 420294 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 420914 -5146
rect 420294 -5466 420914 -5382
rect 420294 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 420914 -5466
rect 420294 -7654 420914 -5702
rect 424794 710598 425414 711590
rect 424794 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 425414 710598
rect 424794 710278 425414 710362
rect 424794 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 425414 710278
rect 424794 678454 425414 710042
rect 424794 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 425414 678454
rect 424794 678134 425414 678218
rect 424794 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 425414 678134
rect 424794 642454 425414 677898
rect 424794 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 425414 642454
rect 424794 642134 425414 642218
rect 424794 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 425414 642134
rect 424794 606454 425414 641898
rect 424794 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 425414 606454
rect 424794 606134 425414 606218
rect 424794 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 425414 606134
rect 424794 570454 425414 605898
rect 424794 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 425414 570454
rect 424794 570134 425414 570218
rect 424794 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 425414 570134
rect 424794 534454 425414 569898
rect 424794 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 425414 534454
rect 424794 534134 425414 534218
rect 424794 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 425414 534134
rect 424794 498454 425414 533898
rect 424794 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 425414 498454
rect 424794 498134 425414 498218
rect 424794 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 425414 498134
rect 424794 462454 425414 497898
rect 424794 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 425414 462454
rect 424794 462134 425414 462218
rect 424794 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 425414 462134
rect 424794 426454 425414 461898
rect 424794 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 425414 426454
rect 424794 426134 425414 426218
rect 424794 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 425414 426134
rect 424794 390454 425414 425898
rect 424794 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 425414 390454
rect 424794 390134 425414 390218
rect 424794 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 425414 390134
rect 424794 354454 425414 389898
rect 424794 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 425414 354454
rect 424794 354134 425414 354218
rect 424794 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 425414 354134
rect 424794 318454 425414 353898
rect 424794 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 425414 318454
rect 424794 318134 425414 318218
rect 424794 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 425414 318134
rect 424794 282454 425414 317898
rect 424794 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 425414 282454
rect 424794 282134 425414 282218
rect 424794 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 425414 282134
rect 424794 246454 425414 281898
rect 424794 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 425414 246454
rect 424794 246134 425414 246218
rect 424794 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 425414 246134
rect 424794 210454 425414 245898
rect 424794 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 425414 210454
rect 424794 210134 425414 210218
rect 424794 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 425414 210134
rect 424794 174454 425414 209898
rect 424794 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 425414 174454
rect 424794 174134 425414 174218
rect 424794 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 425414 174134
rect 424794 138454 425414 173898
rect 424794 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 425414 138454
rect 424794 138134 425414 138218
rect 424794 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 425414 138134
rect 424794 102454 425414 137898
rect 424794 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 425414 102454
rect 424794 102134 425414 102218
rect 424794 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 425414 102134
rect 424794 66454 425414 101898
rect 424794 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 425414 66454
rect 424794 66134 425414 66218
rect 424794 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 425414 66134
rect 424794 30454 425414 65898
rect 424794 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 425414 30454
rect 424794 30134 425414 30218
rect 424794 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 425414 30134
rect 424794 -6106 425414 29898
rect 424794 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 425414 -6106
rect 424794 -6426 425414 -6342
rect 424794 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 425414 -6426
rect 424794 -7654 425414 -6662
rect 429294 711558 429914 711590
rect 429294 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 429914 711558
rect 429294 711238 429914 711322
rect 429294 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 429914 711238
rect 429294 682954 429914 711002
rect 429294 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 429914 682954
rect 429294 682634 429914 682718
rect 429294 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 429914 682634
rect 429294 646954 429914 682398
rect 429294 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 429914 646954
rect 429294 646634 429914 646718
rect 429294 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 429914 646634
rect 429294 610954 429914 646398
rect 429294 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 429914 610954
rect 429294 610634 429914 610718
rect 429294 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 429914 610634
rect 429294 574954 429914 610398
rect 429294 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 429914 574954
rect 429294 574634 429914 574718
rect 429294 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 429914 574634
rect 429294 538954 429914 574398
rect 429294 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 429914 538954
rect 429294 538634 429914 538718
rect 429294 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 429914 538634
rect 429294 502954 429914 538398
rect 429294 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 429914 502954
rect 429294 502634 429914 502718
rect 429294 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 429914 502634
rect 429294 466954 429914 502398
rect 429294 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 429914 466954
rect 429294 466634 429914 466718
rect 429294 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 429914 466634
rect 429294 430954 429914 466398
rect 429294 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 429914 430954
rect 429294 430634 429914 430718
rect 429294 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 429914 430634
rect 429294 394954 429914 430398
rect 429294 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 429914 394954
rect 429294 394634 429914 394718
rect 429294 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 429914 394634
rect 429294 358954 429914 394398
rect 429294 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 429914 358954
rect 429294 358634 429914 358718
rect 429294 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 429914 358634
rect 429294 322954 429914 358398
rect 429294 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 429914 322954
rect 429294 322634 429914 322718
rect 429294 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 429914 322634
rect 429294 286954 429914 322398
rect 429294 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 429914 286954
rect 429294 286634 429914 286718
rect 429294 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 429914 286634
rect 429294 250954 429914 286398
rect 429294 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 429914 250954
rect 429294 250634 429914 250718
rect 429294 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 429914 250634
rect 429294 214954 429914 250398
rect 429294 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 429914 214954
rect 429294 214634 429914 214718
rect 429294 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 429914 214634
rect 429294 178954 429914 214398
rect 429294 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 429914 178954
rect 429294 178634 429914 178718
rect 429294 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 429914 178634
rect 429294 142954 429914 178398
rect 429294 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 429914 142954
rect 429294 142634 429914 142718
rect 429294 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 429914 142634
rect 429294 106954 429914 142398
rect 429294 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 429914 106954
rect 429294 106634 429914 106718
rect 429294 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 429914 106634
rect 429294 70954 429914 106398
rect 429294 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 429914 70954
rect 429294 70634 429914 70718
rect 429294 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 429914 70634
rect 429294 34954 429914 70398
rect 429294 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 429914 34954
rect 429294 34634 429914 34718
rect 429294 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 429914 34634
rect 429294 -7066 429914 34398
rect 429294 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 429914 -7066
rect 429294 -7386 429914 -7302
rect 429294 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 429914 -7386
rect 429294 -7654 429914 -7622
rect 433794 704838 434414 711590
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 438294 705798 438914 711590
rect 438294 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 438914 705798
rect 438294 705478 438914 705562
rect 438294 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 438914 705478
rect 438294 691954 438914 705242
rect 438294 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 438914 691954
rect 438294 691634 438914 691718
rect 438294 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 438914 691634
rect 438294 655954 438914 691398
rect 438294 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 438914 655954
rect 438294 655634 438914 655718
rect 438294 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 438914 655634
rect 438294 619954 438914 655398
rect 438294 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 438914 619954
rect 438294 619634 438914 619718
rect 438294 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 438914 619634
rect 438294 583954 438914 619398
rect 438294 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 438914 583954
rect 438294 583634 438914 583718
rect 438294 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 438914 583634
rect 438294 547954 438914 583398
rect 438294 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 438914 547954
rect 438294 547634 438914 547718
rect 438294 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 438914 547634
rect 438294 511954 438914 547398
rect 438294 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 438914 511954
rect 438294 511634 438914 511718
rect 438294 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 438914 511634
rect 438294 475954 438914 511398
rect 438294 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 438914 475954
rect 438294 475634 438914 475718
rect 438294 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 438914 475634
rect 438294 439954 438914 475398
rect 438294 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 438914 439954
rect 438294 439634 438914 439718
rect 438294 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 438914 439634
rect 438294 403954 438914 439398
rect 438294 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 438914 403954
rect 438294 403634 438914 403718
rect 438294 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 438914 403634
rect 438294 367954 438914 403398
rect 438294 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 438914 367954
rect 438294 367634 438914 367718
rect 438294 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 438914 367634
rect 438294 331954 438914 367398
rect 438294 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 438914 331954
rect 438294 331634 438914 331718
rect 438294 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 438914 331634
rect 438294 295954 438914 331398
rect 438294 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 438914 295954
rect 438294 295634 438914 295718
rect 438294 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 438914 295634
rect 438294 259954 438914 295398
rect 438294 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 438914 259954
rect 438294 259634 438914 259718
rect 438294 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 438914 259634
rect 438294 223954 438914 259398
rect 438294 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 438914 223954
rect 438294 223634 438914 223718
rect 438294 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 438914 223634
rect 438294 187954 438914 223398
rect 438294 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 438914 187954
rect 438294 187634 438914 187718
rect 438294 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 438914 187634
rect 438294 151954 438914 187398
rect 438294 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 438914 151954
rect 438294 151634 438914 151718
rect 438294 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 438914 151634
rect 438294 115954 438914 151398
rect 438294 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 438914 115954
rect 438294 115634 438914 115718
rect 438294 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 438914 115634
rect 438294 79954 438914 115398
rect 438294 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 438914 79954
rect 438294 79634 438914 79718
rect 438294 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 438914 79634
rect 438294 43954 438914 79398
rect 438294 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 438914 43954
rect 438294 43634 438914 43718
rect 438294 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 438914 43634
rect 438294 7954 438914 43398
rect 438294 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 438914 7954
rect 438294 7634 438914 7718
rect 438294 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 438914 7634
rect 438294 -1306 438914 7398
rect 438294 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 438914 -1306
rect 438294 -1626 438914 -1542
rect 438294 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 438914 -1626
rect 438294 -7654 438914 -1862
rect 442794 706758 443414 711590
rect 442794 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 443414 706758
rect 442794 706438 443414 706522
rect 442794 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 443414 706438
rect 442794 696454 443414 706202
rect 442794 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 443414 696454
rect 442794 696134 443414 696218
rect 442794 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 443414 696134
rect 442794 660454 443414 695898
rect 442794 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 443414 660454
rect 442794 660134 443414 660218
rect 442794 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 443414 660134
rect 442794 624454 443414 659898
rect 442794 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 443414 624454
rect 442794 624134 443414 624218
rect 442794 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 443414 624134
rect 442794 588454 443414 623898
rect 442794 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 443414 588454
rect 442794 588134 443414 588218
rect 442794 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 443414 588134
rect 442794 552454 443414 587898
rect 442794 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 443414 552454
rect 442794 552134 443414 552218
rect 442794 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 443414 552134
rect 442794 516454 443414 551898
rect 442794 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 443414 516454
rect 442794 516134 443414 516218
rect 442794 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 443414 516134
rect 442794 480454 443414 515898
rect 442794 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 443414 480454
rect 442794 480134 443414 480218
rect 442794 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 443414 480134
rect 442794 444454 443414 479898
rect 442794 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 443414 444454
rect 442794 444134 443414 444218
rect 442794 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 443414 444134
rect 442794 408454 443414 443898
rect 442794 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 443414 408454
rect 442794 408134 443414 408218
rect 442794 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 443414 408134
rect 442794 372454 443414 407898
rect 442794 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 443414 372454
rect 442794 372134 443414 372218
rect 442794 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 443414 372134
rect 442794 336454 443414 371898
rect 442794 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 443414 336454
rect 442794 336134 443414 336218
rect 442794 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 443414 336134
rect 442794 300454 443414 335898
rect 442794 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 443414 300454
rect 442794 300134 443414 300218
rect 442794 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 443414 300134
rect 442794 264454 443414 299898
rect 442794 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 443414 264454
rect 442794 264134 443414 264218
rect 442794 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 443414 264134
rect 442794 228454 443414 263898
rect 442794 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 443414 228454
rect 442794 228134 443414 228218
rect 442794 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 443414 228134
rect 442794 192454 443414 227898
rect 442794 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 443414 192454
rect 442794 192134 443414 192218
rect 442794 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 443414 192134
rect 442794 156454 443414 191898
rect 442794 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 443414 156454
rect 442794 156134 443414 156218
rect 442794 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 443414 156134
rect 442794 120454 443414 155898
rect 442794 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 443414 120454
rect 442794 120134 443414 120218
rect 442794 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 443414 120134
rect 442794 84454 443414 119898
rect 442794 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 443414 84454
rect 442794 84134 443414 84218
rect 442794 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 443414 84134
rect 442794 48454 443414 83898
rect 442794 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 443414 48454
rect 442794 48134 443414 48218
rect 442794 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 443414 48134
rect 442794 12454 443414 47898
rect 442794 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 443414 12454
rect 442794 12134 443414 12218
rect 442794 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 443414 12134
rect 442794 -2266 443414 11898
rect 442794 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 443414 -2266
rect 442794 -2586 443414 -2502
rect 442794 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 443414 -2586
rect 442794 -7654 443414 -2822
rect 447294 707718 447914 711590
rect 447294 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 447914 707718
rect 447294 707398 447914 707482
rect 447294 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 447914 707398
rect 447294 700954 447914 707162
rect 447294 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 447914 700954
rect 447294 700634 447914 700718
rect 447294 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 447914 700634
rect 447294 664954 447914 700398
rect 447294 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 447914 664954
rect 447294 664634 447914 664718
rect 447294 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 447914 664634
rect 447294 628954 447914 664398
rect 447294 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 447914 628954
rect 447294 628634 447914 628718
rect 447294 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 447914 628634
rect 447294 592954 447914 628398
rect 447294 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 447914 592954
rect 447294 592634 447914 592718
rect 447294 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 447914 592634
rect 447294 556954 447914 592398
rect 447294 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 447914 556954
rect 447294 556634 447914 556718
rect 447294 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 447914 556634
rect 447294 520954 447914 556398
rect 447294 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 447914 520954
rect 447294 520634 447914 520718
rect 447294 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 447914 520634
rect 447294 484954 447914 520398
rect 447294 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 447914 484954
rect 447294 484634 447914 484718
rect 447294 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 447914 484634
rect 447294 448954 447914 484398
rect 447294 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 447914 448954
rect 447294 448634 447914 448718
rect 447294 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 447914 448634
rect 447294 412954 447914 448398
rect 447294 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 447914 412954
rect 447294 412634 447914 412718
rect 447294 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 447914 412634
rect 447294 376954 447914 412398
rect 447294 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 447914 376954
rect 447294 376634 447914 376718
rect 447294 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 447914 376634
rect 447294 340954 447914 376398
rect 447294 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 447914 340954
rect 447294 340634 447914 340718
rect 447294 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 447914 340634
rect 447294 304954 447914 340398
rect 447294 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 447914 304954
rect 447294 304634 447914 304718
rect 447294 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 447914 304634
rect 447294 268954 447914 304398
rect 447294 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 447914 268954
rect 447294 268634 447914 268718
rect 447294 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 447914 268634
rect 447294 232954 447914 268398
rect 447294 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 447914 232954
rect 447294 232634 447914 232718
rect 447294 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 447914 232634
rect 447294 196954 447914 232398
rect 447294 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 447914 196954
rect 447294 196634 447914 196718
rect 447294 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 447914 196634
rect 447294 160954 447914 196398
rect 447294 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 447914 160954
rect 447294 160634 447914 160718
rect 447294 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 447914 160634
rect 447294 124954 447914 160398
rect 447294 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 447914 124954
rect 447294 124634 447914 124718
rect 447294 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 447914 124634
rect 447294 88954 447914 124398
rect 447294 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 447914 88954
rect 447294 88634 447914 88718
rect 447294 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 447914 88634
rect 447294 52954 447914 88398
rect 447294 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 447914 52954
rect 447294 52634 447914 52718
rect 447294 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 447914 52634
rect 447294 16954 447914 52398
rect 447294 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 447914 16954
rect 447294 16634 447914 16718
rect 447294 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 447914 16634
rect 447294 -3226 447914 16398
rect 447294 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 447914 -3226
rect 447294 -3546 447914 -3462
rect 447294 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 447914 -3546
rect 447294 -7654 447914 -3782
rect 451794 708678 452414 711590
rect 451794 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 452414 708678
rect 451794 708358 452414 708442
rect 451794 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 452414 708358
rect 451794 669454 452414 708122
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -4186 452414 20898
rect 451794 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 452414 -4186
rect 451794 -4506 452414 -4422
rect 451794 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 452414 -4506
rect 451794 -7654 452414 -4742
rect 456294 709638 456914 711590
rect 456294 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 456914 709638
rect 456294 709318 456914 709402
rect 456294 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 456914 709318
rect 456294 673954 456914 709082
rect 456294 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 456914 673954
rect 456294 673634 456914 673718
rect 456294 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 456914 673634
rect 456294 637954 456914 673398
rect 456294 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 456914 637954
rect 456294 637634 456914 637718
rect 456294 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 456914 637634
rect 456294 601954 456914 637398
rect 456294 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 456914 601954
rect 456294 601634 456914 601718
rect 456294 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 456914 601634
rect 456294 565954 456914 601398
rect 456294 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 456914 565954
rect 456294 565634 456914 565718
rect 456294 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 456914 565634
rect 456294 529954 456914 565398
rect 456294 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 456914 529954
rect 456294 529634 456914 529718
rect 456294 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 456914 529634
rect 456294 493954 456914 529398
rect 456294 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 456914 493954
rect 456294 493634 456914 493718
rect 456294 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 456914 493634
rect 456294 457954 456914 493398
rect 456294 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 456914 457954
rect 456294 457634 456914 457718
rect 456294 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 456914 457634
rect 456294 421954 456914 457398
rect 456294 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 456914 421954
rect 456294 421634 456914 421718
rect 456294 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 456914 421634
rect 456294 385954 456914 421398
rect 456294 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 456914 385954
rect 456294 385634 456914 385718
rect 456294 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 456914 385634
rect 456294 349954 456914 385398
rect 456294 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 456914 349954
rect 456294 349634 456914 349718
rect 456294 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 456914 349634
rect 456294 313954 456914 349398
rect 456294 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 456914 313954
rect 456294 313634 456914 313718
rect 456294 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 456914 313634
rect 456294 277954 456914 313398
rect 456294 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 456914 277954
rect 456294 277634 456914 277718
rect 456294 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 456914 277634
rect 456294 241954 456914 277398
rect 456294 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 456914 241954
rect 456294 241634 456914 241718
rect 456294 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 456914 241634
rect 456294 205954 456914 241398
rect 456294 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 456914 205954
rect 456294 205634 456914 205718
rect 456294 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 456914 205634
rect 456294 169954 456914 205398
rect 456294 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 456914 169954
rect 456294 169634 456914 169718
rect 456294 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 456914 169634
rect 456294 133954 456914 169398
rect 456294 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 456914 133954
rect 456294 133634 456914 133718
rect 456294 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 456914 133634
rect 456294 97954 456914 133398
rect 456294 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 456914 97954
rect 456294 97634 456914 97718
rect 456294 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 456914 97634
rect 456294 61954 456914 97398
rect 456294 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 456914 61954
rect 456294 61634 456914 61718
rect 456294 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 456914 61634
rect 456294 25954 456914 61398
rect 456294 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 456914 25954
rect 456294 25634 456914 25718
rect 456294 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 456914 25634
rect 456294 -5146 456914 25398
rect 456294 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 456914 -5146
rect 456294 -5466 456914 -5382
rect 456294 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 456914 -5466
rect 456294 -7654 456914 -5702
rect 460794 710598 461414 711590
rect 460794 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 461414 710598
rect 460794 710278 461414 710362
rect 460794 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 461414 710278
rect 460794 678454 461414 710042
rect 460794 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 461414 678454
rect 460794 678134 461414 678218
rect 460794 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 461414 678134
rect 460794 642454 461414 677898
rect 460794 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 461414 642454
rect 460794 642134 461414 642218
rect 460794 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 461414 642134
rect 460794 606454 461414 641898
rect 460794 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 461414 606454
rect 460794 606134 461414 606218
rect 460794 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 461414 606134
rect 460794 570454 461414 605898
rect 460794 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 461414 570454
rect 460794 570134 461414 570218
rect 460794 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 461414 570134
rect 460794 534454 461414 569898
rect 460794 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 461414 534454
rect 460794 534134 461414 534218
rect 460794 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 461414 534134
rect 460794 498454 461414 533898
rect 460794 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 461414 498454
rect 460794 498134 461414 498218
rect 460794 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 461414 498134
rect 460794 462454 461414 497898
rect 460794 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 461414 462454
rect 460794 462134 461414 462218
rect 460794 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 461414 462134
rect 460794 426454 461414 461898
rect 460794 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 461414 426454
rect 460794 426134 461414 426218
rect 460794 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 461414 426134
rect 460794 390454 461414 425898
rect 460794 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 461414 390454
rect 460794 390134 461414 390218
rect 460794 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 461414 390134
rect 460794 354454 461414 389898
rect 460794 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 461414 354454
rect 460794 354134 461414 354218
rect 460794 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 461414 354134
rect 460794 318454 461414 353898
rect 460794 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 461414 318454
rect 460794 318134 461414 318218
rect 460794 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 461414 318134
rect 460794 282454 461414 317898
rect 460794 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 461414 282454
rect 460794 282134 461414 282218
rect 460794 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 461414 282134
rect 460794 246454 461414 281898
rect 460794 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 461414 246454
rect 460794 246134 461414 246218
rect 460794 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 461414 246134
rect 460794 210454 461414 245898
rect 460794 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 461414 210454
rect 460794 210134 461414 210218
rect 460794 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 461414 210134
rect 460794 174454 461414 209898
rect 460794 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 461414 174454
rect 460794 174134 461414 174218
rect 460794 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 461414 174134
rect 460794 138454 461414 173898
rect 460794 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 461414 138454
rect 460794 138134 461414 138218
rect 460794 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 461414 138134
rect 460794 102454 461414 137898
rect 460794 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 461414 102454
rect 460794 102134 461414 102218
rect 460794 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 461414 102134
rect 460794 66454 461414 101898
rect 460794 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 461414 66454
rect 460794 66134 461414 66218
rect 460794 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 461414 66134
rect 460794 30454 461414 65898
rect 460794 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 461414 30454
rect 460794 30134 461414 30218
rect 460794 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 461414 30134
rect 460794 -6106 461414 29898
rect 460794 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 461414 -6106
rect 460794 -6426 461414 -6342
rect 460794 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 461414 -6426
rect 460794 -7654 461414 -6662
rect 465294 711558 465914 711590
rect 465294 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 465914 711558
rect 465294 711238 465914 711322
rect 465294 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 465914 711238
rect 465294 682954 465914 711002
rect 465294 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 465914 682954
rect 465294 682634 465914 682718
rect 465294 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 465914 682634
rect 465294 646954 465914 682398
rect 465294 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 465914 646954
rect 465294 646634 465914 646718
rect 465294 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 465914 646634
rect 465294 610954 465914 646398
rect 465294 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 465914 610954
rect 465294 610634 465914 610718
rect 465294 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 465914 610634
rect 465294 574954 465914 610398
rect 465294 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 465914 574954
rect 465294 574634 465914 574718
rect 465294 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 465914 574634
rect 465294 538954 465914 574398
rect 465294 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 465914 538954
rect 465294 538634 465914 538718
rect 465294 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 465914 538634
rect 465294 502954 465914 538398
rect 465294 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 465914 502954
rect 465294 502634 465914 502718
rect 465294 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 465914 502634
rect 465294 466954 465914 502398
rect 465294 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 465914 466954
rect 465294 466634 465914 466718
rect 465294 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 465914 466634
rect 465294 430954 465914 466398
rect 465294 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 465914 430954
rect 465294 430634 465914 430718
rect 465294 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 465914 430634
rect 465294 394954 465914 430398
rect 465294 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 465914 394954
rect 465294 394634 465914 394718
rect 465294 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 465914 394634
rect 465294 358954 465914 394398
rect 465294 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 465914 358954
rect 465294 358634 465914 358718
rect 465294 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 465914 358634
rect 465294 322954 465914 358398
rect 465294 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 465914 322954
rect 465294 322634 465914 322718
rect 465294 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 465914 322634
rect 465294 286954 465914 322398
rect 465294 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 465914 286954
rect 465294 286634 465914 286718
rect 465294 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 465914 286634
rect 465294 250954 465914 286398
rect 465294 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 465914 250954
rect 465294 250634 465914 250718
rect 465294 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 465914 250634
rect 465294 214954 465914 250398
rect 465294 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 465914 214954
rect 465294 214634 465914 214718
rect 465294 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 465914 214634
rect 465294 178954 465914 214398
rect 465294 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 465914 178954
rect 465294 178634 465914 178718
rect 465294 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 465914 178634
rect 465294 142954 465914 178398
rect 465294 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 465914 142954
rect 465294 142634 465914 142718
rect 465294 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 465914 142634
rect 465294 106954 465914 142398
rect 465294 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 465914 106954
rect 465294 106634 465914 106718
rect 465294 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 465914 106634
rect 465294 70954 465914 106398
rect 465294 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 465914 70954
rect 465294 70634 465914 70718
rect 465294 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 465914 70634
rect 465294 34954 465914 70398
rect 465294 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 465914 34954
rect 465294 34634 465914 34718
rect 465294 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 465914 34634
rect 465294 -7066 465914 34398
rect 465294 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 465914 -7066
rect 465294 -7386 465914 -7302
rect 465294 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 465914 -7386
rect 465294 -7654 465914 -7622
rect 469794 704838 470414 711590
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 474294 705798 474914 711590
rect 474294 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 474914 705798
rect 474294 705478 474914 705562
rect 474294 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 474914 705478
rect 474294 691954 474914 705242
rect 474294 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 474914 691954
rect 474294 691634 474914 691718
rect 474294 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 474914 691634
rect 474294 655954 474914 691398
rect 474294 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 474914 655954
rect 474294 655634 474914 655718
rect 474294 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 474914 655634
rect 474294 619954 474914 655398
rect 474294 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 474914 619954
rect 474294 619634 474914 619718
rect 474294 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 474914 619634
rect 474294 583954 474914 619398
rect 474294 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 474914 583954
rect 474294 583634 474914 583718
rect 474294 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 474914 583634
rect 474294 547954 474914 583398
rect 474294 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 474914 547954
rect 474294 547634 474914 547718
rect 474294 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 474914 547634
rect 474294 511954 474914 547398
rect 474294 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 474914 511954
rect 474294 511634 474914 511718
rect 474294 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 474914 511634
rect 474294 475954 474914 511398
rect 474294 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 474914 475954
rect 474294 475634 474914 475718
rect 474294 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 474914 475634
rect 474294 439954 474914 475398
rect 474294 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 474914 439954
rect 474294 439634 474914 439718
rect 474294 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 474914 439634
rect 474294 403954 474914 439398
rect 474294 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 474914 403954
rect 474294 403634 474914 403718
rect 474294 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 474914 403634
rect 474294 367954 474914 403398
rect 474294 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 474914 367954
rect 474294 367634 474914 367718
rect 474294 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 474914 367634
rect 474294 331954 474914 367398
rect 474294 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 474914 331954
rect 474294 331634 474914 331718
rect 474294 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 474914 331634
rect 474294 295954 474914 331398
rect 474294 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 474914 295954
rect 474294 295634 474914 295718
rect 474294 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 474914 295634
rect 474294 259954 474914 295398
rect 474294 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 474914 259954
rect 474294 259634 474914 259718
rect 474294 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 474914 259634
rect 474294 223954 474914 259398
rect 474294 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 474914 223954
rect 474294 223634 474914 223718
rect 474294 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 474914 223634
rect 474294 187954 474914 223398
rect 474294 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 474914 187954
rect 474294 187634 474914 187718
rect 474294 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 474914 187634
rect 474294 151954 474914 187398
rect 474294 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 474914 151954
rect 474294 151634 474914 151718
rect 474294 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 474914 151634
rect 474294 115954 474914 151398
rect 474294 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 474914 115954
rect 474294 115634 474914 115718
rect 474294 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 474914 115634
rect 474294 79954 474914 115398
rect 474294 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 474914 79954
rect 474294 79634 474914 79718
rect 474294 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 474914 79634
rect 474294 43954 474914 79398
rect 474294 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 474914 43954
rect 474294 43634 474914 43718
rect 474294 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 474914 43634
rect 474294 7954 474914 43398
rect 474294 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 474914 7954
rect 474294 7634 474914 7718
rect 474294 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 474914 7634
rect 474294 -1306 474914 7398
rect 474294 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 474914 -1306
rect 474294 -1626 474914 -1542
rect 474294 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 474914 -1626
rect 474294 -7654 474914 -1862
rect 478794 706758 479414 711590
rect 478794 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 479414 706758
rect 478794 706438 479414 706522
rect 478794 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 479414 706438
rect 478794 696454 479414 706202
rect 478794 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 479414 696454
rect 478794 696134 479414 696218
rect 478794 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 479414 696134
rect 478794 660454 479414 695898
rect 478794 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 479414 660454
rect 478794 660134 479414 660218
rect 478794 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 479414 660134
rect 478794 624454 479414 659898
rect 478794 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 479414 624454
rect 478794 624134 479414 624218
rect 478794 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 479414 624134
rect 478794 588454 479414 623898
rect 478794 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 479414 588454
rect 478794 588134 479414 588218
rect 478794 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 479414 588134
rect 478794 552454 479414 587898
rect 478794 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 479414 552454
rect 478794 552134 479414 552218
rect 478794 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 479414 552134
rect 478794 516454 479414 551898
rect 478794 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 479414 516454
rect 478794 516134 479414 516218
rect 478794 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 479414 516134
rect 478794 480454 479414 515898
rect 478794 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 479414 480454
rect 478794 480134 479414 480218
rect 478794 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 479414 480134
rect 478794 444454 479414 479898
rect 478794 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 479414 444454
rect 478794 444134 479414 444218
rect 478794 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 479414 444134
rect 478794 408454 479414 443898
rect 478794 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 479414 408454
rect 478794 408134 479414 408218
rect 478794 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 479414 408134
rect 478794 372454 479414 407898
rect 478794 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 479414 372454
rect 478794 372134 479414 372218
rect 478794 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 479414 372134
rect 478794 336454 479414 371898
rect 478794 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 479414 336454
rect 478794 336134 479414 336218
rect 478794 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 479414 336134
rect 478794 300454 479414 335898
rect 478794 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 479414 300454
rect 478794 300134 479414 300218
rect 478794 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 479414 300134
rect 478794 264454 479414 299898
rect 478794 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 479414 264454
rect 478794 264134 479414 264218
rect 478794 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 479414 264134
rect 478794 228454 479414 263898
rect 478794 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 479414 228454
rect 478794 228134 479414 228218
rect 478794 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 479414 228134
rect 478794 192454 479414 227898
rect 478794 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 479414 192454
rect 478794 192134 479414 192218
rect 478794 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 479414 192134
rect 478794 156454 479414 191898
rect 478794 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 479414 156454
rect 478794 156134 479414 156218
rect 478794 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 479414 156134
rect 478794 120454 479414 155898
rect 478794 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 479414 120454
rect 478794 120134 479414 120218
rect 478794 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 479414 120134
rect 478794 84454 479414 119898
rect 478794 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 479414 84454
rect 478794 84134 479414 84218
rect 478794 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 479414 84134
rect 478794 48454 479414 83898
rect 478794 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 479414 48454
rect 478794 48134 479414 48218
rect 478794 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 479414 48134
rect 478794 12454 479414 47898
rect 478794 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 479414 12454
rect 478794 12134 479414 12218
rect 478794 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 479414 12134
rect 478794 -2266 479414 11898
rect 478794 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 479414 -2266
rect 478794 -2586 479414 -2502
rect 478794 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 479414 -2586
rect 478794 -7654 479414 -2822
rect 483294 707718 483914 711590
rect 483294 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 483914 707718
rect 483294 707398 483914 707482
rect 483294 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 483914 707398
rect 483294 700954 483914 707162
rect 483294 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 483914 700954
rect 483294 700634 483914 700718
rect 483294 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 483914 700634
rect 483294 664954 483914 700398
rect 483294 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 483914 664954
rect 483294 664634 483914 664718
rect 483294 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 483914 664634
rect 483294 628954 483914 664398
rect 483294 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 483914 628954
rect 483294 628634 483914 628718
rect 483294 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 483914 628634
rect 483294 592954 483914 628398
rect 483294 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 483914 592954
rect 483294 592634 483914 592718
rect 483294 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 483914 592634
rect 483294 556954 483914 592398
rect 483294 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 483914 556954
rect 483294 556634 483914 556718
rect 483294 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 483914 556634
rect 483294 520954 483914 556398
rect 483294 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 483914 520954
rect 483294 520634 483914 520718
rect 483294 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 483914 520634
rect 483294 484954 483914 520398
rect 483294 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 483914 484954
rect 483294 484634 483914 484718
rect 483294 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 483914 484634
rect 483294 448954 483914 484398
rect 483294 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 483914 448954
rect 483294 448634 483914 448718
rect 483294 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 483914 448634
rect 483294 412954 483914 448398
rect 483294 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 483914 412954
rect 483294 412634 483914 412718
rect 483294 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 483914 412634
rect 483294 376954 483914 412398
rect 483294 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 483914 376954
rect 483294 376634 483914 376718
rect 483294 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 483914 376634
rect 483294 340954 483914 376398
rect 483294 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 483914 340954
rect 483294 340634 483914 340718
rect 483294 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 483914 340634
rect 483294 304954 483914 340398
rect 483294 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 483914 304954
rect 483294 304634 483914 304718
rect 483294 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 483914 304634
rect 483294 268954 483914 304398
rect 483294 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 483914 268954
rect 483294 268634 483914 268718
rect 483294 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 483914 268634
rect 483294 232954 483914 268398
rect 483294 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 483914 232954
rect 483294 232634 483914 232718
rect 483294 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 483914 232634
rect 483294 196954 483914 232398
rect 483294 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 483914 196954
rect 483294 196634 483914 196718
rect 483294 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 483914 196634
rect 483294 160954 483914 196398
rect 483294 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 483914 160954
rect 483294 160634 483914 160718
rect 483294 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 483914 160634
rect 483294 124954 483914 160398
rect 483294 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 483914 124954
rect 483294 124634 483914 124718
rect 483294 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 483914 124634
rect 483294 88954 483914 124398
rect 483294 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 483914 88954
rect 483294 88634 483914 88718
rect 483294 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 483914 88634
rect 483294 52954 483914 88398
rect 483294 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 483914 52954
rect 483294 52634 483914 52718
rect 483294 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 483914 52634
rect 483294 16954 483914 52398
rect 483294 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 483914 16954
rect 483294 16634 483914 16718
rect 483294 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 483914 16634
rect 483294 -3226 483914 16398
rect 483294 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 483914 -3226
rect 483294 -3546 483914 -3462
rect 483294 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 483914 -3546
rect 483294 -7654 483914 -3782
rect 487794 708678 488414 711590
rect 487794 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 488414 708678
rect 487794 708358 488414 708442
rect 487794 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 488414 708358
rect 487794 669454 488414 708122
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -4186 488414 20898
rect 487794 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 488414 -4186
rect 487794 -4506 488414 -4422
rect 487794 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 488414 -4506
rect 487794 -7654 488414 -4742
rect 492294 709638 492914 711590
rect 492294 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 492914 709638
rect 492294 709318 492914 709402
rect 492294 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 492914 709318
rect 492294 673954 492914 709082
rect 492294 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 492914 673954
rect 492294 673634 492914 673718
rect 492294 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 492914 673634
rect 492294 637954 492914 673398
rect 492294 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 492914 637954
rect 492294 637634 492914 637718
rect 492294 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 492914 637634
rect 492294 601954 492914 637398
rect 492294 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 492914 601954
rect 492294 601634 492914 601718
rect 492294 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 492914 601634
rect 492294 565954 492914 601398
rect 492294 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 492914 565954
rect 492294 565634 492914 565718
rect 492294 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 492914 565634
rect 492294 529954 492914 565398
rect 492294 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 492914 529954
rect 492294 529634 492914 529718
rect 492294 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 492914 529634
rect 492294 493954 492914 529398
rect 492294 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 492914 493954
rect 492294 493634 492914 493718
rect 492294 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 492914 493634
rect 492294 457954 492914 493398
rect 492294 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 492914 457954
rect 492294 457634 492914 457718
rect 492294 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 492914 457634
rect 492294 421954 492914 457398
rect 492294 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 492914 421954
rect 492294 421634 492914 421718
rect 492294 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 492914 421634
rect 492294 385954 492914 421398
rect 492294 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 492914 385954
rect 492294 385634 492914 385718
rect 492294 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 492914 385634
rect 492294 349954 492914 385398
rect 492294 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 492914 349954
rect 492294 349634 492914 349718
rect 492294 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 492914 349634
rect 492294 313954 492914 349398
rect 492294 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 492914 313954
rect 492294 313634 492914 313718
rect 492294 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 492914 313634
rect 492294 277954 492914 313398
rect 492294 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 492914 277954
rect 492294 277634 492914 277718
rect 492294 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 492914 277634
rect 492294 241954 492914 277398
rect 492294 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 492914 241954
rect 492294 241634 492914 241718
rect 492294 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 492914 241634
rect 492294 205954 492914 241398
rect 492294 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 492914 205954
rect 492294 205634 492914 205718
rect 492294 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 492914 205634
rect 492294 169954 492914 205398
rect 492294 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 492914 169954
rect 492294 169634 492914 169718
rect 492294 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 492914 169634
rect 492294 133954 492914 169398
rect 492294 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 492914 133954
rect 492294 133634 492914 133718
rect 492294 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 492914 133634
rect 492294 97954 492914 133398
rect 492294 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 492914 97954
rect 492294 97634 492914 97718
rect 492294 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 492914 97634
rect 492294 61954 492914 97398
rect 492294 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 492914 61954
rect 492294 61634 492914 61718
rect 492294 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 492914 61634
rect 492294 25954 492914 61398
rect 492294 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 492914 25954
rect 492294 25634 492914 25718
rect 492294 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 492914 25634
rect 492294 -5146 492914 25398
rect 492294 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 492914 -5146
rect 492294 -5466 492914 -5382
rect 492294 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 492914 -5466
rect 492294 -7654 492914 -5702
rect 496794 710598 497414 711590
rect 496794 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 497414 710598
rect 496794 710278 497414 710362
rect 496794 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 497414 710278
rect 496794 678454 497414 710042
rect 496794 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 497414 678454
rect 496794 678134 497414 678218
rect 496794 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 497414 678134
rect 496794 642454 497414 677898
rect 496794 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 497414 642454
rect 496794 642134 497414 642218
rect 496794 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 497414 642134
rect 496794 606454 497414 641898
rect 496794 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 497414 606454
rect 496794 606134 497414 606218
rect 496794 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 497414 606134
rect 496794 570454 497414 605898
rect 496794 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 497414 570454
rect 496794 570134 497414 570218
rect 496794 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 497414 570134
rect 496794 534454 497414 569898
rect 496794 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 497414 534454
rect 496794 534134 497414 534218
rect 496794 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 497414 534134
rect 496794 498454 497414 533898
rect 496794 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 497414 498454
rect 496794 498134 497414 498218
rect 496794 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 497414 498134
rect 496794 462454 497414 497898
rect 496794 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 497414 462454
rect 496794 462134 497414 462218
rect 496794 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 497414 462134
rect 496794 426454 497414 461898
rect 496794 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 497414 426454
rect 496794 426134 497414 426218
rect 496794 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 497414 426134
rect 496794 390454 497414 425898
rect 496794 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 497414 390454
rect 496794 390134 497414 390218
rect 496794 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 497414 390134
rect 496794 354454 497414 389898
rect 496794 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 497414 354454
rect 496794 354134 497414 354218
rect 496794 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 497414 354134
rect 496794 318454 497414 353898
rect 496794 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 497414 318454
rect 496794 318134 497414 318218
rect 496794 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 497414 318134
rect 496794 282454 497414 317898
rect 496794 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 497414 282454
rect 496794 282134 497414 282218
rect 496794 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 497414 282134
rect 496794 246454 497414 281898
rect 496794 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 497414 246454
rect 496794 246134 497414 246218
rect 496794 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 497414 246134
rect 496794 210454 497414 245898
rect 496794 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 497414 210454
rect 496794 210134 497414 210218
rect 496794 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 497414 210134
rect 496794 174454 497414 209898
rect 496794 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 497414 174454
rect 496794 174134 497414 174218
rect 496794 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 497414 174134
rect 496794 138454 497414 173898
rect 496794 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 497414 138454
rect 496794 138134 497414 138218
rect 496794 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 497414 138134
rect 496794 102454 497414 137898
rect 496794 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 497414 102454
rect 496794 102134 497414 102218
rect 496794 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 497414 102134
rect 496794 66454 497414 101898
rect 496794 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 497414 66454
rect 496794 66134 497414 66218
rect 496794 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 497414 66134
rect 496794 30454 497414 65898
rect 496794 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 497414 30454
rect 496794 30134 497414 30218
rect 496794 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 497414 30134
rect 496794 -6106 497414 29898
rect 496794 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 497414 -6106
rect 496794 -6426 497414 -6342
rect 496794 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 497414 -6426
rect 496794 -7654 497414 -6662
rect 501294 711558 501914 711590
rect 501294 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 501914 711558
rect 501294 711238 501914 711322
rect 501294 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 501914 711238
rect 501294 682954 501914 711002
rect 501294 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 501914 682954
rect 501294 682634 501914 682718
rect 501294 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 501914 682634
rect 501294 646954 501914 682398
rect 501294 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 501914 646954
rect 501294 646634 501914 646718
rect 501294 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 501914 646634
rect 501294 610954 501914 646398
rect 501294 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 501914 610954
rect 501294 610634 501914 610718
rect 501294 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 501914 610634
rect 501294 574954 501914 610398
rect 501294 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 501914 574954
rect 501294 574634 501914 574718
rect 501294 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 501914 574634
rect 501294 538954 501914 574398
rect 501294 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 501914 538954
rect 501294 538634 501914 538718
rect 501294 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 501914 538634
rect 501294 502954 501914 538398
rect 501294 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 501914 502954
rect 501294 502634 501914 502718
rect 501294 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 501914 502634
rect 501294 466954 501914 502398
rect 501294 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 501914 466954
rect 501294 466634 501914 466718
rect 501294 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 501914 466634
rect 501294 430954 501914 466398
rect 501294 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 501914 430954
rect 501294 430634 501914 430718
rect 501294 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 501914 430634
rect 501294 394954 501914 430398
rect 501294 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 501914 394954
rect 501294 394634 501914 394718
rect 501294 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 501914 394634
rect 501294 358954 501914 394398
rect 501294 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 501914 358954
rect 501294 358634 501914 358718
rect 501294 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 501914 358634
rect 501294 322954 501914 358398
rect 501294 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 501914 322954
rect 501294 322634 501914 322718
rect 501294 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 501914 322634
rect 501294 286954 501914 322398
rect 501294 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 501914 286954
rect 501294 286634 501914 286718
rect 501294 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 501914 286634
rect 501294 250954 501914 286398
rect 501294 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 501914 250954
rect 501294 250634 501914 250718
rect 501294 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 501914 250634
rect 501294 214954 501914 250398
rect 501294 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 501914 214954
rect 501294 214634 501914 214718
rect 501294 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 501914 214634
rect 501294 178954 501914 214398
rect 501294 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 501914 178954
rect 501294 178634 501914 178718
rect 501294 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 501914 178634
rect 501294 142954 501914 178398
rect 501294 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 501914 142954
rect 501294 142634 501914 142718
rect 501294 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 501914 142634
rect 501294 106954 501914 142398
rect 501294 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 501914 106954
rect 501294 106634 501914 106718
rect 501294 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 501914 106634
rect 501294 70954 501914 106398
rect 501294 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 501914 70954
rect 501294 70634 501914 70718
rect 501294 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 501914 70634
rect 501294 34954 501914 70398
rect 501294 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 501914 34954
rect 501294 34634 501914 34718
rect 501294 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 501914 34634
rect 501294 -7066 501914 34398
rect 501294 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 501914 -7066
rect 501294 -7386 501914 -7302
rect 501294 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 501914 -7386
rect 501294 -7654 501914 -7622
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 510294 705798 510914 711590
rect 510294 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 510914 705798
rect 510294 705478 510914 705562
rect 510294 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 510914 705478
rect 510294 691954 510914 705242
rect 510294 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 510914 691954
rect 510294 691634 510914 691718
rect 510294 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 510914 691634
rect 510294 655954 510914 691398
rect 510294 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 510914 655954
rect 510294 655634 510914 655718
rect 510294 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 510914 655634
rect 510294 619954 510914 655398
rect 510294 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 510914 619954
rect 510294 619634 510914 619718
rect 510294 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 510914 619634
rect 510294 583954 510914 619398
rect 510294 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 510914 583954
rect 510294 583634 510914 583718
rect 510294 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 510914 583634
rect 510294 547954 510914 583398
rect 510294 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 510914 547954
rect 510294 547634 510914 547718
rect 510294 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 510914 547634
rect 510294 511954 510914 547398
rect 510294 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 510914 511954
rect 510294 511634 510914 511718
rect 510294 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 510914 511634
rect 510294 475954 510914 511398
rect 510294 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 510914 475954
rect 510294 475634 510914 475718
rect 510294 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 510914 475634
rect 510294 439954 510914 475398
rect 510294 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 510914 439954
rect 510294 439634 510914 439718
rect 510294 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 510914 439634
rect 510294 403954 510914 439398
rect 510294 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 510914 403954
rect 510294 403634 510914 403718
rect 510294 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 510914 403634
rect 510294 367954 510914 403398
rect 510294 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 510914 367954
rect 510294 367634 510914 367718
rect 510294 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 510914 367634
rect 510294 331954 510914 367398
rect 510294 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 510914 331954
rect 510294 331634 510914 331718
rect 510294 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 510914 331634
rect 510294 295954 510914 331398
rect 510294 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 510914 295954
rect 510294 295634 510914 295718
rect 510294 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 510914 295634
rect 510294 259954 510914 295398
rect 510294 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 510914 259954
rect 510294 259634 510914 259718
rect 510294 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 510914 259634
rect 510294 223954 510914 259398
rect 510294 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 510914 223954
rect 510294 223634 510914 223718
rect 510294 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 510914 223634
rect 510294 187954 510914 223398
rect 510294 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 510914 187954
rect 510294 187634 510914 187718
rect 510294 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 510914 187634
rect 510294 151954 510914 187398
rect 510294 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 510914 151954
rect 510294 151634 510914 151718
rect 510294 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 510914 151634
rect 510294 115954 510914 151398
rect 510294 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 510914 115954
rect 510294 115634 510914 115718
rect 510294 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 510914 115634
rect 510294 79954 510914 115398
rect 510294 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 510914 79954
rect 510294 79634 510914 79718
rect 510294 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 510914 79634
rect 510294 43954 510914 79398
rect 510294 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 510914 43954
rect 510294 43634 510914 43718
rect 510294 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 510914 43634
rect 510294 7954 510914 43398
rect 510294 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 510914 7954
rect 510294 7634 510914 7718
rect 510294 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 510914 7634
rect 510294 -1306 510914 7398
rect 510294 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 510914 -1306
rect 510294 -1626 510914 -1542
rect 510294 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 510914 -1626
rect 510294 -7654 510914 -1862
rect 514794 706758 515414 711590
rect 514794 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 515414 706758
rect 514794 706438 515414 706522
rect 514794 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 515414 706438
rect 514794 696454 515414 706202
rect 514794 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 515414 696454
rect 514794 696134 515414 696218
rect 514794 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 515414 696134
rect 514794 660454 515414 695898
rect 514794 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 515414 660454
rect 514794 660134 515414 660218
rect 514794 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 515414 660134
rect 514794 624454 515414 659898
rect 514794 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 515414 624454
rect 514794 624134 515414 624218
rect 514794 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 515414 624134
rect 514794 588454 515414 623898
rect 514794 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 515414 588454
rect 514794 588134 515414 588218
rect 514794 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 515414 588134
rect 514794 552454 515414 587898
rect 514794 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 515414 552454
rect 514794 552134 515414 552218
rect 514794 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 515414 552134
rect 514794 516454 515414 551898
rect 514794 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 515414 516454
rect 514794 516134 515414 516218
rect 514794 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 515414 516134
rect 514794 480454 515414 515898
rect 514794 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 515414 480454
rect 514794 480134 515414 480218
rect 514794 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 515414 480134
rect 514794 444454 515414 479898
rect 514794 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 515414 444454
rect 514794 444134 515414 444218
rect 514794 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 515414 444134
rect 514794 408454 515414 443898
rect 514794 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 515414 408454
rect 514794 408134 515414 408218
rect 514794 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 515414 408134
rect 514794 372454 515414 407898
rect 514794 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 515414 372454
rect 514794 372134 515414 372218
rect 514794 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 515414 372134
rect 514794 336454 515414 371898
rect 514794 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 515414 336454
rect 514794 336134 515414 336218
rect 514794 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 515414 336134
rect 514794 300454 515414 335898
rect 514794 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 515414 300454
rect 514794 300134 515414 300218
rect 514794 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 515414 300134
rect 514794 264454 515414 299898
rect 514794 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 515414 264454
rect 514794 264134 515414 264218
rect 514794 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 515414 264134
rect 514794 228454 515414 263898
rect 514794 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 515414 228454
rect 514794 228134 515414 228218
rect 514794 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 515414 228134
rect 514794 192454 515414 227898
rect 514794 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 515414 192454
rect 514794 192134 515414 192218
rect 514794 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 515414 192134
rect 514794 156454 515414 191898
rect 514794 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 515414 156454
rect 514794 156134 515414 156218
rect 514794 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 515414 156134
rect 514794 120454 515414 155898
rect 514794 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 515414 120454
rect 514794 120134 515414 120218
rect 514794 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 515414 120134
rect 514794 84454 515414 119898
rect 514794 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 515414 84454
rect 514794 84134 515414 84218
rect 514794 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 515414 84134
rect 514794 48454 515414 83898
rect 514794 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 515414 48454
rect 514794 48134 515414 48218
rect 514794 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 515414 48134
rect 514794 12454 515414 47898
rect 514794 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 515414 12454
rect 514794 12134 515414 12218
rect 514794 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 515414 12134
rect 514794 -2266 515414 11898
rect 514794 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 515414 -2266
rect 514794 -2586 515414 -2502
rect 514794 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 515414 -2586
rect 514794 -7654 515414 -2822
rect 519294 707718 519914 711590
rect 519294 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 519914 707718
rect 519294 707398 519914 707482
rect 519294 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 519914 707398
rect 519294 700954 519914 707162
rect 519294 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 519914 700954
rect 519294 700634 519914 700718
rect 519294 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 519914 700634
rect 519294 664954 519914 700398
rect 519294 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 519914 664954
rect 519294 664634 519914 664718
rect 519294 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 519914 664634
rect 519294 628954 519914 664398
rect 519294 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 519914 628954
rect 519294 628634 519914 628718
rect 519294 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 519914 628634
rect 519294 592954 519914 628398
rect 519294 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 519914 592954
rect 519294 592634 519914 592718
rect 519294 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 519914 592634
rect 519294 556954 519914 592398
rect 519294 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 519914 556954
rect 519294 556634 519914 556718
rect 519294 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 519914 556634
rect 519294 520954 519914 556398
rect 519294 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 519914 520954
rect 519294 520634 519914 520718
rect 519294 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 519914 520634
rect 519294 484954 519914 520398
rect 519294 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 519914 484954
rect 519294 484634 519914 484718
rect 519294 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 519914 484634
rect 519294 448954 519914 484398
rect 519294 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 519914 448954
rect 519294 448634 519914 448718
rect 519294 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 519914 448634
rect 519294 412954 519914 448398
rect 519294 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 519914 412954
rect 519294 412634 519914 412718
rect 519294 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 519914 412634
rect 519294 376954 519914 412398
rect 519294 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 519914 376954
rect 519294 376634 519914 376718
rect 519294 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 519914 376634
rect 519294 340954 519914 376398
rect 519294 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 519914 340954
rect 519294 340634 519914 340718
rect 519294 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 519914 340634
rect 519294 304954 519914 340398
rect 519294 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 519914 304954
rect 519294 304634 519914 304718
rect 519294 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 519914 304634
rect 519294 268954 519914 304398
rect 519294 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 519914 268954
rect 519294 268634 519914 268718
rect 519294 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 519914 268634
rect 519294 232954 519914 268398
rect 519294 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 519914 232954
rect 519294 232634 519914 232718
rect 519294 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 519914 232634
rect 519294 196954 519914 232398
rect 519294 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 519914 196954
rect 519294 196634 519914 196718
rect 519294 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 519914 196634
rect 519294 160954 519914 196398
rect 519294 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 519914 160954
rect 519294 160634 519914 160718
rect 519294 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 519914 160634
rect 519294 124954 519914 160398
rect 519294 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 519914 124954
rect 519294 124634 519914 124718
rect 519294 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 519914 124634
rect 519294 88954 519914 124398
rect 519294 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 519914 88954
rect 519294 88634 519914 88718
rect 519294 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 519914 88634
rect 519294 52954 519914 88398
rect 519294 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 519914 52954
rect 519294 52634 519914 52718
rect 519294 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 519914 52634
rect 519294 16954 519914 52398
rect 519294 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 519914 16954
rect 519294 16634 519914 16718
rect 519294 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 519914 16634
rect 519294 -3226 519914 16398
rect 519294 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 519914 -3226
rect 519294 -3546 519914 -3462
rect 519294 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 519914 -3546
rect 519294 -7654 519914 -3782
rect 523794 708678 524414 711590
rect 523794 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 524414 708678
rect 523794 708358 524414 708442
rect 523794 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 524414 708358
rect 523794 669454 524414 708122
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -4186 524414 20898
rect 523794 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 524414 -4186
rect 523794 -4506 524414 -4422
rect 523794 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 524414 -4506
rect 523794 -7654 524414 -4742
rect 528294 709638 528914 711590
rect 528294 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 528914 709638
rect 528294 709318 528914 709402
rect 528294 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 528914 709318
rect 528294 673954 528914 709082
rect 528294 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 528914 673954
rect 528294 673634 528914 673718
rect 528294 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 528914 673634
rect 528294 637954 528914 673398
rect 528294 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 528914 637954
rect 528294 637634 528914 637718
rect 528294 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 528914 637634
rect 528294 601954 528914 637398
rect 528294 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 528914 601954
rect 528294 601634 528914 601718
rect 528294 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 528914 601634
rect 528294 565954 528914 601398
rect 528294 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 528914 565954
rect 528294 565634 528914 565718
rect 528294 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 528914 565634
rect 528294 529954 528914 565398
rect 528294 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 528914 529954
rect 528294 529634 528914 529718
rect 528294 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 528914 529634
rect 528294 493954 528914 529398
rect 528294 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 528914 493954
rect 528294 493634 528914 493718
rect 528294 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 528914 493634
rect 528294 457954 528914 493398
rect 528294 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 528914 457954
rect 528294 457634 528914 457718
rect 528294 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 528914 457634
rect 528294 421954 528914 457398
rect 528294 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 528914 421954
rect 528294 421634 528914 421718
rect 528294 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 528914 421634
rect 528294 385954 528914 421398
rect 528294 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 528914 385954
rect 528294 385634 528914 385718
rect 528294 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 528914 385634
rect 528294 349954 528914 385398
rect 528294 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 528914 349954
rect 528294 349634 528914 349718
rect 528294 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 528914 349634
rect 528294 313954 528914 349398
rect 528294 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 528914 313954
rect 528294 313634 528914 313718
rect 528294 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 528914 313634
rect 528294 277954 528914 313398
rect 528294 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 528914 277954
rect 528294 277634 528914 277718
rect 528294 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 528914 277634
rect 528294 241954 528914 277398
rect 528294 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 528914 241954
rect 528294 241634 528914 241718
rect 528294 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 528914 241634
rect 528294 205954 528914 241398
rect 528294 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 528914 205954
rect 528294 205634 528914 205718
rect 528294 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 528914 205634
rect 528294 169954 528914 205398
rect 528294 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 528914 169954
rect 528294 169634 528914 169718
rect 528294 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 528914 169634
rect 528294 133954 528914 169398
rect 528294 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 528914 133954
rect 528294 133634 528914 133718
rect 528294 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 528914 133634
rect 528294 97954 528914 133398
rect 528294 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 528914 97954
rect 528294 97634 528914 97718
rect 528294 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 528914 97634
rect 528294 61954 528914 97398
rect 528294 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 528914 61954
rect 528294 61634 528914 61718
rect 528294 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 528914 61634
rect 528294 25954 528914 61398
rect 528294 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 528914 25954
rect 528294 25634 528914 25718
rect 528294 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 528914 25634
rect 528294 -5146 528914 25398
rect 528294 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 528914 -5146
rect 528294 -5466 528914 -5382
rect 528294 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 528914 -5466
rect 528294 -7654 528914 -5702
rect 532794 710598 533414 711590
rect 532794 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 533414 710598
rect 532794 710278 533414 710362
rect 532794 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 533414 710278
rect 532794 678454 533414 710042
rect 532794 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 533414 678454
rect 532794 678134 533414 678218
rect 532794 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 533414 678134
rect 532794 642454 533414 677898
rect 532794 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 533414 642454
rect 532794 642134 533414 642218
rect 532794 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 533414 642134
rect 532794 606454 533414 641898
rect 532794 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 533414 606454
rect 532794 606134 533414 606218
rect 532794 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 533414 606134
rect 532794 570454 533414 605898
rect 532794 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 533414 570454
rect 532794 570134 533414 570218
rect 532794 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 533414 570134
rect 532794 534454 533414 569898
rect 532794 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 533414 534454
rect 532794 534134 533414 534218
rect 532794 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 533414 534134
rect 532794 498454 533414 533898
rect 532794 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 533414 498454
rect 532794 498134 533414 498218
rect 532794 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 533414 498134
rect 532794 462454 533414 497898
rect 532794 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 533414 462454
rect 532794 462134 533414 462218
rect 532794 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 533414 462134
rect 532794 426454 533414 461898
rect 532794 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 533414 426454
rect 532794 426134 533414 426218
rect 532794 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 533414 426134
rect 532794 390454 533414 425898
rect 532794 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 533414 390454
rect 532794 390134 533414 390218
rect 532794 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 533414 390134
rect 532794 354454 533414 389898
rect 532794 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 533414 354454
rect 532794 354134 533414 354218
rect 532794 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 533414 354134
rect 532794 318454 533414 353898
rect 532794 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 533414 318454
rect 532794 318134 533414 318218
rect 532794 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 533414 318134
rect 532794 282454 533414 317898
rect 532794 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 533414 282454
rect 532794 282134 533414 282218
rect 532794 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 533414 282134
rect 532794 246454 533414 281898
rect 532794 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 533414 246454
rect 532794 246134 533414 246218
rect 532794 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 533414 246134
rect 532794 210454 533414 245898
rect 532794 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 533414 210454
rect 532794 210134 533414 210218
rect 532794 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 533414 210134
rect 532794 174454 533414 209898
rect 532794 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 533414 174454
rect 532794 174134 533414 174218
rect 532794 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 533414 174134
rect 532794 138454 533414 173898
rect 532794 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 533414 138454
rect 532794 138134 533414 138218
rect 532794 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 533414 138134
rect 532794 102454 533414 137898
rect 532794 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 533414 102454
rect 532794 102134 533414 102218
rect 532794 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 533414 102134
rect 532794 66454 533414 101898
rect 532794 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 533414 66454
rect 532794 66134 533414 66218
rect 532794 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 533414 66134
rect 532794 30454 533414 65898
rect 532794 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 533414 30454
rect 532794 30134 533414 30218
rect 532794 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 533414 30134
rect 532794 -6106 533414 29898
rect 532794 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 533414 -6106
rect 532794 -6426 533414 -6342
rect 532794 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 533414 -6426
rect 532794 -7654 533414 -6662
rect 537294 711558 537914 711590
rect 537294 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 537914 711558
rect 537294 711238 537914 711322
rect 537294 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 537914 711238
rect 537294 682954 537914 711002
rect 537294 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 537914 682954
rect 537294 682634 537914 682718
rect 537294 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 537914 682634
rect 537294 646954 537914 682398
rect 537294 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 537914 646954
rect 537294 646634 537914 646718
rect 537294 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 537914 646634
rect 537294 610954 537914 646398
rect 537294 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 537914 610954
rect 537294 610634 537914 610718
rect 537294 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 537914 610634
rect 537294 574954 537914 610398
rect 537294 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 537914 574954
rect 537294 574634 537914 574718
rect 537294 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 537914 574634
rect 537294 538954 537914 574398
rect 537294 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 537914 538954
rect 537294 538634 537914 538718
rect 537294 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 537914 538634
rect 537294 502954 537914 538398
rect 537294 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 537914 502954
rect 537294 502634 537914 502718
rect 537294 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 537914 502634
rect 537294 466954 537914 502398
rect 537294 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 537914 466954
rect 537294 466634 537914 466718
rect 537294 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 537914 466634
rect 537294 430954 537914 466398
rect 537294 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 537914 430954
rect 537294 430634 537914 430718
rect 537294 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 537914 430634
rect 537294 394954 537914 430398
rect 537294 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 537914 394954
rect 537294 394634 537914 394718
rect 537294 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 537914 394634
rect 537294 358954 537914 394398
rect 537294 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 537914 358954
rect 537294 358634 537914 358718
rect 537294 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 537914 358634
rect 537294 322954 537914 358398
rect 537294 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 537914 322954
rect 537294 322634 537914 322718
rect 537294 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 537914 322634
rect 537294 286954 537914 322398
rect 537294 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 537914 286954
rect 537294 286634 537914 286718
rect 537294 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 537914 286634
rect 537294 250954 537914 286398
rect 537294 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 537914 250954
rect 537294 250634 537914 250718
rect 537294 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 537914 250634
rect 537294 214954 537914 250398
rect 537294 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 537914 214954
rect 537294 214634 537914 214718
rect 537294 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 537914 214634
rect 537294 178954 537914 214398
rect 537294 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 537914 178954
rect 537294 178634 537914 178718
rect 537294 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 537914 178634
rect 537294 142954 537914 178398
rect 537294 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 537914 142954
rect 537294 142634 537914 142718
rect 537294 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 537914 142634
rect 537294 106954 537914 142398
rect 537294 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 537914 106954
rect 537294 106634 537914 106718
rect 537294 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 537914 106634
rect 537294 70954 537914 106398
rect 537294 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 537914 70954
rect 537294 70634 537914 70718
rect 537294 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 537914 70634
rect 537294 34954 537914 70398
rect 537294 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 537914 34954
rect 537294 34634 537914 34718
rect 537294 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 537914 34634
rect 537294 -7066 537914 34398
rect 537294 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 537914 -7066
rect 537294 -7386 537914 -7302
rect 537294 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 537914 -7386
rect 537294 -7654 537914 -7622
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 546294 705798 546914 711590
rect 546294 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 546914 705798
rect 546294 705478 546914 705562
rect 546294 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 546914 705478
rect 546294 691954 546914 705242
rect 546294 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 546914 691954
rect 546294 691634 546914 691718
rect 546294 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 546914 691634
rect 546294 655954 546914 691398
rect 546294 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 546914 655954
rect 546294 655634 546914 655718
rect 546294 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 546914 655634
rect 546294 619954 546914 655398
rect 546294 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 546914 619954
rect 546294 619634 546914 619718
rect 546294 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 546914 619634
rect 546294 583954 546914 619398
rect 546294 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 546914 583954
rect 546294 583634 546914 583718
rect 546294 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 546914 583634
rect 546294 547954 546914 583398
rect 546294 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 546914 547954
rect 546294 547634 546914 547718
rect 546294 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 546914 547634
rect 546294 511954 546914 547398
rect 546294 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 546914 511954
rect 546294 511634 546914 511718
rect 546294 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 546914 511634
rect 546294 475954 546914 511398
rect 546294 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 546914 475954
rect 546294 475634 546914 475718
rect 546294 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 546914 475634
rect 546294 439954 546914 475398
rect 546294 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 546914 439954
rect 546294 439634 546914 439718
rect 546294 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 546914 439634
rect 546294 403954 546914 439398
rect 546294 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 546914 403954
rect 546294 403634 546914 403718
rect 546294 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 546914 403634
rect 546294 367954 546914 403398
rect 546294 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 546914 367954
rect 546294 367634 546914 367718
rect 546294 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 546914 367634
rect 546294 331954 546914 367398
rect 546294 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 546914 331954
rect 546294 331634 546914 331718
rect 546294 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 546914 331634
rect 546294 295954 546914 331398
rect 546294 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 546914 295954
rect 546294 295634 546914 295718
rect 546294 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 546914 295634
rect 546294 259954 546914 295398
rect 546294 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 546914 259954
rect 546294 259634 546914 259718
rect 546294 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 546914 259634
rect 546294 223954 546914 259398
rect 546294 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 546914 223954
rect 546294 223634 546914 223718
rect 546294 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 546914 223634
rect 546294 187954 546914 223398
rect 546294 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 546914 187954
rect 546294 187634 546914 187718
rect 546294 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 546914 187634
rect 546294 151954 546914 187398
rect 546294 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 546914 151954
rect 546294 151634 546914 151718
rect 546294 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 546914 151634
rect 546294 115954 546914 151398
rect 546294 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 546914 115954
rect 546294 115634 546914 115718
rect 546294 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 546914 115634
rect 546294 79954 546914 115398
rect 546294 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 546914 79954
rect 546294 79634 546914 79718
rect 546294 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 546914 79634
rect 546294 43954 546914 79398
rect 546294 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 546914 43954
rect 546294 43634 546914 43718
rect 546294 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 546914 43634
rect 546294 7954 546914 43398
rect 546294 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 546914 7954
rect 546294 7634 546914 7718
rect 546294 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 546914 7634
rect 546294 -1306 546914 7398
rect 546294 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 546914 -1306
rect 546294 -1626 546914 -1542
rect 546294 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 546914 -1626
rect 546294 -7654 546914 -1862
rect 550794 706758 551414 711590
rect 550794 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 551414 706758
rect 550794 706438 551414 706522
rect 550794 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 551414 706438
rect 550794 696454 551414 706202
rect 550794 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 551414 696454
rect 550794 696134 551414 696218
rect 550794 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 551414 696134
rect 550794 660454 551414 695898
rect 550794 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 551414 660454
rect 550794 660134 551414 660218
rect 550794 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 551414 660134
rect 550794 624454 551414 659898
rect 550794 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 551414 624454
rect 550794 624134 551414 624218
rect 550794 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 551414 624134
rect 550794 588454 551414 623898
rect 550794 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 551414 588454
rect 550794 588134 551414 588218
rect 550794 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 551414 588134
rect 550794 552454 551414 587898
rect 550794 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 551414 552454
rect 550794 552134 551414 552218
rect 550794 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 551414 552134
rect 550794 516454 551414 551898
rect 550794 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 551414 516454
rect 550794 516134 551414 516218
rect 550794 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 551414 516134
rect 550794 480454 551414 515898
rect 550794 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 551414 480454
rect 550794 480134 551414 480218
rect 550794 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 551414 480134
rect 550794 444454 551414 479898
rect 550794 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 551414 444454
rect 550794 444134 551414 444218
rect 550794 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 551414 444134
rect 550794 408454 551414 443898
rect 550794 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 551414 408454
rect 550794 408134 551414 408218
rect 550794 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 551414 408134
rect 550794 372454 551414 407898
rect 550794 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 551414 372454
rect 550794 372134 551414 372218
rect 550794 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 551414 372134
rect 550794 336454 551414 371898
rect 550794 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 551414 336454
rect 550794 336134 551414 336218
rect 550794 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 551414 336134
rect 550794 300454 551414 335898
rect 550794 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 551414 300454
rect 550794 300134 551414 300218
rect 550794 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 551414 300134
rect 550794 264454 551414 299898
rect 550794 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 551414 264454
rect 550794 264134 551414 264218
rect 550794 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 551414 264134
rect 550794 228454 551414 263898
rect 550794 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 551414 228454
rect 550794 228134 551414 228218
rect 550794 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 551414 228134
rect 550794 192454 551414 227898
rect 550794 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 551414 192454
rect 550794 192134 551414 192218
rect 550794 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 551414 192134
rect 550794 156454 551414 191898
rect 550794 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 551414 156454
rect 550794 156134 551414 156218
rect 550794 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 551414 156134
rect 550794 120454 551414 155898
rect 550794 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 551414 120454
rect 550794 120134 551414 120218
rect 550794 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 551414 120134
rect 550794 84454 551414 119898
rect 550794 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 551414 84454
rect 550794 84134 551414 84218
rect 550794 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 551414 84134
rect 550794 48454 551414 83898
rect 550794 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 551414 48454
rect 550794 48134 551414 48218
rect 550794 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 551414 48134
rect 550794 12454 551414 47898
rect 550794 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 551414 12454
rect 550794 12134 551414 12218
rect 550794 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 551414 12134
rect 550794 -2266 551414 11898
rect 550794 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 551414 -2266
rect 550794 -2586 551414 -2502
rect 550794 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 551414 -2586
rect 550794 -7654 551414 -2822
rect 555294 707718 555914 711590
rect 555294 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 555914 707718
rect 555294 707398 555914 707482
rect 555294 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 555914 707398
rect 555294 700954 555914 707162
rect 555294 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 555914 700954
rect 555294 700634 555914 700718
rect 555294 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 555914 700634
rect 555294 664954 555914 700398
rect 555294 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 555914 664954
rect 555294 664634 555914 664718
rect 555294 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 555914 664634
rect 555294 628954 555914 664398
rect 555294 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 555914 628954
rect 555294 628634 555914 628718
rect 555294 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 555914 628634
rect 555294 592954 555914 628398
rect 555294 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 555914 592954
rect 555294 592634 555914 592718
rect 555294 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 555914 592634
rect 555294 556954 555914 592398
rect 555294 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 555914 556954
rect 555294 556634 555914 556718
rect 555294 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 555914 556634
rect 555294 520954 555914 556398
rect 555294 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 555914 520954
rect 555294 520634 555914 520718
rect 555294 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 555914 520634
rect 555294 484954 555914 520398
rect 555294 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 555914 484954
rect 555294 484634 555914 484718
rect 555294 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 555914 484634
rect 555294 448954 555914 484398
rect 555294 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 555914 448954
rect 555294 448634 555914 448718
rect 555294 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 555914 448634
rect 555294 412954 555914 448398
rect 555294 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 555914 412954
rect 555294 412634 555914 412718
rect 555294 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 555914 412634
rect 555294 376954 555914 412398
rect 555294 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 555914 376954
rect 555294 376634 555914 376718
rect 555294 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 555914 376634
rect 555294 340954 555914 376398
rect 555294 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 555914 340954
rect 555294 340634 555914 340718
rect 555294 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 555914 340634
rect 555294 304954 555914 340398
rect 555294 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 555914 304954
rect 555294 304634 555914 304718
rect 555294 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 555914 304634
rect 555294 268954 555914 304398
rect 555294 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 555914 268954
rect 555294 268634 555914 268718
rect 555294 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 555914 268634
rect 555294 232954 555914 268398
rect 555294 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 555914 232954
rect 555294 232634 555914 232718
rect 555294 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 555914 232634
rect 555294 196954 555914 232398
rect 555294 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 555914 196954
rect 555294 196634 555914 196718
rect 555294 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 555914 196634
rect 555294 160954 555914 196398
rect 555294 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 555914 160954
rect 555294 160634 555914 160718
rect 555294 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 555914 160634
rect 555294 124954 555914 160398
rect 555294 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 555914 124954
rect 555294 124634 555914 124718
rect 555294 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 555914 124634
rect 555294 88954 555914 124398
rect 555294 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 555914 88954
rect 555294 88634 555914 88718
rect 555294 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 555914 88634
rect 555294 52954 555914 88398
rect 555294 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 555914 52954
rect 555294 52634 555914 52718
rect 555294 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 555914 52634
rect 555294 16954 555914 52398
rect 555294 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 555914 16954
rect 555294 16634 555914 16718
rect 555294 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 555914 16634
rect 555294 -3226 555914 16398
rect 555294 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 555914 -3226
rect 555294 -3546 555914 -3462
rect 555294 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 555914 -3546
rect 555294 -7654 555914 -3782
rect 559794 708678 560414 711590
rect 559794 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 560414 708678
rect 559794 708358 560414 708442
rect 559794 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 560414 708358
rect 559794 669454 560414 708122
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -4186 560414 20898
rect 559794 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 560414 -4186
rect 559794 -4506 560414 -4422
rect 559794 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 560414 -4506
rect 559794 -7654 560414 -4742
rect 564294 709638 564914 711590
rect 564294 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 564914 709638
rect 564294 709318 564914 709402
rect 564294 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 564914 709318
rect 564294 673954 564914 709082
rect 564294 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 564914 673954
rect 564294 673634 564914 673718
rect 564294 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 564914 673634
rect 564294 637954 564914 673398
rect 564294 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 564914 637954
rect 564294 637634 564914 637718
rect 564294 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 564914 637634
rect 564294 601954 564914 637398
rect 564294 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 564914 601954
rect 564294 601634 564914 601718
rect 564294 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 564914 601634
rect 564294 565954 564914 601398
rect 564294 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 564914 565954
rect 564294 565634 564914 565718
rect 564294 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 564914 565634
rect 564294 529954 564914 565398
rect 564294 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 564914 529954
rect 564294 529634 564914 529718
rect 564294 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 564914 529634
rect 564294 493954 564914 529398
rect 564294 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 564914 493954
rect 564294 493634 564914 493718
rect 564294 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 564914 493634
rect 564294 457954 564914 493398
rect 564294 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 564914 457954
rect 564294 457634 564914 457718
rect 564294 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 564914 457634
rect 564294 421954 564914 457398
rect 564294 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 564914 421954
rect 564294 421634 564914 421718
rect 564294 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 564914 421634
rect 564294 385954 564914 421398
rect 564294 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 564914 385954
rect 564294 385634 564914 385718
rect 564294 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 564914 385634
rect 564294 349954 564914 385398
rect 564294 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 564914 349954
rect 564294 349634 564914 349718
rect 564294 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 564914 349634
rect 564294 313954 564914 349398
rect 564294 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 564914 313954
rect 564294 313634 564914 313718
rect 564294 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 564914 313634
rect 564294 277954 564914 313398
rect 564294 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 564914 277954
rect 564294 277634 564914 277718
rect 564294 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 564914 277634
rect 564294 241954 564914 277398
rect 564294 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 564914 241954
rect 564294 241634 564914 241718
rect 564294 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 564914 241634
rect 564294 205954 564914 241398
rect 564294 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 564914 205954
rect 564294 205634 564914 205718
rect 564294 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 564914 205634
rect 564294 169954 564914 205398
rect 564294 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 564914 169954
rect 564294 169634 564914 169718
rect 564294 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 564914 169634
rect 564294 133954 564914 169398
rect 564294 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 564914 133954
rect 564294 133634 564914 133718
rect 564294 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 564914 133634
rect 564294 97954 564914 133398
rect 564294 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 564914 97954
rect 564294 97634 564914 97718
rect 564294 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 564914 97634
rect 564294 61954 564914 97398
rect 564294 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 564914 61954
rect 564294 61634 564914 61718
rect 564294 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 564914 61634
rect 564294 25954 564914 61398
rect 564294 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 564914 25954
rect 564294 25634 564914 25718
rect 564294 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 564914 25634
rect 564294 -5146 564914 25398
rect 564294 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 564914 -5146
rect 564294 -5466 564914 -5382
rect 564294 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 564914 -5466
rect 564294 -7654 564914 -5702
rect 568794 710598 569414 711590
rect 568794 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 569414 710598
rect 568794 710278 569414 710362
rect 568794 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 569414 710278
rect 568794 678454 569414 710042
rect 568794 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 569414 678454
rect 568794 678134 569414 678218
rect 568794 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 569414 678134
rect 568794 642454 569414 677898
rect 568794 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 569414 642454
rect 568794 642134 569414 642218
rect 568794 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 569414 642134
rect 568794 606454 569414 641898
rect 568794 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 569414 606454
rect 568794 606134 569414 606218
rect 568794 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 569414 606134
rect 568794 570454 569414 605898
rect 568794 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 569414 570454
rect 568794 570134 569414 570218
rect 568794 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 569414 570134
rect 568794 534454 569414 569898
rect 568794 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 569414 534454
rect 568794 534134 569414 534218
rect 568794 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 569414 534134
rect 568794 498454 569414 533898
rect 568794 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 569414 498454
rect 568794 498134 569414 498218
rect 568794 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 569414 498134
rect 568794 462454 569414 497898
rect 568794 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 569414 462454
rect 568794 462134 569414 462218
rect 568794 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 569414 462134
rect 568794 426454 569414 461898
rect 568794 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 569414 426454
rect 568794 426134 569414 426218
rect 568794 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 569414 426134
rect 568794 390454 569414 425898
rect 568794 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 569414 390454
rect 568794 390134 569414 390218
rect 568794 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 569414 390134
rect 568794 354454 569414 389898
rect 568794 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 569414 354454
rect 568794 354134 569414 354218
rect 568794 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 569414 354134
rect 568794 318454 569414 353898
rect 568794 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 569414 318454
rect 568794 318134 569414 318218
rect 568794 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 569414 318134
rect 568794 282454 569414 317898
rect 568794 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 569414 282454
rect 568794 282134 569414 282218
rect 568794 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 569414 282134
rect 568794 246454 569414 281898
rect 568794 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 569414 246454
rect 568794 246134 569414 246218
rect 568794 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 569414 246134
rect 568794 210454 569414 245898
rect 568794 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 569414 210454
rect 568794 210134 569414 210218
rect 568794 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 569414 210134
rect 568794 174454 569414 209898
rect 568794 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 569414 174454
rect 568794 174134 569414 174218
rect 568794 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 569414 174134
rect 568794 138454 569414 173898
rect 568794 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 569414 138454
rect 568794 138134 569414 138218
rect 568794 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 569414 138134
rect 568794 102454 569414 137898
rect 568794 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 569414 102454
rect 568794 102134 569414 102218
rect 568794 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 569414 102134
rect 568794 66454 569414 101898
rect 568794 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 569414 66454
rect 568794 66134 569414 66218
rect 568794 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 569414 66134
rect 568794 30454 569414 65898
rect 568794 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 569414 30454
rect 568794 30134 569414 30218
rect 568794 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 569414 30134
rect 568794 -6106 569414 29898
rect 568794 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 569414 -6106
rect 568794 -6426 569414 -6342
rect 568794 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 569414 -6426
rect 568794 -7654 569414 -6662
rect 573294 711558 573914 711590
rect 573294 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 573914 711558
rect 573294 711238 573914 711322
rect 573294 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 573914 711238
rect 573294 682954 573914 711002
rect 573294 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 573914 682954
rect 573294 682634 573914 682718
rect 573294 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 573914 682634
rect 573294 646954 573914 682398
rect 573294 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 573914 646954
rect 573294 646634 573914 646718
rect 573294 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 573914 646634
rect 573294 610954 573914 646398
rect 573294 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 573914 610954
rect 573294 610634 573914 610718
rect 573294 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 573914 610634
rect 573294 574954 573914 610398
rect 573294 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 573914 574954
rect 573294 574634 573914 574718
rect 573294 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 573914 574634
rect 573294 538954 573914 574398
rect 573294 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 573914 538954
rect 573294 538634 573914 538718
rect 573294 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 573914 538634
rect 573294 502954 573914 538398
rect 573294 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 573914 502954
rect 573294 502634 573914 502718
rect 573294 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 573914 502634
rect 573294 466954 573914 502398
rect 573294 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 573914 466954
rect 573294 466634 573914 466718
rect 573294 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 573914 466634
rect 573294 430954 573914 466398
rect 573294 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 573914 430954
rect 573294 430634 573914 430718
rect 573294 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 573914 430634
rect 573294 394954 573914 430398
rect 573294 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 573914 394954
rect 573294 394634 573914 394718
rect 573294 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 573914 394634
rect 573294 358954 573914 394398
rect 573294 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 573914 358954
rect 573294 358634 573914 358718
rect 573294 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 573914 358634
rect 573294 322954 573914 358398
rect 573294 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 573914 322954
rect 573294 322634 573914 322718
rect 573294 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 573914 322634
rect 573294 286954 573914 322398
rect 573294 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 573914 286954
rect 573294 286634 573914 286718
rect 573294 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 573914 286634
rect 573294 250954 573914 286398
rect 573294 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 573914 250954
rect 573294 250634 573914 250718
rect 573294 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 573914 250634
rect 573294 214954 573914 250398
rect 573294 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 573914 214954
rect 573294 214634 573914 214718
rect 573294 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 573914 214634
rect 573294 178954 573914 214398
rect 573294 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 573914 178954
rect 573294 178634 573914 178718
rect 573294 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 573914 178634
rect 573294 142954 573914 178398
rect 573294 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 573914 142954
rect 573294 142634 573914 142718
rect 573294 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 573914 142634
rect 573294 106954 573914 142398
rect 573294 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 573914 106954
rect 573294 106634 573914 106718
rect 573294 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 573914 106634
rect 573294 70954 573914 106398
rect 573294 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 573914 70954
rect 573294 70634 573914 70718
rect 573294 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 573914 70634
rect 573294 34954 573914 70398
rect 573294 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 573914 34954
rect 573294 34634 573914 34718
rect 573294 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 573914 34634
rect 573294 -7066 573914 34398
rect 573294 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 573914 -7066
rect 573294 -7386 573914 -7302
rect 573294 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 573914 -7386
rect 573294 -7654 573914 -7622
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 582294 705798 582914 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 582294 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 582914 705798
rect 582294 705478 582914 705562
rect 582294 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 582914 705478
rect 580763 697236 580829 697237
rect 580763 697172 580764 697236
rect 580828 697172 580829 697236
rect 580763 697171 580829 697172
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 580766 75309 580826 697171
rect 582294 691954 582914 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 582294 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 582914 691954
rect 582294 691634 582914 691718
rect 582294 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 582914 691634
rect 582294 655954 582914 691398
rect 582294 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 582914 655954
rect 582294 655634 582914 655718
rect 582294 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 582914 655634
rect 582294 619954 582914 655398
rect 582294 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 582914 619954
rect 582294 619634 582914 619718
rect 582294 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 582914 619634
rect 582294 583954 582914 619398
rect 582294 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 582914 583954
rect 582294 583634 582914 583718
rect 582294 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 582914 583634
rect 582294 547954 582914 583398
rect 582294 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 582914 547954
rect 582294 547634 582914 547718
rect 582294 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 582914 547634
rect 582294 511954 582914 547398
rect 582294 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 582914 511954
rect 582294 511634 582914 511718
rect 582294 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 582914 511634
rect 582294 475954 582914 511398
rect 582294 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 582914 475954
rect 582294 475634 582914 475718
rect 582294 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 582914 475634
rect 582294 439954 582914 475398
rect 582294 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 582914 439954
rect 582294 439634 582914 439718
rect 582294 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 582914 439634
rect 582294 403954 582914 439398
rect 582294 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 582914 403954
rect 582294 403634 582914 403718
rect 582294 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 582914 403634
rect 582294 367954 582914 403398
rect 582294 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 582914 367954
rect 582294 367634 582914 367718
rect 582294 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 582914 367634
rect 582294 331954 582914 367398
rect 582294 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 582914 331954
rect 582294 331634 582914 331718
rect 582294 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 582914 331634
rect 582294 295954 582914 331398
rect 582294 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 582914 295954
rect 582294 295634 582914 295718
rect 582294 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 582914 295634
rect 582294 259954 582914 295398
rect 582294 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 582914 259954
rect 582294 259634 582914 259718
rect 582294 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 582914 259634
rect 582294 223954 582914 259398
rect 582294 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 582914 223954
rect 582294 223634 582914 223718
rect 582294 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 582914 223634
rect 582294 187954 582914 223398
rect 582294 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 582914 187954
rect 582294 187634 582914 187718
rect 582294 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 582914 187634
rect 582294 151954 582914 187398
rect 582294 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 582914 151954
rect 582294 151634 582914 151718
rect 582294 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 582914 151634
rect 582294 115954 582914 151398
rect 582294 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 582914 115954
rect 582294 115634 582914 115718
rect 582294 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 582914 115634
rect 582294 79954 582914 115398
rect 582294 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 582914 79954
rect 582294 79634 582914 79718
rect 582294 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 582914 79634
rect 580763 75308 580829 75309
rect 580763 75244 580764 75308
rect 580828 75244 580829 75308
rect 580763 75243 580829 75244
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 582294 43954 582914 79398
rect 582294 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 582914 43954
rect 582294 43634 582914 43718
rect 582294 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 582914 43634
rect 582294 7954 582914 43398
rect 582294 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 582914 7954
rect 582294 7634 582914 7718
rect 582294 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 582914 7634
rect 582294 -1306 582914 7398
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691954 586890 705242
rect 586270 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 586890 691954
rect 586270 691634 586890 691718
rect 586270 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 586890 691634
rect 586270 655954 586890 691398
rect 586270 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 586890 655954
rect 586270 655634 586890 655718
rect 586270 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 586890 655634
rect 586270 619954 586890 655398
rect 586270 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 586890 619954
rect 586270 619634 586890 619718
rect 586270 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 586890 619634
rect 586270 583954 586890 619398
rect 586270 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 586890 583954
rect 586270 583634 586890 583718
rect 586270 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 586890 583634
rect 586270 547954 586890 583398
rect 586270 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 586890 547954
rect 586270 547634 586890 547718
rect 586270 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 586890 547634
rect 586270 511954 586890 547398
rect 586270 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 586890 511954
rect 586270 511634 586890 511718
rect 586270 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 586890 511634
rect 586270 475954 586890 511398
rect 586270 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 586890 475954
rect 586270 475634 586890 475718
rect 586270 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 586890 475634
rect 586270 439954 586890 475398
rect 586270 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 586890 439954
rect 586270 439634 586890 439718
rect 586270 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 586890 439634
rect 586270 403954 586890 439398
rect 586270 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 586890 403954
rect 586270 403634 586890 403718
rect 586270 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 586890 403634
rect 586270 367954 586890 403398
rect 586270 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 586890 367954
rect 586270 367634 586890 367718
rect 586270 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 586890 367634
rect 586270 331954 586890 367398
rect 586270 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 586890 331954
rect 586270 331634 586890 331718
rect 586270 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 586890 331634
rect 586270 295954 586890 331398
rect 586270 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 586890 295954
rect 586270 295634 586890 295718
rect 586270 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 586890 295634
rect 586270 259954 586890 295398
rect 586270 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 586890 259954
rect 586270 259634 586890 259718
rect 586270 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 586890 259634
rect 586270 223954 586890 259398
rect 586270 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 586890 223954
rect 586270 223634 586890 223718
rect 586270 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 586890 223634
rect 586270 187954 586890 223398
rect 586270 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 586890 187954
rect 586270 187634 586890 187718
rect 586270 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 586890 187634
rect 586270 151954 586890 187398
rect 586270 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 586890 151954
rect 586270 151634 586890 151718
rect 586270 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 586890 151634
rect 586270 115954 586890 151398
rect 586270 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 586890 115954
rect 586270 115634 586890 115718
rect 586270 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 586890 115634
rect 586270 79954 586890 115398
rect 586270 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 586890 79954
rect 586270 79634 586890 79718
rect 586270 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 586890 79634
rect 586270 43954 586890 79398
rect 586270 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 586890 43954
rect 586270 43634 586890 43718
rect 586270 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 586890 43634
rect 586270 7954 586890 43398
rect 586270 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 586890 7954
rect 586270 7634 586890 7718
rect 586270 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 586890 7634
rect 582294 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 582914 -1306
rect 582294 -1626 582914 -1542
rect 582294 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 582914 -1626
rect 582294 -7654 582914 -1862
rect 586270 -1306 586890 7398
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 696454 587850 706202
rect 587230 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 587850 696454
rect 587230 696134 587850 696218
rect 587230 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 587850 696134
rect 587230 660454 587850 695898
rect 587230 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 587850 660454
rect 587230 660134 587850 660218
rect 587230 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 587850 660134
rect 587230 624454 587850 659898
rect 587230 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 587850 624454
rect 587230 624134 587850 624218
rect 587230 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 587850 624134
rect 587230 588454 587850 623898
rect 587230 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 587850 588454
rect 587230 588134 587850 588218
rect 587230 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 587850 588134
rect 587230 552454 587850 587898
rect 587230 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 587850 552454
rect 587230 552134 587850 552218
rect 587230 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 587850 552134
rect 587230 516454 587850 551898
rect 587230 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 587850 516454
rect 587230 516134 587850 516218
rect 587230 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 587850 516134
rect 587230 480454 587850 515898
rect 587230 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 587850 480454
rect 587230 480134 587850 480218
rect 587230 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 587850 480134
rect 587230 444454 587850 479898
rect 587230 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 587850 444454
rect 587230 444134 587850 444218
rect 587230 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 587850 444134
rect 587230 408454 587850 443898
rect 587230 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 587850 408454
rect 587230 408134 587850 408218
rect 587230 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 587850 408134
rect 587230 372454 587850 407898
rect 587230 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 587850 372454
rect 587230 372134 587850 372218
rect 587230 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 587850 372134
rect 587230 336454 587850 371898
rect 587230 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 587850 336454
rect 587230 336134 587850 336218
rect 587230 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 587850 336134
rect 587230 300454 587850 335898
rect 587230 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 587850 300454
rect 587230 300134 587850 300218
rect 587230 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 587850 300134
rect 587230 264454 587850 299898
rect 587230 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 587850 264454
rect 587230 264134 587850 264218
rect 587230 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 587850 264134
rect 587230 228454 587850 263898
rect 587230 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 587850 228454
rect 587230 228134 587850 228218
rect 587230 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 587850 228134
rect 587230 192454 587850 227898
rect 587230 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 587850 192454
rect 587230 192134 587850 192218
rect 587230 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 587850 192134
rect 587230 156454 587850 191898
rect 587230 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 587850 156454
rect 587230 156134 587850 156218
rect 587230 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 587850 156134
rect 587230 120454 587850 155898
rect 587230 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 587850 120454
rect 587230 120134 587850 120218
rect 587230 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 587850 120134
rect 587230 84454 587850 119898
rect 587230 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 587850 84454
rect 587230 84134 587850 84218
rect 587230 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 587850 84134
rect 587230 48454 587850 83898
rect 587230 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 587850 48454
rect 587230 48134 587850 48218
rect 587230 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 587850 48134
rect 587230 12454 587850 47898
rect 587230 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 587850 12454
rect 587230 12134 587850 12218
rect 587230 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 587850 12134
rect 587230 -2266 587850 11898
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 700954 588810 707162
rect 588190 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 588810 700954
rect 588190 700634 588810 700718
rect 588190 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 588810 700634
rect 588190 664954 588810 700398
rect 588190 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 588810 664954
rect 588190 664634 588810 664718
rect 588190 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 588810 664634
rect 588190 628954 588810 664398
rect 588190 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 588810 628954
rect 588190 628634 588810 628718
rect 588190 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 588810 628634
rect 588190 592954 588810 628398
rect 588190 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 588810 592954
rect 588190 592634 588810 592718
rect 588190 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 588810 592634
rect 588190 556954 588810 592398
rect 588190 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 588810 556954
rect 588190 556634 588810 556718
rect 588190 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 588810 556634
rect 588190 520954 588810 556398
rect 588190 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 588810 520954
rect 588190 520634 588810 520718
rect 588190 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 588810 520634
rect 588190 484954 588810 520398
rect 588190 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 588810 484954
rect 588190 484634 588810 484718
rect 588190 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 588810 484634
rect 588190 448954 588810 484398
rect 588190 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 588810 448954
rect 588190 448634 588810 448718
rect 588190 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 588810 448634
rect 588190 412954 588810 448398
rect 588190 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 588810 412954
rect 588190 412634 588810 412718
rect 588190 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 588810 412634
rect 588190 376954 588810 412398
rect 588190 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 588810 376954
rect 588190 376634 588810 376718
rect 588190 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 588810 376634
rect 588190 340954 588810 376398
rect 588190 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 588810 340954
rect 588190 340634 588810 340718
rect 588190 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 588810 340634
rect 588190 304954 588810 340398
rect 588190 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 588810 304954
rect 588190 304634 588810 304718
rect 588190 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 588810 304634
rect 588190 268954 588810 304398
rect 588190 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 588810 268954
rect 588190 268634 588810 268718
rect 588190 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 588810 268634
rect 588190 232954 588810 268398
rect 588190 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 588810 232954
rect 588190 232634 588810 232718
rect 588190 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 588810 232634
rect 588190 196954 588810 232398
rect 588190 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 588810 196954
rect 588190 196634 588810 196718
rect 588190 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 588810 196634
rect 588190 160954 588810 196398
rect 588190 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 588810 160954
rect 588190 160634 588810 160718
rect 588190 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 588810 160634
rect 588190 124954 588810 160398
rect 588190 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 588810 124954
rect 588190 124634 588810 124718
rect 588190 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 588810 124634
rect 588190 88954 588810 124398
rect 588190 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 588810 88954
rect 588190 88634 588810 88718
rect 588190 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 588810 88634
rect 588190 52954 588810 88398
rect 588190 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 588810 52954
rect 588190 52634 588810 52718
rect 588190 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 588810 52634
rect 588190 16954 588810 52398
rect 588190 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 588810 16954
rect 588190 16634 588810 16718
rect 588190 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 588810 16634
rect 588190 -3226 588810 16398
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 669454 589770 708122
rect 589150 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 589770 669454
rect 589150 669134 589770 669218
rect 589150 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 589770 669134
rect 589150 633454 589770 668898
rect 589150 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 589770 633454
rect 589150 633134 589770 633218
rect 589150 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 589770 633134
rect 589150 597454 589770 632898
rect 589150 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 589770 597454
rect 589150 597134 589770 597218
rect 589150 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 589770 597134
rect 589150 561454 589770 596898
rect 589150 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 589770 561454
rect 589150 561134 589770 561218
rect 589150 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 589770 561134
rect 589150 525454 589770 560898
rect 589150 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 589770 525454
rect 589150 525134 589770 525218
rect 589150 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 589770 525134
rect 589150 489454 589770 524898
rect 589150 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 589770 489454
rect 589150 489134 589770 489218
rect 589150 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 589770 489134
rect 589150 453454 589770 488898
rect 589150 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 589770 453454
rect 589150 453134 589770 453218
rect 589150 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 589770 453134
rect 589150 417454 589770 452898
rect 589150 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 589770 417454
rect 589150 417134 589770 417218
rect 589150 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 589770 417134
rect 589150 381454 589770 416898
rect 589150 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 589770 381454
rect 589150 381134 589770 381218
rect 589150 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 589770 381134
rect 589150 345454 589770 380898
rect 589150 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 589770 345454
rect 589150 345134 589770 345218
rect 589150 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 589770 345134
rect 589150 309454 589770 344898
rect 589150 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 589770 309454
rect 589150 309134 589770 309218
rect 589150 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 589770 309134
rect 589150 273454 589770 308898
rect 589150 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 589770 273454
rect 589150 273134 589770 273218
rect 589150 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 589770 273134
rect 589150 237454 589770 272898
rect 589150 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 589770 237454
rect 589150 237134 589770 237218
rect 589150 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 589770 237134
rect 589150 201454 589770 236898
rect 589150 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 589770 201454
rect 589150 201134 589770 201218
rect 589150 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 589770 201134
rect 589150 165454 589770 200898
rect 589150 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 589770 165454
rect 589150 165134 589770 165218
rect 589150 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 589770 165134
rect 589150 129454 589770 164898
rect 589150 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 589770 129454
rect 589150 129134 589770 129218
rect 589150 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 589770 129134
rect 589150 93454 589770 128898
rect 589150 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 589770 93454
rect 589150 93134 589770 93218
rect 589150 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 589770 93134
rect 589150 57454 589770 92898
rect 589150 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 589770 57454
rect 589150 57134 589770 57218
rect 589150 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 589770 57134
rect 589150 21454 589770 56898
rect 589150 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 589770 21454
rect 589150 21134 589770 21218
rect 589150 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 589770 21134
rect 589150 -4186 589770 20898
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 673954 590730 709082
rect 590110 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 590730 673954
rect 590110 673634 590730 673718
rect 590110 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 590730 673634
rect 590110 637954 590730 673398
rect 590110 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 590730 637954
rect 590110 637634 590730 637718
rect 590110 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 590730 637634
rect 590110 601954 590730 637398
rect 590110 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 590730 601954
rect 590110 601634 590730 601718
rect 590110 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 590730 601634
rect 590110 565954 590730 601398
rect 590110 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 590730 565954
rect 590110 565634 590730 565718
rect 590110 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 590730 565634
rect 590110 529954 590730 565398
rect 590110 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 590730 529954
rect 590110 529634 590730 529718
rect 590110 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 590730 529634
rect 590110 493954 590730 529398
rect 590110 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 590730 493954
rect 590110 493634 590730 493718
rect 590110 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 590730 493634
rect 590110 457954 590730 493398
rect 590110 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 590730 457954
rect 590110 457634 590730 457718
rect 590110 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 590730 457634
rect 590110 421954 590730 457398
rect 590110 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 590730 421954
rect 590110 421634 590730 421718
rect 590110 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 590730 421634
rect 590110 385954 590730 421398
rect 590110 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 590730 385954
rect 590110 385634 590730 385718
rect 590110 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 590730 385634
rect 590110 349954 590730 385398
rect 590110 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 590730 349954
rect 590110 349634 590730 349718
rect 590110 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 590730 349634
rect 590110 313954 590730 349398
rect 590110 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 590730 313954
rect 590110 313634 590730 313718
rect 590110 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 590730 313634
rect 590110 277954 590730 313398
rect 590110 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 590730 277954
rect 590110 277634 590730 277718
rect 590110 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 590730 277634
rect 590110 241954 590730 277398
rect 590110 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 590730 241954
rect 590110 241634 590730 241718
rect 590110 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 590730 241634
rect 590110 205954 590730 241398
rect 590110 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 590730 205954
rect 590110 205634 590730 205718
rect 590110 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 590730 205634
rect 590110 169954 590730 205398
rect 590110 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 590730 169954
rect 590110 169634 590730 169718
rect 590110 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 590730 169634
rect 590110 133954 590730 169398
rect 590110 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 590730 133954
rect 590110 133634 590730 133718
rect 590110 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 590730 133634
rect 590110 97954 590730 133398
rect 590110 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 590730 97954
rect 590110 97634 590730 97718
rect 590110 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 590730 97634
rect 590110 61954 590730 97398
rect 590110 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 590730 61954
rect 590110 61634 590730 61718
rect 590110 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 590730 61634
rect 590110 25954 590730 61398
rect 590110 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 590730 25954
rect 590110 25634 590730 25718
rect 590110 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 590730 25634
rect 590110 -5146 590730 25398
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 678454 591690 710042
rect 591070 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 591690 678454
rect 591070 678134 591690 678218
rect 591070 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 591690 678134
rect 591070 642454 591690 677898
rect 591070 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 591690 642454
rect 591070 642134 591690 642218
rect 591070 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 591690 642134
rect 591070 606454 591690 641898
rect 591070 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 591690 606454
rect 591070 606134 591690 606218
rect 591070 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 591690 606134
rect 591070 570454 591690 605898
rect 591070 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 591690 570454
rect 591070 570134 591690 570218
rect 591070 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 591690 570134
rect 591070 534454 591690 569898
rect 591070 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 591690 534454
rect 591070 534134 591690 534218
rect 591070 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 591690 534134
rect 591070 498454 591690 533898
rect 591070 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 591690 498454
rect 591070 498134 591690 498218
rect 591070 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 591690 498134
rect 591070 462454 591690 497898
rect 591070 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 591690 462454
rect 591070 462134 591690 462218
rect 591070 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 591690 462134
rect 591070 426454 591690 461898
rect 591070 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 591690 426454
rect 591070 426134 591690 426218
rect 591070 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 591690 426134
rect 591070 390454 591690 425898
rect 591070 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 591690 390454
rect 591070 390134 591690 390218
rect 591070 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 591690 390134
rect 591070 354454 591690 389898
rect 591070 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 591690 354454
rect 591070 354134 591690 354218
rect 591070 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 591690 354134
rect 591070 318454 591690 353898
rect 591070 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 591690 318454
rect 591070 318134 591690 318218
rect 591070 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 591690 318134
rect 591070 282454 591690 317898
rect 591070 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 591690 282454
rect 591070 282134 591690 282218
rect 591070 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 591690 282134
rect 591070 246454 591690 281898
rect 591070 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 591690 246454
rect 591070 246134 591690 246218
rect 591070 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 591690 246134
rect 591070 210454 591690 245898
rect 591070 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 591690 210454
rect 591070 210134 591690 210218
rect 591070 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 591690 210134
rect 591070 174454 591690 209898
rect 591070 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 591690 174454
rect 591070 174134 591690 174218
rect 591070 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 591690 174134
rect 591070 138454 591690 173898
rect 591070 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 591690 138454
rect 591070 138134 591690 138218
rect 591070 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 591690 138134
rect 591070 102454 591690 137898
rect 591070 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 591690 102454
rect 591070 102134 591690 102218
rect 591070 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 591690 102134
rect 591070 66454 591690 101898
rect 591070 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 591690 66454
rect 591070 66134 591690 66218
rect 591070 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 591690 66134
rect 591070 30454 591690 65898
rect 591070 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 591690 30454
rect 591070 30134 591690 30218
rect 591070 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 591690 30134
rect 591070 -6106 591690 29898
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 682954 592650 711002
rect 592030 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect 592030 682634 592650 682718
rect 592030 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect 592030 646954 592650 682398
rect 592030 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect 592030 646634 592650 646718
rect 592030 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect 592030 610954 592650 646398
rect 592030 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect 592030 610634 592650 610718
rect 592030 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect 592030 574954 592650 610398
rect 592030 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect 592030 574634 592650 574718
rect 592030 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect 592030 538954 592650 574398
rect 592030 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect 592030 538634 592650 538718
rect 592030 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect 592030 502954 592650 538398
rect 592030 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect 592030 502634 592650 502718
rect 592030 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect 592030 466954 592650 502398
rect 592030 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect 592030 466634 592650 466718
rect 592030 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect 592030 430954 592650 466398
rect 592030 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect 592030 430634 592650 430718
rect 592030 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect 592030 394954 592650 430398
rect 592030 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect 592030 394634 592650 394718
rect 592030 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect 592030 358954 592650 394398
rect 592030 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect 592030 358634 592650 358718
rect 592030 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect 592030 322954 592650 358398
rect 592030 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect 592030 322634 592650 322718
rect 592030 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect 592030 286954 592650 322398
rect 592030 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect 592030 286634 592650 286718
rect 592030 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect 592030 250954 592650 286398
rect 592030 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect 592030 250634 592650 250718
rect 592030 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect 592030 214954 592650 250398
rect 592030 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect 592030 214634 592650 214718
rect 592030 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect 592030 178954 592650 214398
rect 592030 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect 592030 178634 592650 178718
rect 592030 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect 592030 142954 592650 178398
rect 592030 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect 592030 142634 592650 142718
rect 592030 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect 592030 106954 592650 142398
rect 592030 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect 592030 106634 592650 106718
rect 592030 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect 592030 70954 592650 106398
rect 592030 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect 592030 70634 592650 70718
rect 592030 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect 592030 34954 592650 70398
rect 592030 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect 592030 34634 592650 34718
rect 592030 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect 592030 -7066 592650 34398
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 682718 -8458 682954
rect -8374 682718 -8138 682954
rect -8694 682398 -8458 682634
rect -8374 682398 -8138 682634
rect -8694 646718 -8458 646954
rect -8374 646718 -8138 646954
rect -8694 646398 -8458 646634
rect -8374 646398 -8138 646634
rect -8694 610718 -8458 610954
rect -8374 610718 -8138 610954
rect -8694 610398 -8458 610634
rect -8374 610398 -8138 610634
rect -8694 574718 -8458 574954
rect -8374 574718 -8138 574954
rect -8694 574398 -8458 574634
rect -8374 574398 -8138 574634
rect -8694 538718 -8458 538954
rect -8374 538718 -8138 538954
rect -8694 538398 -8458 538634
rect -8374 538398 -8138 538634
rect -8694 502718 -8458 502954
rect -8374 502718 -8138 502954
rect -8694 502398 -8458 502634
rect -8374 502398 -8138 502634
rect -8694 466718 -8458 466954
rect -8374 466718 -8138 466954
rect -8694 466398 -8458 466634
rect -8374 466398 -8138 466634
rect -8694 430718 -8458 430954
rect -8374 430718 -8138 430954
rect -8694 430398 -8458 430634
rect -8374 430398 -8138 430634
rect -8694 394718 -8458 394954
rect -8374 394718 -8138 394954
rect -8694 394398 -8458 394634
rect -8374 394398 -8138 394634
rect -8694 358718 -8458 358954
rect -8374 358718 -8138 358954
rect -8694 358398 -8458 358634
rect -8374 358398 -8138 358634
rect -8694 322718 -8458 322954
rect -8374 322718 -8138 322954
rect -8694 322398 -8458 322634
rect -8374 322398 -8138 322634
rect -8694 286718 -8458 286954
rect -8374 286718 -8138 286954
rect -8694 286398 -8458 286634
rect -8374 286398 -8138 286634
rect -8694 250718 -8458 250954
rect -8374 250718 -8138 250954
rect -8694 250398 -8458 250634
rect -8374 250398 -8138 250634
rect -8694 214718 -8458 214954
rect -8374 214718 -8138 214954
rect -8694 214398 -8458 214634
rect -8374 214398 -8138 214634
rect -8694 178718 -8458 178954
rect -8374 178718 -8138 178954
rect -8694 178398 -8458 178634
rect -8374 178398 -8138 178634
rect -8694 142718 -8458 142954
rect -8374 142718 -8138 142954
rect -8694 142398 -8458 142634
rect -8374 142398 -8138 142634
rect -8694 106718 -8458 106954
rect -8374 106718 -8138 106954
rect -8694 106398 -8458 106634
rect -8374 106398 -8138 106634
rect -8694 70718 -8458 70954
rect -8374 70718 -8138 70954
rect -8694 70398 -8458 70634
rect -8374 70398 -8138 70634
rect -8694 34718 -8458 34954
rect -8374 34718 -8138 34954
rect -8694 34398 -8458 34634
rect -8374 34398 -8138 34634
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 678218 -7498 678454
rect -7414 678218 -7178 678454
rect -7734 677898 -7498 678134
rect -7414 677898 -7178 678134
rect -7734 642218 -7498 642454
rect -7414 642218 -7178 642454
rect -7734 641898 -7498 642134
rect -7414 641898 -7178 642134
rect -7734 606218 -7498 606454
rect -7414 606218 -7178 606454
rect -7734 605898 -7498 606134
rect -7414 605898 -7178 606134
rect -7734 570218 -7498 570454
rect -7414 570218 -7178 570454
rect -7734 569898 -7498 570134
rect -7414 569898 -7178 570134
rect -7734 534218 -7498 534454
rect -7414 534218 -7178 534454
rect -7734 533898 -7498 534134
rect -7414 533898 -7178 534134
rect -7734 498218 -7498 498454
rect -7414 498218 -7178 498454
rect -7734 497898 -7498 498134
rect -7414 497898 -7178 498134
rect -7734 462218 -7498 462454
rect -7414 462218 -7178 462454
rect -7734 461898 -7498 462134
rect -7414 461898 -7178 462134
rect -7734 426218 -7498 426454
rect -7414 426218 -7178 426454
rect -7734 425898 -7498 426134
rect -7414 425898 -7178 426134
rect -7734 390218 -7498 390454
rect -7414 390218 -7178 390454
rect -7734 389898 -7498 390134
rect -7414 389898 -7178 390134
rect -7734 354218 -7498 354454
rect -7414 354218 -7178 354454
rect -7734 353898 -7498 354134
rect -7414 353898 -7178 354134
rect -7734 318218 -7498 318454
rect -7414 318218 -7178 318454
rect -7734 317898 -7498 318134
rect -7414 317898 -7178 318134
rect -7734 282218 -7498 282454
rect -7414 282218 -7178 282454
rect -7734 281898 -7498 282134
rect -7414 281898 -7178 282134
rect -7734 246218 -7498 246454
rect -7414 246218 -7178 246454
rect -7734 245898 -7498 246134
rect -7414 245898 -7178 246134
rect -7734 210218 -7498 210454
rect -7414 210218 -7178 210454
rect -7734 209898 -7498 210134
rect -7414 209898 -7178 210134
rect -7734 174218 -7498 174454
rect -7414 174218 -7178 174454
rect -7734 173898 -7498 174134
rect -7414 173898 -7178 174134
rect -7734 138218 -7498 138454
rect -7414 138218 -7178 138454
rect -7734 137898 -7498 138134
rect -7414 137898 -7178 138134
rect -7734 102218 -7498 102454
rect -7414 102218 -7178 102454
rect -7734 101898 -7498 102134
rect -7414 101898 -7178 102134
rect -7734 66218 -7498 66454
rect -7414 66218 -7178 66454
rect -7734 65898 -7498 66134
rect -7414 65898 -7178 66134
rect -7734 30218 -7498 30454
rect -7414 30218 -7178 30454
rect -7734 29898 -7498 30134
rect -7414 29898 -7178 30134
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 673718 -6538 673954
rect -6454 673718 -6218 673954
rect -6774 673398 -6538 673634
rect -6454 673398 -6218 673634
rect -6774 637718 -6538 637954
rect -6454 637718 -6218 637954
rect -6774 637398 -6538 637634
rect -6454 637398 -6218 637634
rect -6774 601718 -6538 601954
rect -6454 601718 -6218 601954
rect -6774 601398 -6538 601634
rect -6454 601398 -6218 601634
rect -6774 565718 -6538 565954
rect -6454 565718 -6218 565954
rect -6774 565398 -6538 565634
rect -6454 565398 -6218 565634
rect -6774 529718 -6538 529954
rect -6454 529718 -6218 529954
rect -6774 529398 -6538 529634
rect -6454 529398 -6218 529634
rect -6774 493718 -6538 493954
rect -6454 493718 -6218 493954
rect -6774 493398 -6538 493634
rect -6454 493398 -6218 493634
rect -6774 457718 -6538 457954
rect -6454 457718 -6218 457954
rect -6774 457398 -6538 457634
rect -6454 457398 -6218 457634
rect -6774 421718 -6538 421954
rect -6454 421718 -6218 421954
rect -6774 421398 -6538 421634
rect -6454 421398 -6218 421634
rect -6774 385718 -6538 385954
rect -6454 385718 -6218 385954
rect -6774 385398 -6538 385634
rect -6454 385398 -6218 385634
rect -6774 349718 -6538 349954
rect -6454 349718 -6218 349954
rect -6774 349398 -6538 349634
rect -6454 349398 -6218 349634
rect -6774 313718 -6538 313954
rect -6454 313718 -6218 313954
rect -6774 313398 -6538 313634
rect -6454 313398 -6218 313634
rect -6774 277718 -6538 277954
rect -6454 277718 -6218 277954
rect -6774 277398 -6538 277634
rect -6454 277398 -6218 277634
rect -6774 241718 -6538 241954
rect -6454 241718 -6218 241954
rect -6774 241398 -6538 241634
rect -6454 241398 -6218 241634
rect -6774 205718 -6538 205954
rect -6454 205718 -6218 205954
rect -6774 205398 -6538 205634
rect -6454 205398 -6218 205634
rect -6774 169718 -6538 169954
rect -6454 169718 -6218 169954
rect -6774 169398 -6538 169634
rect -6454 169398 -6218 169634
rect -6774 133718 -6538 133954
rect -6454 133718 -6218 133954
rect -6774 133398 -6538 133634
rect -6454 133398 -6218 133634
rect -6774 97718 -6538 97954
rect -6454 97718 -6218 97954
rect -6774 97398 -6538 97634
rect -6454 97398 -6218 97634
rect -6774 61718 -6538 61954
rect -6454 61718 -6218 61954
rect -6774 61398 -6538 61634
rect -6454 61398 -6218 61634
rect -6774 25718 -6538 25954
rect -6454 25718 -6218 25954
rect -6774 25398 -6538 25634
rect -6454 25398 -6218 25634
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 669218 -5578 669454
rect -5494 669218 -5258 669454
rect -5814 668898 -5578 669134
rect -5494 668898 -5258 669134
rect -5814 633218 -5578 633454
rect -5494 633218 -5258 633454
rect -5814 632898 -5578 633134
rect -5494 632898 -5258 633134
rect -5814 597218 -5578 597454
rect -5494 597218 -5258 597454
rect -5814 596898 -5578 597134
rect -5494 596898 -5258 597134
rect -5814 561218 -5578 561454
rect -5494 561218 -5258 561454
rect -5814 560898 -5578 561134
rect -5494 560898 -5258 561134
rect -5814 525218 -5578 525454
rect -5494 525218 -5258 525454
rect -5814 524898 -5578 525134
rect -5494 524898 -5258 525134
rect -5814 489218 -5578 489454
rect -5494 489218 -5258 489454
rect -5814 488898 -5578 489134
rect -5494 488898 -5258 489134
rect -5814 453218 -5578 453454
rect -5494 453218 -5258 453454
rect -5814 452898 -5578 453134
rect -5494 452898 -5258 453134
rect -5814 417218 -5578 417454
rect -5494 417218 -5258 417454
rect -5814 416898 -5578 417134
rect -5494 416898 -5258 417134
rect -5814 381218 -5578 381454
rect -5494 381218 -5258 381454
rect -5814 380898 -5578 381134
rect -5494 380898 -5258 381134
rect -5814 345218 -5578 345454
rect -5494 345218 -5258 345454
rect -5814 344898 -5578 345134
rect -5494 344898 -5258 345134
rect -5814 309218 -5578 309454
rect -5494 309218 -5258 309454
rect -5814 308898 -5578 309134
rect -5494 308898 -5258 309134
rect -5814 273218 -5578 273454
rect -5494 273218 -5258 273454
rect -5814 272898 -5578 273134
rect -5494 272898 -5258 273134
rect -5814 237218 -5578 237454
rect -5494 237218 -5258 237454
rect -5814 236898 -5578 237134
rect -5494 236898 -5258 237134
rect -5814 201218 -5578 201454
rect -5494 201218 -5258 201454
rect -5814 200898 -5578 201134
rect -5494 200898 -5258 201134
rect -5814 165218 -5578 165454
rect -5494 165218 -5258 165454
rect -5814 164898 -5578 165134
rect -5494 164898 -5258 165134
rect -5814 129218 -5578 129454
rect -5494 129218 -5258 129454
rect -5814 128898 -5578 129134
rect -5494 128898 -5258 129134
rect -5814 93218 -5578 93454
rect -5494 93218 -5258 93454
rect -5814 92898 -5578 93134
rect -5494 92898 -5258 93134
rect -5814 57218 -5578 57454
rect -5494 57218 -5258 57454
rect -5814 56898 -5578 57134
rect -5494 56898 -5258 57134
rect -5814 21218 -5578 21454
rect -5494 21218 -5258 21454
rect -5814 20898 -5578 21134
rect -5494 20898 -5258 21134
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 700718 -4618 700954
rect -4534 700718 -4298 700954
rect -4854 700398 -4618 700634
rect -4534 700398 -4298 700634
rect -4854 664718 -4618 664954
rect -4534 664718 -4298 664954
rect -4854 664398 -4618 664634
rect -4534 664398 -4298 664634
rect -4854 628718 -4618 628954
rect -4534 628718 -4298 628954
rect -4854 628398 -4618 628634
rect -4534 628398 -4298 628634
rect -4854 592718 -4618 592954
rect -4534 592718 -4298 592954
rect -4854 592398 -4618 592634
rect -4534 592398 -4298 592634
rect -4854 556718 -4618 556954
rect -4534 556718 -4298 556954
rect -4854 556398 -4618 556634
rect -4534 556398 -4298 556634
rect -4854 520718 -4618 520954
rect -4534 520718 -4298 520954
rect -4854 520398 -4618 520634
rect -4534 520398 -4298 520634
rect -4854 484718 -4618 484954
rect -4534 484718 -4298 484954
rect -4854 484398 -4618 484634
rect -4534 484398 -4298 484634
rect -4854 448718 -4618 448954
rect -4534 448718 -4298 448954
rect -4854 448398 -4618 448634
rect -4534 448398 -4298 448634
rect -4854 412718 -4618 412954
rect -4534 412718 -4298 412954
rect -4854 412398 -4618 412634
rect -4534 412398 -4298 412634
rect -4854 376718 -4618 376954
rect -4534 376718 -4298 376954
rect -4854 376398 -4618 376634
rect -4534 376398 -4298 376634
rect -4854 340718 -4618 340954
rect -4534 340718 -4298 340954
rect -4854 340398 -4618 340634
rect -4534 340398 -4298 340634
rect -4854 304718 -4618 304954
rect -4534 304718 -4298 304954
rect -4854 304398 -4618 304634
rect -4534 304398 -4298 304634
rect -4854 268718 -4618 268954
rect -4534 268718 -4298 268954
rect -4854 268398 -4618 268634
rect -4534 268398 -4298 268634
rect -4854 232718 -4618 232954
rect -4534 232718 -4298 232954
rect -4854 232398 -4618 232634
rect -4534 232398 -4298 232634
rect -4854 196718 -4618 196954
rect -4534 196718 -4298 196954
rect -4854 196398 -4618 196634
rect -4534 196398 -4298 196634
rect -4854 160718 -4618 160954
rect -4534 160718 -4298 160954
rect -4854 160398 -4618 160634
rect -4534 160398 -4298 160634
rect -4854 124718 -4618 124954
rect -4534 124718 -4298 124954
rect -4854 124398 -4618 124634
rect -4534 124398 -4298 124634
rect -4854 88718 -4618 88954
rect -4534 88718 -4298 88954
rect -4854 88398 -4618 88634
rect -4534 88398 -4298 88634
rect -4854 52718 -4618 52954
rect -4534 52718 -4298 52954
rect -4854 52398 -4618 52634
rect -4534 52398 -4298 52634
rect -4854 16718 -4618 16954
rect -4534 16718 -4298 16954
rect -4854 16398 -4618 16634
rect -4534 16398 -4298 16634
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 696218 -3658 696454
rect -3574 696218 -3338 696454
rect -3894 695898 -3658 696134
rect -3574 695898 -3338 696134
rect -3894 660218 -3658 660454
rect -3574 660218 -3338 660454
rect -3894 659898 -3658 660134
rect -3574 659898 -3338 660134
rect -3894 624218 -3658 624454
rect -3574 624218 -3338 624454
rect -3894 623898 -3658 624134
rect -3574 623898 -3338 624134
rect -3894 588218 -3658 588454
rect -3574 588218 -3338 588454
rect -3894 587898 -3658 588134
rect -3574 587898 -3338 588134
rect -3894 552218 -3658 552454
rect -3574 552218 -3338 552454
rect -3894 551898 -3658 552134
rect -3574 551898 -3338 552134
rect -3894 516218 -3658 516454
rect -3574 516218 -3338 516454
rect -3894 515898 -3658 516134
rect -3574 515898 -3338 516134
rect -3894 480218 -3658 480454
rect -3574 480218 -3338 480454
rect -3894 479898 -3658 480134
rect -3574 479898 -3338 480134
rect -3894 444218 -3658 444454
rect -3574 444218 -3338 444454
rect -3894 443898 -3658 444134
rect -3574 443898 -3338 444134
rect -3894 408218 -3658 408454
rect -3574 408218 -3338 408454
rect -3894 407898 -3658 408134
rect -3574 407898 -3338 408134
rect -3894 372218 -3658 372454
rect -3574 372218 -3338 372454
rect -3894 371898 -3658 372134
rect -3574 371898 -3338 372134
rect -3894 336218 -3658 336454
rect -3574 336218 -3338 336454
rect -3894 335898 -3658 336134
rect -3574 335898 -3338 336134
rect -3894 300218 -3658 300454
rect -3574 300218 -3338 300454
rect -3894 299898 -3658 300134
rect -3574 299898 -3338 300134
rect -3894 264218 -3658 264454
rect -3574 264218 -3338 264454
rect -3894 263898 -3658 264134
rect -3574 263898 -3338 264134
rect -3894 228218 -3658 228454
rect -3574 228218 -3338 228454
rect -3894 227898 -3658 228134
rect -3574 227898 -3338 228134
rect -3894 192218 -3658 192454
rect -3574 192218 -3338 192454
rect -3894 191898 -3658 192134
rect -3574 191898 -3338 192134
rect -3894 156218 -3658 156454
rect -3574 156218 -3338 156454
rect -3894 155898 -3658 156134
rect -3574 155898 -3338 156134
rect -3894 120218 -3658 120454
rect -3574 120218 -3338 120454
rect -3894 119898 -3658 120134
rect -3574 119898 -3338 120134
rect -3894 84218 -3658 84454
rect -3574 84218 -3338 84454
rect -3894 83898 -3658 84134
rect -3574 83898 -3338 84134
rect -3894 48218 -3658 48454
rect -3574 48218 -3338 48454
rect -3894 47898 -3658 48134
rect -3574 47898 -3338 48134
rect -3894 12218 -3658 12454
rect -3574 12218 -3338 12454
rect -3894 11898 -3658 12134
rect -3574 11898 -3338 12134
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 691718 -2698 691954
rect -2614 691718 -2378 691954
rect -2934 691398 -2698 691634
rect -2614 691398 -2378 691634
rect -2934 655718 -2698 655954
rect -2614 655718 -2378 655954
rect -2934 655398 -2698 655634
rect -2614 655398 -2378 655634
rect -2934 619718 -2698 619954
rect -2614 619718 -2378 619954
rect -2934 619398 -2698 619634
rect -2614 619398 -2378 619634
rect -2934 583718 -2698 583954
rect -2614 583718 -2378 583954
rect -2934 583398 -2698 583634
rect -2614 583398 -2378 583634
rect -2934 547718 -2698 547954
rect -2614 547718 -2378 547954
rect -2934 547398 -2698 547634
rect -2614 547398 -2378 547634
rect -2934 511718 -2698 511954
rect -2614 511718 -2378 511954
rect -2934 511398 -2698 511634
rect -2614 511398 -2378 511634
rect -2934 475718 -2698 475954
rect -2614 475718 -2378 475954
rect -2934 475398 -2698 475634
rect -2614 475398 -2378 475634
rect -2934 439718 -2698 439954
rect -2614 439718 -2378 439954
rect -2934 439398 -2698 439634
rect -2614 439398 -2378 439634
rect -2934 403718 -2698 403954
rect -2614 403718 -2378 403954
rect -2934 403398 -2698 403634
rect -2614 403398 -2378 403634
rect -2934 367718 -2698 367954
rect -2614 367718 -2378 367954
rect -2934 367398 -2698 367634
rect -2614 367398 -2378 367634
rect -2934 331718 -2698 331954
rect -2614 331718 -2378 331954
rect -2934 331398 -2698 331634
rect -2614 331398 -2378 331634
rect -2934 295718 -2698 295954
rect -2614 295718 -2378 295954
rect -2934 295398 -2698 295634
rect -2614 295398 -2378 295634
rect -2934 259718 -2698 259954
rect -2614 259718 -2378 259954
rect -2934 259398 -2698 259634
rect -2614 259398 -2378 259634
rect -2934 223718 -2698 223954
rect -2614 223718 -2378 223954
rect -2934 223398 -2698 223634
rect -2614 223398 -2378 223634
rect -2934 187718 -2698 187954
rect -2614 187718 -2378 187954
rect -2934 187398 -2698 187634
rect -2614 187398 -2378 187634
rect -2934 151718 -2698 151954
rect -2614 151718 -2378 151954
rect -2934 151398 -2698 151634
rect -2614 151398 -2378 151634
rect -2934 115718 -2698 115954
rect -2614 115718 -2378 115954
rect -2934 115398 -2698 115634
rect -2614 115398 -2378 115634
rect -2934 79718 -2698 79954
rect -2614 79718 -2378 79954
rect -2934 79398 -2698 79634
rect -2614 79398 -2378 79634
rect -2934 43718 -2698 43954
rect -2614 43718 -2378 43954
rect -2934 43398 -2698 43634
rect -2614 43398 -2378 43634
rect -2934 7718 -2698 7954
rect -2614 7718 -2378 7954
rect -2934 7398 -2698 7634
rect -2614 7398 -2378 7634
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 6326 705562 6562 705798
rect 6646 705562 6882 705798
rect 6326 705242 6562 705478
rect 6646 705242 6882 705478
rect 6326 691718 6562 691954
rect 6646 691718 6882 691954
rect 6326 691398 6562 691634
rect 6646 691398 6882 691634
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 6326 655718 6562 655954
rect 6646 655718 6882 655954
rect 6326 655398 6562 655634
rect 6646 655398 6882 655634
rect 6326 619718 6562 619954
rect 6646 619718 6882 619954
rect 6326 619398 6562 619634
rect 6646 619398 6882 619634
rect 6326 583718 6562 583954
rect 6646 583718 6882 583954
rect 6326 583398 6562 583634
rect 6646 583398 6882 583634
rect 6326 547718 6562 547954
rect 6646 547718 6882 547954
rect 6326 547398 6562 547634
rect 6646 547398 6882 547634
rect 6326 511718 6562 511954
rect 6646 511718 6882 511954
rect 6326 511398 6562 511634
rect 6646 511398 6882 511634
rect 6326 475718 6562 475954
rect 6646 475718 6882 475954
rect 6326 475398 6562 475634
rect 6646 475398 6882 475634
rect 6326 439718 6562 439954
rect 6646 439718 6882 439954
rect 6326 439398 6562 439634
rect 6646 439398 6882 439634
rect 6326 403718 6562 403954
rect 6646 403718 6882 403954
rect 6326 403398 6562 403634
rect 6646 403398 6882 403634
rect 6326 367718 6562 367954
rect 6646 367718 6882 367954
rect 6326 367398 6562 367634
rect 6646 367398 6882 367634
rect 6326 331718 6562 331954
rect 6646 331718 6882 331954
rect 6326 331398 6562 331634
rect 6646 331398 6882 331634
rect 6326 295718 6562 295954
rect 6646 295718 6882 295954
rect 6326 295398 6562 295634
rect 6646 295398 6882 295634
rect 6326 259718 6562 259954
rect 6646 259718 6882 259954
rect 6326 259398 6562 259634
rect 6646 259398 6882 259634
rect 6326 223718 6562 223954
rect 6646 223718 6882 223954
rect 6326 223398 6562 223634
rect 6646 223398 6882 223634
rect 6326 187718 6562 187954
rect 6646 187718 6882 187954
rect 6326 187398 6562 187634
rect 6646 187398 6882 187634
rect 6326 151718 6562 151954
rect 6646 151718 6882 151954
rect 6326 151398 6562 151634
rect 6646 151398 6882 151634
rect 6326 115718 6562 115954
rect 6646 115718 6882 115954
rect 6326 115398 6562 115634
rect 6646 115398 6882 115634
rect 6326 79718 6562 79954
rect 6646 79718 6882 79954
rect 6326 79398 6562 79634
rect 6646 79398 6882 79634
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 6326 43718 6562 43954
rect 6646 43718 6882 43954
rect 6326 43398 6562 43634
rect 6646 43398 6882 43634
rect 6326 7718 6562 7954
rect 6646 7718 6882 7954
rect 6326 7398 6562 7634
rect 6646 7398 6882 7634
rect 6326 -1542 6562 -1306
rect 6646 -1542 6882 -1306
rect 6326 -1862 6562 -1626
rect 6646 -1862 6882 -1626
rect 10826 706522 11062 706758
rect 11146 706522 11382 706758
rect 10826 706202 11062 706438
rect 11146 706202 11382 706438
rect 10826 696218 11062 696454
rect 11146 696218 11382 696454
rect 10826 695898 11062 696134
rect 11146 695898 11382 696134
rect 10826 660218 11062 660454
rect 11146 660218 11382 660454
rect 10826 659898 11062 660134
rect 11146 659898 11382 660134
rect 10826 624218 11062 624454
rect 11146 624218 11382 624454
rect 10826 623898 11062 624134
rect 11146 623898 11382 624134
rect 10826 588218 11062 588454
rect 11146 588218 11382 588454
rect 10826 587898 11062 588134
rect 11146 587898 11382 588134
rect 10826 552218 11062 552454
rect 11146 552218 11382 552454
rect 10826 551898 11062 552134
rect 11146 551898 11382 552134
rect 10826 516218 11062 516454
rect 11146 516218 11382 516454
rect 10826 515898 11062 516134
rect 11146 515898 11382 516134
rect 10826 480218 11062 480454
rect 11146 480218 11382 480454
rect 10826 479898 11062 480134
rect 11146 479898 11382 480134
rect 10826 444218 11062 444454
rect 11146 444218 11382 444454
rect 10826 443898 11062 444134
rect 11146 443898 11382 444134
rect 10826 408218 11062 408454
rect 11146 408218 11382 408454
rect 10826 407898 11062 408134
rect 11146 407898 11382 408134
rect 10826 372218 11062 372454
rect 11146 372218 11382 372454
rect 10826 371898 11062 372134
rect 11146 371898 11382 372134
rect 10826 336218 11062 336454
rect 11146 336218 11382 336454
rect 10826 335898 11062 336134
rect 11146 335898 11382 336134
rect 10826 300218 11062 300454
rect 11146 300218 11382 300454
rect 10826 299898 11062 300134
rect 11146 299898 11382 300134
rect 10826 264218 11062 264454
rect 11146 264218 11382 264454
rect 10826 263898 11062 264134
rect 11146 263898 11382 264134
rect 10826 228218 11062 228454
rect 11146 228218 11382 228454
rect 10826 227898 11062 228134
rect 11146 227898 11382 228134
rect 10826 192218 11062 192454
rect 11146 192218 11382 192454
rect 10826 191898 11062 192134
rect 11146 191898 11382 192134
rect 10826 156218 11062 156454
rect 11146 156218 11382 156454
rect 10826 155898 11062 156134
rect 11146 155898 11382 156134
rect 10826 120218 11062 120454
rect 11146 120218 11382 120454
rect 10826 119898 11062 120134
rect 11146 119898 11382 120134
rect 10826 84218 11062 84454
rect 11146 84218 11382 84454
rect 10826 83898 11062 84134
rect 11146 83898 11382 84134
rect 10826 48218 11062 48454
rect 11146 48218 11382 48454
rect 10826 47898 11062 48134
rect 11146 47898 11382 48134
rect 10826 12218 11062 12454
rect 11146 12218 11382 12454
rect 10826 11898 11062 12134
rect 11146 11898 11382 12134
rect 10826 -2502 11062 -2266
rect 11146 -2502 11382 -2266
rect 10826 -2822 11062 -2586
rect 11146 -2822 11382 -2586
rect 15326 707482 15562 707718
rect 15646 707482 15882 707718
rect 15326 707162 15562 707398
rect 15646 707162 15882 707398
rect 15326 700718 15562 700954
rect 15646 700718 15882 700954
rect 15326 700398 15562 700634
rect 15646 700398 15882 700634
rect 15326 664718 15562 664954
rect 15646 664718 15882 664954
rect 15326 664398 15562 664634
rect 15646 664398 15882 664634
rect 15326 628718 15562 628954
rect 15646 628718 15882 628954
rect 15326 628398 15562 628634
rect 15646 628398 15882 628634
rect 15326 592718 15562 592954
rect 15646 592718 15882 592954
rect 15326 592398 15562 592634
rect 15646 592398 15882 592634
rect 15326 556718 15562 556954
rect 15646 556718 15882 556954
rect 15326 556398 15562 556634
rect 15646 556398 15882 556634
rect 15326 520718 15562 520954
rect 15646 520718 15882 520954
rect 15326 520398 15562 520634
rect 15646 520398 15882 520634
rect 15326 484718 15562 484954
rect 15646 484718 15882 484954
rect 15326 484398 15562 484634
rect 15646 484398 15882 484634
rect 15326 448718 15562 448954
rect 15646 448718 15882 448954
rect 15326 448398 15562 448634
rect 15646 448398 15882 448634
rect 15326 412718 15562 412954
rect 15646 412718 15882 412954
rect 15326 412398 15562 412634
rect 15646 412398 15882 412634
rect 15326 376718 15562 376954
rect 15646 376718 15882 376954
rect 15326 376398 15562 376634
rect 15646 376398 15882 376634
rect 15326 340718 15562 340954
rect 15646 340718 15882 340954
rect 15326 340398 15562 340634
rect 15646 340398 15882 340634
rect 15326 304718 15562 304954
rect 15646 304718 15882 304954
rect 15326 304398 15562 304634
rect 15646 304398 15882 304634
rect 15326 268718 15562 268954
rect 15646 268718 15882 268954
rect 15326 268398 15562 268634
rect 15646 268398 15882 268634
rect 15326 232718 15562 232954
rect 15646 232718 15882 232954
rect 15326 232398 15562 232634
rect 15646 232398 15882 232634
rect 15326 196718 15562 196954
rect 15646 196718 15882 196954
rect 15326 196398 15562 196634
rect 15646 196398 15882 196634
rect 15326 160718 15562 160954
rect 15646 160718 15882 160954
rect 15326 160398 15562 160634
rect 15646 160398 15882 160634
rect 15326 124718 15562 124954
rect 15646 124718 15882 124954
rect 15326 124398 15562 124634
rect 15646 124398 15882 124634
rect 15326 88718 15562 88954
rect 15646 88718 15882 88954
rect 15326 88398 15562 88634
rect 15646 88398 15882 88634
rect 15326 52718 15562 52954
rect 15646 52718 15882 52954
rect 15326 52398 15562 52634
rect 15646 52398 15882 52634
rect 15326 16718 15562 16954
rect 15646 16718 15882 16954
rect 15326 16398 15562 16634
rect 15646 16398 15882 16634
rect 15326 -3462 15562 -3226
rect 15646 -3462 15882 -3226
rect 15326 -3782 15562 -3546
rect 15646 -3782 15882 -3546
rect 19826 708442 20062 708678
rect 20146 708442 20382 708678
rect 19826 708122 20062 708358
rect 20146 708122 20382 708358
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -4422 20062 -4186
rect 20146 -4422 20382 -4186
rect 19826 -4742 20062 -4506
rect 20146 -4742 20382 -4506
rect 24326 709402 24562 709638
rect 24646 709402 24882 709638
rect 24326 709082 24562 709318
rect 24646 709082 24882 709318
rect 24326 673718 24562 673954
rect 24646 673718 24882 673954
rect 24326 673398 24562 673634
rect 24646 673398 24882 673634
rect 24326 637718 24562 637954
rect 24646 637718 24882 637954
rect 24326 637398 24562 637634
rect 24646 637398 24882 637634
rect 24326 601718 24562 601954
rect 24646 601718 24882 601954
rect 24326 601398 24562 601634
rect 24646 601398 24882 601634
rect 24326 565718 24562 565954
rect 24646 565718 24882 565954
rect 24326 565398 24562 565634
rect 24646 565398 24882 565634
rect 24326 529718 24562 529954
rect 24646 529718 24882 529954
rect 24326 529398 24562 529634
rect 24646 529398 24882 529634
rect 24326 493718 24562 493954
rect 24646 493718 24882 493954
rect 24326 493398 24562 493634
rect 24646 493398 24882 493634
rect 24326 457718 24562 457954
rect 24646 457718 24882 457954
rect 24326 457398 24562 457634
rect 24646 457398 24882 457634
rect 24326 421718 24562 421954
rect 24646 421718 24882 421954
rect 24326 421398 24562 421634
rect 24646 421398 24882 421634
rect 24326 385718 24562 385954
rect 24646 385718 24882 385954
rect 24326 385398 24562 385634
rect 24646 385398 24882 385634
rect 24326 349718 24562 349954
rect 24646 349718 24882 349954
rect 24326 349398 24562 349634
rect 24646 349398 24882 349634
rect 24326 313718 24562 313954
rect 24646 313718 24882 313954
rect 24326 313398 24562 313634
rect 24646 313398 24882 313634
rect 24326 277718 24562 277954
rect 24646 277718 24882 277954
rect 24326 277398 24562 277634
rect 24646 277398 24882 277634
rect 24326 241718 24562 241954
rect 24646 241718 24882 241954
rect 24326 241398 24562 241634
rect 24646 241398 24882 241634
rect 24326 205718 24562 205954
rect 24646 205718 24882 205954
rect 24326 205398 24562 205634
rect 24646 205398 24882 205634
rect 24326 169718 24562 169954
rect 24646 169718 24882 169954
rect 24326 169398 24562 169634
rect 24646 169398 24882 169634
rect 24326 133718 24562 133954
rect 24646 133718 24882 133954
rect 24326 133398 24562 133634
rect 24646 133398 24882 133634
rect 24326 97718 24562 97954
rect 24646 97718 24882 97954
rect 24326 97398 24562 97634
rect 24646 97398 24882 97634
rect 24326 61718 24562 61954
rect 24646 61718 24882 61954
rect 24326 61398 24562 61634
rect 24646 61398 24882 61634
rect 24326 25718 24562 25954
rect 24646 25718 24882 25954
rect 24326 25398 24562 25634
rect 24646 25398 24882 25634
rect 24326 -5382 24562 -5146
rect 24646 -5382 24882 -5146
rect 24326 -5702 24562 -5466
rect 24646 -5702 24882 -5466
rect 28826 710362 29062 710598
rect 29146 710362 29382 710598
rect 28826 710042 29062 710278
rect 29146 710042 29382 710278
rect 28826 678218 29062 678454
rect 29146 678218 29382 678454
rect 28826 677898 29062 678134
rect 29146 677898 29382 678134
rect 28826 642218 29062 642454
rect 29146 642218 29382 642454
rect 28826 641898 29062 642134
rect 29146 641898 29382 642134
rect 28826 606218 29062 606454
rect 29146 606218 29382 606454
rect 28826 605898 29062 606134
rect 29146 605898 29382 606134
rect 28826 570218 29062 570454
rect 29146 570218 29382 570454
rect 28826 569898 29062 570134
rect 29146 569898 29382 570134
rect 28826 534218 29062 534454
rect 29146 534218 29382 534454
rect 28826 533898 29062 534134
rect 29146 533898 29382 534134
rect 28826 498218 29062 498454
rect 29146 498218 29382 498454
rect 28826 497898 29062 498134
rect 29146 497898 29382 498134
rect 28826 462218 29062 462454
rect 29146 462218 29382 462454
rect 28826 461898 29062 462134
rect 29146 461898 29382 462134
rect 28826 426218 29062 426454
rect 29146 426218 29382 426454
rect 28826 425898 29062 426134
rect 29146 425898 29382 426134
rect 28826 390218 29062 390454
rect 29146 390218 29382 390454
rect 28826 389898 29062 390134
rect 29146 389898 29382 390134
rect 28826 354218 29062 354454
rect 29146 354218 29382 354454
rect 28826 353898 29062 354134
rect 29146 353898 29382 354134
rect 28826 318218 29062 318454
rect 29146 318218 29382 318454
rect 28826 317898 29062 318134
rect 29146 317898 29382 318134
rect 28826 282218 29062 282454
rect 29146 282218 29382 282454
rect 28826 281898 29062 282134
rect 29146 281898 29382 282134
rect 28826 246218 29062 246454
rect 29146 246218 29382 246454
rect 28826 245898 29062 246134
rect 29146 245898 29382 246134
rect 28826 210218 29062 210454
rect 29146 210218 29382 210454
rect 28826 209898 29062 210134
rect 29146 209898 29382 210134
rect 28826 174218 29062 174454
rect 29146 174218 29382 174454
rect 28826 173898 29062 174134
rect 29146 173898 29382 174134
rect 28826 138218 29062 138454
rect 29146 138218 29382 138454
rect 28826 137898 29062 138134
rect 29146 137898 29382 138134
rect 28826 102218 29062 102454
rect 29146 102218 29382 102454
rect 28826 101898 29062 102134
rect 29146 101898 29382 102134
rect 28826 66218 29062 66454
rect 29146 66218 29382 66454
rect 28826 65898 29062 66134
rect 29146 65898 29382 66134
rect 28826 30218 29062 30454
rect 29146 30218 29382 30454
rect 28826 29898 29062 30134
rect 29146 29898 29382 30134
rect 28826 -6342 29062 -6106
rect 29146 -6342 29382 -6106
rect 28826 -6662 29062 -6426
rect 29146 -6662 29382 -6426
rect 33326 711322 33562 711558
rect 33646 711322 33882 711558
rect 33326 711002 33562 711238
rect 33646 711002 33882 711238
rect 33326 682718 33562 682954
rect 33646 682718 33882 682954
rect 33326 682398 33562 682634
rect 33646 682398 33882 682634
rect 33326 646718 33562 646954
rect 33646 646718 33882 646954
rect 33326 646398 33562 646634
rect 33646 646398 33882 646634
rect 33326 610718 33562 610954
rect 33646 610718 33882 610954
rect 33326 610398 33562 610634
rect 33646 610398 33882 610634
rect 33326 574718 33562 574954
rect 33646 574718 33882 574954
rect 33326 574398 33562 574634
rect 33646 574398 33882 574634
rect 33326 538718 33562 538954
rect 33646 538718 33882 538954
rect 33326 538398 33562 538634
rect 33646 538398 33882 538634
rect 33326 502718 33562 502954
rect 33646 502718 33882 502954
rect 33326 502398 33562 502634
rect 33646 502398 33882 502634
rect 33326 466718 33562 466954
rect 33646 466718 33882 466954
rect 33326 466398 33562 466634
rect 33646 466398 33882 466634
rect 33326 430718 33562 430954
rect 33646 430718 33882 430954
rect 33326 430398 33562 430634
rect 33646 430398 33882 430634
rect 33326 394718 33562 394954
rect 33646 394718 33882 394954
rect 33326 394398 33562 394634
rect 33646 394398 33882 394634
rect 33326 358718 33562 358954
rect 33646 358718 33882 358954
rect 33326 358398 33562 358634
rect 33646 358398 33882 358634
rect 33326 322718 33562 322954
rect 33646 322718 33882 322954
rect 33326 322398 33562 322634
rect 33646 322398 33882 322634
rect 33326 286718 33562 286954
rect 33646 286718 33882 286954
rect 33326 286398 33562 286634
rect 33646 286398 33882 286634
rect 33326 250718 33562 250954
rect 33646 250718 33882 250954
rect 33326 250398 33562 250634
rect 33646 250398 33882 250634
rect 33326 214718 33562 214954
rect 33646 214718 33882 214954
rect 33326 214398 33562 214634
rect 33646 214398 33882 214634
rect 33326 178718 33562 178954
rect 33646 178718 33882 178954
rect 33326 178398 33562 178634
rect 33646 178398 33882 178634
rect 33326 142718 33562 142954
rect 33646 142718 33882 142954
rect 33326 142398 33562 142634
rect 33646 142398 33882 142634
rect 33326 106718 33562 106954
rect 33646 106718 33882 106954
rect 33326 106398 33562 106634
rect 33646 106398 33882 106634
rect 33326 70718 33562 70954
rect 33646 70718 33882 70954
rect 33326 70398 33562 70634
rect 33646 70398 33882 70634
rect 33326 34718 33562 34954
rect 33646 34718 33882 34954
rect 33326 34398 33562 34634
rect 33646 34398 33882 34634
rect 33326 -7302 33562 -7066
rect 33646 -7302 33882 -7066
rect 33326 -7622 33562 -7386
rect 33646 -7622 33882 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 42326 705562 42562 705798
rect 42646 705562 42882 705798
rect 42326 705242 42562 705478
rect 42646 705242 42882 705478
rect 42326 691718 42562 691954
rect 42646 691718 42882 691954
rect 42326 691398 42562 691634
rect 42646 691398 42882 691634
rect 42326 655718 42562 655954
rect 42646 655718 42882 655954
rect 42326 655398 42562 655634
rect 42646 655398 42882 655634
rect 42326 619718 42562 619954
rect 42646 619718 42882 619954
rect 42326 619398 42562 619634
rect 42646 619398 42882 619634
rect 42326 583718 42562 583954
rect 42646 583718 42882 583954
rect 42326 583398 42562 583634
rect 42646 583398 42882 583634
rect 42326 547718 42562 547954
rect 42646 547718 42882 547954
rect 42326 547398 42562 547634
rect 42646 547398 42882 547634
rect 42326 511718 42562 511954
rect 42646 511718 42882 511954
rect 42326 511398 42562 511634
rect 42646 511398 42882 511634
rect 42326 475718 42562 475954
rect 42646 475718 42882 475954
rect 42326 475398 42562 475634
rect 42646 475398 42882 475634
rect 42326 439718 42562 439954
rect 42646 439718 42882 439954
rect 42326 439398 42562 439634
rect 42646 439398 42882 439634
rect 42326 403718 42562 403954
rect 42646 403718 42882 403954
rect 42326 403398 42562 403634
rect 42646 403398 42882 403634
rect 42326 367718 42562 367954
rect 42646 367718 42882 367954
rect 42326 367398 42562 367634
rect 42646 367398 42882 367634
rect 42326 331718 42562 331954
rect 42646 331718 42882 331954
rect 42326 331398 42562 331634
rect 42646 331398 42882 331634
rect 42326 295718 42562 295954
rect 42646 295718 42882 295954
rect 42326 295398 42562 295634
rect 42646 295398 42882 295634
rect 42326 259718 42562 259954
rect 42646 259718 42882 259954
rect 42326 259398 42562 259634
rect 42646 259398 42882 259634
rect 46826 706522 47062 706758
rect 47146 706522 47382 706758
rect 46826 706202 47062 706438
rect 47146 706202 47382 706438
rect 46826 696218 47062 696454
rect 47146 696218 47382 696454
rect 46826 695898 47062 696134
rect 47146 695898 47382 696134
rect 46826 660218 47062 660454
rect 47146 660218 47382 660454
rect 46826 659898 47062 660134
rect 47146 659898 47382 660134
rect 46826 624218 47062 624454
rect 47146 624218 47382 624454
rect 46826 623898 47062 624134
rect 47146 623898 47382 624134
rect 46826 588218 47062 588454
rect 47146 588218 47382 588454
rect 46826 587898 47062 588134
rect 47146 587898 47382 588134
rect 46826 552218 47062 552454
rect 47146 552218 47382 552454
rect 46826 551898 47062 552134
rect 47146 551898 47382 552134
rect 46826 516218 47062 516454
rect 47146 516218 47382 516454
rect 46826 515898 47062 516134
rect 47146 515898 47382 516134
rect 46826 480218 47062 480454
rect 47146 480218 47382 480454
rect 46826 479898 47062 480134
rect 47146 479898 47382 480134
rect 46826 444218 47062 444454
rect 47146 444218 47382 444454
rect 46826 443898 47062 444134
rect 47146 443898 47382 444134
rect 46826 408218 47062 408454
rect 47146 408218 47382 408454
rect 46826 407898 47062 408134
rect 47146 407898 47382 408134
rect 46826 372218 47062 372454
rect 47146 372218 47382 372454
rect 46826 371898 47062 372134
rect 47146 371898 47382 372134
rect 46826 336218 47062 336454
rect 47146 336218 47382 336454
rect 46826 335898 47062 336134
rect 47146 335898 47382 336134
rect 46826 300218 47062 300454
rect 47146 300218 47382 300454
rect 46826 299898 47062 300134
rect 47146 299898 47382 300134
rect 46826 264218 47062 264454
rect 47146 264218 47382 264454
rect 46826 263898 47062 264134
rect 47146 263898 47382 264134
rect 51326 707482 51562 707718
rect 51646 707482 51882 707718
rect 51326 707162 51562 707398
rect 51646 707162 51882 707398
rect 51326 700718 51562 700954
rect 51646 700718 51882 700954
rect 51326 700398 51562 700634
rect 51646 700398 51882 700634
rect 51326 664718 51562 664954
rect 51646 664718 51882 664954
rect 51326 664398 51562 664634
rect 51646 664398 51882 664634
rect 51326 628718 51562 628954
rect 51646 628718 51882 628954
rect 51326 628398 51562 628634
rect 51646 628398 51882 628634
rect 51326 592718 51562 592954
rect 51646 592718 51882 592954
rect 51326 592398 51562 592634
rect 51646 592398 51882 592634
rect 51326 556718 51562 556954
rect 51646 556718 51882 556954
rect 51326 556398 51562 556634
rect 51646 556398 51882 556634
rect 51326 520718 51562 520954
rect 51646 520718 51882 520954
rect 51326 520398 51562 520634
rect 51646 520398 51882 520634
rect 51326 484718 51562 484954
rect 51646 484718 51882 484954
rect 51326 484398 51562 484634
rect 51646 484398 51882 484634
rect 51326 448718 51562 448954
rect 51646 448718 51882 448954
rect 51326 448398 51562 448634
rect 51646 448398 51882 448634
rect 51326 412718 51562 412954
rect 51646 412718 51882 412954
rect 51326 412398 51562 412634
rect 51646 412398 51882 412634
rect 51326 376718 51562 376954
rect 51646 376718 51882 376954
rect 51326 376398 51562 376634
rect 51646 376398 51882 376634
rect 51326 340718 51562 340954
rect 51646 340718 51882 340954
rect 51326 340398 51562 340634
rect 51646 340398 51882 340634
rect 51326 304718 51562 304954
rect 51646 304718 51882 304954
rect 51326 304398 51562 304634
rect 51646 304398 51882 304634
rect 51326 268718 51562 268954
rect 51646 268718 51882 268954
rect 51326 268398 51562 268634
rect 51646 268398 51882 268634
rect 55826 708442 56062 708678
rect 56146 708442 56382 708678
rect 55826 708122 56062 708358
rect 56146 708122 56382 708358
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 60326 709402 60562 709638
rect 60646 709402 60882 709638
rect 60326 709082 60562 709318
rect 60646 709082 60882 709318
rect 60326 673718 60562 673954
rect 60646 673718 60882 673954
rect 60326 673398 60562 673634
rect 60646 673398 60882 673634
rect 60326 637718 60562 637954
rect 60646 637718 60882 637954
rect 60326 637398 60562 637634
rect 60646 637398 60882 637634
rect 60326 601718 60562 601954
rect 60646 601718 60882 601954
rect 60326 601398 60562 601634
rect 60646 601398 60882 601634
rect 60326 565718 60562 565954
rect 60646 565718 60882 565954
rect 60326 565398 60562 565634
rect 60646 565398 60882 565634
rect 60326 529718 60562 529954
rect 60646 529718 60882 529954
rect 60326 529398 60562 529634
rect 60646 529398 60882 529634
rect 60326 493718 60562 493954
rect 60646 493718 60882 493954
rect 60326 493398 60562 493634
rect 60646 493398 60882 493634
rect 60326 457718 60562 457954
rect 60646 457718 60882 457954
rect 60326 457398 60562 457634
rect 60646 457398 60882 457634
rect 60326 421718 60562 421954
rect 60646 421718 60882 421954
rect 60326 421398 60562 421634
rect 60646 421398 60882 421634
rect 60326 385718 60562 385954
rect 60646 385718 60882 385954
rect 60326 385398 60562 385634
rect 60646 385398 60882 385634
rect 60326 349718 60562 349954
rect 60646 349718 60882 349954
rect 60326 349398 60562 349634
rect 60646 349398 60882 349634
rect 60326 313718 60562 313954
rect 60646 313718 60882 313954
rect 60326 313398 60562 313634
rect 60646 313398 60882 313634
rect 60326 277718 60562 277954
rect 60646 277718 60882 277954
rect 60326 277398 60562 277634
rect 60646 277398 60882 277634
rect 64826 710362 65062 710598
rect 65146 710362 65382 710598
rect 64826 710042 65062 710278
rect 65146 710042 65382 710278
rect 64826 678218 65062 678454
rect 65146 678218 65382 678454
rect 64826 677898 65062 678134
rect 65146 677898 65382 678134
rect 64826 642218 65062 642454
rect 65146 642218 65382 642454
rect 64826 641898 65062 642134
rect 65146 641898 65382 642134
rect 64826 606218 65062 606454
rect 65146 606218 65382 606454
rect 64826 605898 65062 606134
rect 65146 605898 65382 606134
rect 64826 570218 65062 570454
rect 65146 570218 65382 570454
rect 64826 569898 65062 570134
rect 65146 569898 65382 570134
rect 64826 534218 65062 534454
rect 65146 534218 65382 534454
rect 64826 533898 65062 534134
rect 65146 533898 65382 534134
rect 64826 498218 65062 498454
rect 65146 498218 65382 498454
rect 64826 497898 65062 498134
rect 65146 497898 65382 498134
rect 64826 462218 65062 462454
rect 65146 462218 65382 462454
rect 64826 461898 65062 462134
rect 65146 461898 65382 462134
rect 64826 426218 65062 426454
rect 65146 426218 65382 426454
rect 64826 425898 65062 426134
rect 65146 425898 65382 426134
rect 64826 390218 65062 390454
rect 65146 390218 65382 390454
rect 64826 389898 65062 390134
rect 65146 389898 65382 390134
rect 64826 354218 65062 354454
rect 65146 354218 65382 354454
rect 64826 353898 65062 354134
rect 65146 353898 65382 354134
rect 64826 318218 65062 318454
rect 65146 318218 65382 318454
rect 64826 317898 65062 318134
rect 65146 317898 65382 318134
rect 64826 282218 65062 282454
rect 65146 282218 65382 282454
rect 64826 281898 65062 282134
rect 65146 281898 65382 282134
rect 69326 711322 69562 711558
rect 69646 711322 69882 711558
rect 69326 711002 69562 711238
rect 69646 711002 69882 711238
rect 69326 682718 69562 682954
rect 69646 682718 69882 682954
rect 69326 682398 69562 682634
rect 69646 682398 69882 682634
rect 69326 646718 69562 646954
rect 69646 646718 69882 646954
rect 69326 646398 69562 646634
rect 69646 646398 69882 646634
rect 69326 610718 69562 610954
rect 69646 610718 69882 610954
rect 69326 610398 69562 610634
rect 69646 610398 69882 610634
rect 69326 574718 69562 574954
rect 69646 574718 69882 574954
rect 69326 574398 69562 574634
rect 69646 574398 69882 574634
rect 69326 538718 69562 538954
rect 69646 538718 69882 538954
rect 69326 538398 69562 538634
rect 69646 538398 69882 538634
rect 69326 502718 69562 502954
rect 69646 502718 69882 502954
rect 69326 502398 69562 502634
rect 69646 502398 69882 502634
rect 69326 466718 69562 466954
rect 69646 466718 69882 466954
rect 69326 466398 69562 466634
rect 69646 466398 69882 466634
rect 69326 430718 69562 430954
rect 69646 430718 69882 430954
rect 69326 430398 69562 430634
rect 69646 430398 69882 430634
rect 69326 394718 69562 394954
rect 69646 394718 69882 394954
rect 69326 394398 69562 394634
rect 69646 394398 69882 394634
rect 69326 358718 69562 358954
rect 69646 358718 69882 358954
rect 69326 358398 69562 358634
rect 69646 358398 69882 358634
rect 69326 322718 69562 322954
rect 69646 322718 69882 322954
rect 69326 322398 69562 322634
rect 69646 322398 69882 322634
rect 69326 286718 69562 286954
rect 69646 286718 69882 286954
rect 69326 286398 69562 286634
rect 69646 286398 69882 286634
rect 69326 250718 69562 250954
rect 69646 250718 69882 250954
rect 69326 250398 69562 250634
rect 69646 250398 69882 250634
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 78326 705562 78562 705798
rect 78646 705562 78882 705798
rect 78326 705242 78562 705478
rect 78646 705242 78882 705478
rect 78326 691718 78562 691954
rect 78646 691718 78882 691954
rect 78326 691398 78562 691634
rect 78646 691398 78882 691634
rect 78326 655718 78562 655954
rect 78646 655718 78882 655954
rect 78326 655398 78562 655634
rect 78646 655398 78882 655634
rect 78326 619718 78562 619954
rect 78646 619718 78882 619954
rect 78326 619398 78562 619634
rect 78646 619398 78882 619634
rect 78326 583718 78562 583954
rect 78646 583718 78882 583954
rect 78326 583398 78562 583634
rect 78646 583398 78882 583634
rect 78326 547718 78562 547954
rect 78646 547718 78882 547954
rect 78326 547398 78562 547634
rect 78646 547398 78882 547634
rect 78326 511718 78562 511954
rect 78646 511718 78882 511954
rect 78326 511398 78562 511634
rect 78646 511398 78882 511634
rect 78326 475718 78562 475954
rect 78646 475718 78882 475954
rect 78326 475398 78562 475634
rect 78646 475398 78882 475634
rect 78326 439718 78562 439954
rect 78646 439718 78882 439954
rect 78326 439398 78562 439634
rect 78646 439398 78882 439634
rect 78326 403718 78562 403954
rect 78646 403718 78882 403954
rect 78326 403398 78562 403634
rect 78646 403398 78882 403634
rect 78326 367718 78562 367954
rect 78646 367718 78882 367954
rect 78326 367398 78562 367634
rect 78646 367398 78882 367634
rect 78326 331718 78562 331954
rect 78646 331718 78882 331954
rect 78326 331398 78562 331634
rect 78646 331398 78882 331634
rect 78326 295718 78562 295954
rect 78646 295718 78882 295954
rect 78326 295398 78562 295634
rect 78646 295398 78882 295634
rect 78326 259718 78562 259954
rect 78646 259718 78882 259954
rect 78326 259398 78562 259634
rect 78646 259398 78882 259634
rect 82826 706522 83062 706758
rect 83146 706522 83382 706758
rect 82826 706202 83062 706438
rect 83146 706202 83382 706438
rect 82826 696218 83062 696454
rect 83146 696218 83382 696454
rect 82826 695898 83062 696134
rect 83146 695898 83382 696134
rect 82826 660218 83062 660454
rect 83146 660218 83382 660454
rect 82826 659898 83062 660134
rect 83146 659898 83382 660134
rect 82826 624218 83062 624454
rect 83146 624218 83382 624454
rect 82826 623898 83062 624134
rect 83146 623898 83382 624134
rect 82826 588218 83062 588454
rect 83146 588218 83382 588454
rect 82826 587898 83062 588134
rect 83146 587898 83382 588134
rect 82826 552218 83062 552454
rect 83146 552218 83382 552454
rect 82826 551898 83062 552134
rect 83146 551898 83382 552134
rect 82826 516218 83062 516454
rect 83146 516218 83382 516454
rect 82826 515898 83062 516134
rect 83146 515898 83382 516134
rect 82826 480218 83062 480454
rect 83146 480218 83382 480454
rect 82826 479898 83062 480134
rect 83146 479898 83382 480134
rect 82826 444218 83062 444454
rect 83146 444218 83382 444454
rect 82826 443898 83062 444134
rect 83146 443898 83382 444134
rect 82826 408218 83062 408454
rect 83146 408218 83382 408454
rect 82826 407898 83062 408134
rect 83146 407898 83382 408134
rect 82826 372218 83062 372454
rect 83146 372218 83382 372454
rect 82826 371898 83062 372134
rect 83146 371898 83382 372134
rect 82826 336218 83062 336454
rect 83146 336218 83382 336454
rect 82826 335898 83062 336134
rect 83146 335898 83382 336134
rect 82826 300218 83062 300454
rect 83146 300218 83382 300454
rect 82826 299898 83062 300134
rect 83146 299898 83382 300134
rect 82826 264218 83062 264454
rect 83146 264218 83382 264454
rect 82826 263898 83062 264134
rect 83146 263898 83382 264134
rect 87326 707482 87562 707718
rect 87646 707482 87882 707718
rect 87326 707162 87562 707398
rect 87646 707162 87882 707398
rect 87326 700718 87562 700954
rect 87646 700718 87882 700954
rect 87326 700398 87562 700634
rect 87646 700398 87882 700634
rect 87326 664718 87562 664954
rect 87646 664718 87882 664954
rect 87326 664398 87562 664634
rect 87646 664398 87882 664634
rect 87326 628718 87562 628954
rect 87646 628718 87882 628954
rect 87326 628398 87562 628634
rect 87646 628398 87882 628634
rect 87326 592718 87562 592954
rect 87646 592718 87882 592954
rect 87326 592398 87562 592634
rect 87646 592398 87882 592634
rect 87326 556718 87562 556954
rect 87646 556718 87882 556954
rect 87326 556398 87562 556634
rect 87646 556398 87882 556634
rect 87326 520718 87562 520954
rect 87646 520718 87882 520954
rect 87326 520398 87562 520634
rect 87646 520398 87882 520634
rect 87326 484718 87562 484954
rect 87646 484718 87882 484954
rect 87326 484398 87562 484634
rect 87646 484398 87882 484634
rect 87326 448718 87562 448954
rect 87646 448718 87882 448954
rect 87326 448398 87562 448634
rect 87646 448398 87882 448634
rect 87326 412718 87562 412954
rect 87646 412718 87882 412954
rect 87326 412398 87562 412634
rect 87646 412398 87882 412634
rect 87326 376718 87562 376954
rect 87646 376718 87882 376954
rect 87326 376398 87562 376634
rect 87646 376398 87882 376634
rect 87326 340718 87562 340954
rect 87646 340718 87882 340954
rect 87326 340398 87562 340634
rect 87646 340398 87882 340634
rect 87326 304718 87562 304954
rect 87646 304718 87882 304954
rect 87326 304398 87562 304634
rect 87646 304398 87882 304634
rect 87326 268718 87562 268954
rect 87646 268718 87882 268954
rect 87326 268398 87562 268634
rect 87646 268398 87882 268634
rect 91826 708442 92062 708678
rect 92146 708442 92382 708678
rect 91826 708122 92062 708358
rect 92146 708122 92382 708358
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 96326 709402 96562 709638
rect 96646 709402 96882 709638
rect 96326 709082 96562 709318
rect 96646 709082 96882 709318
rect 96326 673718 96562 673954
rect 96646 673718 96882 673954
rect 96326 673398 96562 673634
rect 96646 673398 96882 673634
rect 96326 637718 96562 637954
rect 96646 637718 96882 637954
rect 96326 637398 96562 637634
rect 96646 637398 96882 637634
rect 96326 601718 96562 601954
rect 96646 601718 96882 601954
rect 96326 601398 96562 601634
rect 96646 601398 96882 601634
rect 96326 565718 96562 565954
rect 96646 565718 96882 565954
rect 96326 565398 96562 565634
rect 96646 565398 96882 565634
rect 96326 529718 96562 529954
rect 96646 529718 96882 529954
rect 96326 529398 96562 529634
rect 96646 529398 96882 529634
rect 96326 493718 96562 493954
rect 96646 493718 96882 493954
rect 96326 493398 96562 493634
rect 96646 493398 96882 493634
rect 96326 457718 96562 457954
rect 96646 457718 96882 457954
rect 96326 457398 96562 457634
rect 96646 457398 96882 457634
rect 96326 421718 96562 421954
rect 96646 421718 96882 421954
rect 96326 421398 96562 421634
rect 96646 421398 96882 421634
rect 96326 385718 96562 385954
rect 96646 385718 96882 385954
rect 96326 385398 96562 385634
rect 96646 385398 96882 385634
rect 96326 349718 96562 349954
rect 96646 349718 96882 349954
rect 96326 349398 96562 349634
rect 96646 349398 96882 349634
rect 96326 313718 96562 313954
rect 96646 313718 96882 313954
rect 96326 313398 96562 313634
rect 96646 313398 96882 313634
rect 96326 277718 96562 277954
rect 96646 277718 96882 277954
rect 96326 277398 96562 277634
rect 96646 277398 96882 277634
rect 100826 710362 101062 710598
rect 101146 710362 101382 710598
rect 100826 710042 101062 710278
rect 101146 710042 101382 710278
rect 100826 678218 101062 678454
rect 101146 678218 101382 678454
rect 100826 677898 101062 678134
rect 101146 677898 101382 678134
rect 100826 642218 101062 642454
rect 101146 642218 101382 642454
rect 100826 641898 101062 642134
rect 101146 641898 101382 642134
rect 100826 606218 101062 606454
rect 101146 606218 101382 606454
rect 100826 605898 101062 606134
rect 101146 605898 101382 606134
rect 100826 570218 101062 570454
rect 101146 570218 101382 570454
rect 100826 569898 101062 570134
rect 101146 569898 101382 570134
rect 100826 534218 101062 534454
rect 101146 534218 101382 534454
rect 100826 533898 101062 534134
rect 101146 533898 101382 534134
rect 100826 498218 101062 498454
rect 101146 498218 101382 498454
rect 100826 497898 101062 498134
rect 101146 497898 101382 498134
rect 100826 462218 101062 462454
rect 101146 462218 101382 462454
rect 100826 461898 101062 462134
rect 101146 461898 101382 462134
rect 100826 426218 101062 426454
rect 101146 426218 101382 426454
rect 100826 425898 101062 426134
rect 101146 425898 101382 426134
rect 100826 390218 101062 390454
rect 101146 390218 101382 390454
rect 100826 389898 101062 390134
rect 101146 389898 101382 390134
rect 100826 354218 101062 354454
rect 101146 354218 101382 354454
rect 100826 353898 101062 354134
rect 101146 353898 101382 354134
rect 100826 318218 101062 318454
rect 101146 318218 101382 318454
rect 100826 317898 101062 318134
rect 101146 317898 101382 318134
rect 100826 282218 101062 282454
rect 101146 282218 101382 282454
rect 100826 281898 101062 282134
rect 101146 281898 101382 282134
rect 105326 711322 105562 711558
rect 105646 711322 105882 711558
rect 105326 711002 105562 711238
rect 105646 711002 105882 711238
rect 105326 682718 105562 682954
rect 105646 682718 105882 682954
rect 105326 682398 105562 682634
rect 105646 682398 105882 682634
rect 105326 646718 105562 646954
rect 105646 646718 105882 646954
rect 105326 646398 105562 646634
rect 105646 646398 105882 646634
rect 105326 610718 105562 610954
rect 105646 610718 105882 610954
rect 105326 610398 105562 610634
rect 105646 610398 105882 610634
rect 105326 574718 105562 574954
rect 105646 574718 105882 574954
rect 105326 574398 105562 574634
rect 105646 574398 105882 574634
rect 105326 538718 105562 538954
rect 105646 538718 105882 538954
rect 105326 538398 105562 538634
rect 105646 538398 105882 538634
rect 105326 502718 105562 502954
rect 105646 502718 105882 502954
rect 105326 502398 105562 502634
rect 105646 502398 105882 502634
rect 105326 466718 105562 466954
rect 105646 466718 105882 466954
rect 105326 466398 105562 466634
rect 105646 466398 105882 466634
rect 105326 430718 105562 430954
rect 105646 430718 105882 430954
rect 105326 430398 105562 430634
rect 105646 430398 105882 430634
rect 105326 394718 105562 394954
rect 105646 394718 105882 394954
rect 105326 394398 105562 394634
rect 105646 394398 105882 394634
rect 105326 358718 105562 358954
rect 105646 358718 105882 358954
rect 105326 358398 105562 358634
rect 105646 358398 105882 358634
rect 105326 322718 105562 322954
rect 105646 322718 105882 322954
rect 105326 322398 105562 322634
rect 105646 322398 105882 322634
rect 105326 286718 105562 286954
rect 105646 286718 105882 286954
rect 105326 286398 105562 286634
rect 105646 286398 105882 286634
rect 105326 250718 105562 250954
rect 105646 250718 105882 250954
rect 105326 250398 105562 250634
rect 105646 250398 105882 250634
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 114326 705562 114562 705798
rect 114646 705562 114882 705798
rect 114326 705242 114562 705478
rect 114646 705242 114882 705478
rect 114326 691718 114562 691954
rect 114646 691718 114882 691954
rect 114326 691398 114562 691634
rect 114646 691398 114882 691634
rect 114326 655718 114562 655954
rect 114646 655718 114882 655954
rect 114326 655398 114562 655634
rect 114646 655398 114882 655634
rect 114326 619718 114562 619954
rect 114646 619718 114882 619954
rect 114326 619398 114562 619634
rect 114646 619398 114882 619634
rect 114326 583718 114562 583954
rect 114646 583718 114882 583954
rect 114326 583398 114562 583634
rect 114646 583398 114882 583634
rect 114326 547718 114562 547954
rect 114646 547718 114882 547954
rect 114326 547398 114562 547634
rect 114646 547398 114882 547634
rect 114326 511718 114562 511954
rect 114646 511718 114882 511954
rect 114326 511398 114562 511634
rect 114646 511398 114882 511634
rect 114326 475718 114562 475954
rect 114646 475718 114882 475954
rect 114326 475398 114562 475634
rect 114646 475398 114882 475634
rect 114326 439718 114562 439954
rect 114646 439718 114882 439954
rect 114326 439398 114562 439634
rect 114646 439398 114882 439634
rect 114326 403718 114562 403954
rect 114646 403718 114882 403954
rect 114326 403398 114562 403634
rect 114646 403398 114882 403634
rect 114326 367718 114562 367954
rect 114646 367718 114882 367954
rect 114326 367398 114562 367634
rect 114646 367398 114882 367634
rect 114326 331718 114562 331954
rect 114646 331718 114882 331954
rect 114326 331398 114562 331634
rect 114646 331398 114882 331634
rect 114326 295718 114562 295954
rect 114646 295718 114882 295954
rect 114326 295398 114562 295634
rect 114646 295398 114882 295634
rect 114326 259718 114562 259954
rect 114646 259718 114882 259954
rect 114326 259398 114562 259634
rect 114646 259398 114882 259634
rect 118826 706522 119062 706758
rect 119146 706522 119382 706758
rect 118826 706202 119062 706438
rect 119146 706202 119382 706438
rect 118826 696218 119062 696454
rect 119146 696218 119382 696454
rect 118826 695898 119062 696134
rect 119146 695898 119382 696134
rect 118826 660218 119062 660454
rect 119146 660218 119382 660454
rect 118826 659898 119062 660134
rect 119146 659898 119382 660134
rect 118826 624218 119062 624454
rect 119146 624218 119382 624454
rect 118826 623898 119062 624134
rect 119146 623898 119382 624134
rect 118826 588218 119062 588454
rect 119146 588218 119382 588454
rect 118826 587898 119062 588134
rect 119146 587898 119382 588134
rect 118826 552218 119062 552454
rect 119146 552218 119382 552454
rect 118826 551898 119062 552134
rect 119146 551898 119382 552134
rect 118826 516218 119062 516454
rect 119146 516218 119382 516454
rect 118826 515898 119062 516134
rect 119146 515898 119382 516134
rect 118826 480218 119062 480454
rect 119146 480218 119382 480454
rect 118826 479898 119062 480134
rect 119146 479898 119382 480134
rect 118826 444218 119062 444454
rect 119146 444218 119382 444454
rect 118826 443898 119062 444134
rect 119146 443898 119382 444134
rect 118826 408218 119062 408454
rect 119146 408218 119382 408454
rect 118826 407898 119062 408134
rect 119146 407898 119382 408134
rect 118826 372218 119062 372454
rect 119146 372218 119382 372454
rect 118826 371898 119062 372134
rect 119146 371898 119382 372134
rect 118826 336218 119062 336454
rect 119146 336218 119382 336454
rect 118826 335898 119062 336134
rect 119146 335898 119382 336134
rect 118826 300218 119062 300454
rect 119146 300218 119382 300454
rect 118826 299898 119062 300134
rect 119146 299898 119382 300134
rect 118826 264218 119062 264454
rect 119146 264218 119382 264454
rect 118826 263898 119062 264134
rect 119146 263898 119382 264134
rect 123326 707482 123562 707718
rect 123646 707482 123882 707718
rect 123326 707162 123562 707398
rect 123646 707162 123882 707398
rect 123326 700718 123562 700954
rect 123646 700718 123882 700954
rect 123326 700398 123562 700634
rect 123646 700398 123882 700634
rect 123326 664718 123562 664954
rect 123646 664718 123882 664954
rect 123326 664398 123562 664634
rect 123646 664398 123882 664634
rect 123326 628718 123562 628954
rect 123646 628718 123882 628954
rect 123326 628398 123562 628634
rect 123646 628398 123882 628634
rect 123326 592718 123562 592954
rect 123646 592718 123882 592954
rect 123326 592398 123562 592634
rect 123646 592398 123882 592634
rect 123326 556718 123562 556954
rect 123646 556718 123882 556954
rect 123326 556398 123562 556634
rect 123646 556398 123882 556634
rect 123326 520718 123562 520954
rect 123646 520718 123882 520954
rect 123326 520398 123562 520634
rect 123646 520398 123882 520634
rect 123326 484718 123562 484954
rect 123646 484718 123882 484954
rect 123326 484398 123562 484634
rect 123646 484398 123882 484634
rect 123326 448718 123562 448954
rect 123646 448718 123882 448954
rect 123326 448398 123562 448634
rect 123646 448398 123882 448634
rect 123326 412718 123562 412954
rect 123646 412718 123882 412954
rect 123326 412398 123562 412634
rect 123646 412398 123882 412634
rect 123326 376718 123562 376954
rect 123646 376718 123882 376954
rect 123326 376398 123562 376634
rect 123646 376398 123882 376634
rect 123326 340718 123562 340954
rect 123646 340718 123882 340954
rect 123326 340398 123562 340634
rect 123646 340398 123882 340634
rect 123326 304718 123562 304954
rect 123646 304718 123882 304954
rect 123326 304398 123562 304634
rect 123646 304398 123882 304634
rect 123326 268718 123562 268954
rect 123646 268718 123882 268954
rect 123326 268398 123562 268634
rect 123646 268398 123882 268634
rect 127826 708442 128062 708678
rect 128146 708442 128382 708678
rect 127826 708122 128062 708358
rect 128146 708122 128382 708358
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 132326 709402 132562 709638
rect 132646 709402 132882 709638
rect 132326 709082 132562 709318
rect 132646 709082 132882 709318
rect 132326 673718 132562 673954
rect 132646 673718 132882 673954
rect 132326 673398 132562 673634
rect 132646 673398 132882 673634
rect 132326 637718 132562 637954
rect 132646 637718 132882 637954
rect 132326 637398 132562 637634
rect 132646 637398 132882 637634
rect 132326 601718 132562 601954
rect 132646 601718 132882 601954
rect 132326 601398 132562 601634
rect 132646 601398 132882 601634
rect 132326 565718 132562 565954
rect 132646 565718 132882 565954
rect 132326 565398 132562 565634
rect 132646 565398 132882 565634
rect 132326 529718 132562 529954
rect 132646 529718 132882 529954
rect 132326 529398 132562 529634
rect 132646 529398 132882 529634
rect 132326 493718 132562 493954
rect 132646 493718 132882 493954
rect 132326 493398 132562 493634
rect 132646 493398 132882 493634
rect 132326 457718 132562 457954
rect 132646 457718 132882 457954
rect 132326 457398 132562 457634
rect 132646 457398 132882 457634
rect 132326 421718 132562 421954
rect 132646 421718 132882 421954
rect 132326 421398 132562 421634
rect 132646 421398 132882 421634
rect 132326 385718 132562 385954
rect 132646 385718 132882 385954
rect 132326 385398 132562 385634
rect 132646 385398 132882 385634
rect 132326 349718 132562 349954
rect 132646 349718 132882 349954
rect 132326 349398 132562 349634
rect 132646 349398 132882 349634
rect 132326 313718 132562 313954
rect 132646 313718 132882 313954
rect 132326 313398 132562 313634
rect 132646 313398 132882 313634
rect 132326 277718 132562 277954
rect 132646 277718 132882 277954
rect 132326 277398 132562 277634
rect 132646 277398 132882 277634
rect 136826 710362 137062 710598
rect 137146 710362 137382 710598
rect 136826 710042 137062 710278
rect 137146 710042 137382 710278
rect 136826 678218 137062 678454
rect 137146 678218 137382 678454
rect 136826 677898 137062 678134
rect 137146 677898 137382 678134
rect 136826 642218 137062 642454
rect 137146 642218 137382 642454
rect 136826 641898 137062 642134
rect 137146 641898 137382 642134
rect 136826 606218 137062 606454
rect 137146 606218 137382 606454
rect 136826 605898 137062 606134
rect 137146 605898 137382 606134
rect 136826 570218 137062 570454
rect 137146 570218 137382 570454
rect 136826 569898 137062 570134
rect 137146 569898 137382 570134
rect 136826 534218 137062 534454
rect 137146 534218 137382 534454
rect 136826 533898 137062 534134
rect 137146 533898 137382 534134
rect 136826 498218 137062 498454
rect 137146 498218 137382 498454
rect 136826 497898 137062 498134
rect 137146 497898 137382 498134
rect 136826 462218 137062 462454
rect 137146 462218 137382 462454
rect 136826 461898 137062 462134
rect 137146 461898 137382 462134
rect 136826 426218 137062 426454
rect 137146 426218 137382 426454
rect 136826 425898 137062 426134
rect 137146 425898 137382 426134
rect 136826 390218 137062 390454
rect 137146 390218 137382 390454
rect 136826 389898 137062 390134
rect 137146 389898 137382 390134
rect 136826 354218 137062 354454
rect 137146 354218 137382 354454
rect 136826 353898 137062 354134
rect 137146 353898 137382 354134
rect 136826 318218 137062 318454
rect 137146 318218 137382 318454
rect 136826 317898 137062 318134
rect 137146 317898 137382 318134
rect 136826 282218 137062 282454
rect 137146 282218 137382 282454
rect 136826 281898 137062 282134
rect 137146 281898 137382 282134
rect 141326 711322 141562 711558
rect 141646 711322 141882 711558
rect 141326 711002 141562 711238
rect 141646 711002 141882 711238
rect 141326 682718 141562 682954
rect 141646 682718 141882 682954
rect 141326 682398 141562 682634
rect 141646 682398 141882 682634
rect 141326 646718 141562 646954
rect 141646 646718 141882 646954
rect 141326 646398 141562 646634
rect 141646 646398 141882 646634
rect 141326 610718 141562 610954
rect 141646 610718 141882 610954
rect 141326 610398 141562 610634
rect 141646 610398 141882 610634
rect 141326 574718 141562 574954
rect 141646 574718 141882 574954
rect 141326 574398 141562 574634
rect 141646 574398 141882 574634
rect 141326 538718 141562 538954
rect 141646 538718 141882 538954
rect 141326 538398 141562 538634
rect 141646 538398 141882 538634
rect 141326 502718 141562 502954
rect 141646 502718 141882 502954
rect 141326 502398 141562 502634
rect 141646 502398 141882 502634
rect 141326 466718 141562 466954
rect 141646 466718 141882 466954
rect 141326 466398 141562 466634
rect 141646 466398 141882 466634
rect 141326 430718 141562 430954
rect 141646 430718 141882 430954
rect 141326 430398 141562 430634
rect 141646 430398 141882 430634
rect 141326 394718 141562 394954
rect 141646 394718 141882 394954
rect 141326 394398 141562 394634
rect 141646 394398 141882 394634
rect 141326 358718 141562 358954
rect 141646 358718 141882 358954
rect 141326 358398 141562 358634
rect 141646 358398 141882 358634
rect 141326 322718 141562 322954
rect 141646 322718 141882 322954
rect 141326 322398 141562 322634
rect 141646 322398 141882 322634
rect 141326 286718 141562 286954
rect 141646 286718 141882 286954
rect 141326 286398 141562 286634
rect 141646 286398 141882 286634
rect 141326 250718 141562 250954
rect 141646 250718 141882 250954
rect 141326 250398 141562 250634
rect 141646 250398 141882 250634
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 150326 705562 150562 705798
rect 150646 705562 150882 705798
rect 150326 705242 150562 705478
rect 150646 705242 150882 705478
rect 150326 691718 150562 691954
rect 150646 691718 150882 691954
rect 150326 691398 150562 691634
rect 150646 691398 150882 691634
rect 150326 655718 150562 655954
rect 150646 655718 150882 655954
rect 150326 655398 150562 655634
rect 150646 655398 150882 655634
rect 150326 619718 150562 619954
rect 150646 619718 150882 619954
rect 150326 619398 150562 619634
rect 150646 619398 150882 619634
rect 150326 583718 150562 583954
rect 150646 583718 150882 583954
rect 150326 583398 150562 583634
rect 150646 583398 150882 583634
rect 150326 547718 150562 547954
rect 150646 547718 150882 547954
rect 150326 547398 150562 547634
rect 150646 547398 150882 547634
rect 150326 511718 150562 511954
rect 150646 511718 150882 511954
rect 150326 511398 150562 511634
rect 150646 511398 150882 511634
rect 150326 475718 150562 475954
rect 150646 475718 150882 475954
rect 150326 475398 150562 475634
rect 150646 475398 150882 475634
rect 150326 439718 150562 439954
rect 150646 439718 150882 439954
rect 150326 439398 150562 439634
rect 150646 439398 150882 439634
rect 150326 403718 150562 403954
rect 150646 403718 150882 403954
rect 150326 403398 150562 403634
rect 150646 403398 150882 403634
rect 150326 367718 150562 367954
rect 150646 367718 150882 367954
rect 150326 367398 150562 367634
rect 150646 367398 150882 367634
rect 150326 331718 150562 331954
rect 150646 331718 150882 331954
rect 150326 331398 150562 331634
rect 150646 331398 150882 331634
rect 150326 295718 150562 295954
rect 150646 295718 150882 295954
rect 150326 295398 150562 295634
rect 150646 295398 150882 295634
rect 150326 259718 150562 259954
rect 150646 259718 150882 259954
rect 150326 259398 150562 259634
rect 150646 259398 150882 259634
rect 154826 706522 155062 706758
rect 155146 706522 155382 706758
rect 154826 706202 155062 706438
rect 155146 706202 155382 706438
rect 154826 696218 155062 696454
rect 155146 696218 155382 696454
rect 154826 695898 155062 696134
rect 155146 695898 155382 696134
rect 154826 660218 155062 660454
rect 155146 660218 155382 660454
rect 154826 659898 155062 660134
rect 155146 659898 155382 660134
rect 154826 624218 155062 624454
rect 155146 624218 155382 624454
rect 154826 623898 155062 624134
rect 155146 623898 155382 624134
rect 154826 588218 155062 588454
rect 155146 588218 155382 588454
rect 154826 587898 155062 588134
rect 155146 587898 155382 588134
rect 154826 552218 155062 552454
rect 155146 552218 155382 552454
rect 154826 551898 155062 552134
rect 155146 551898 155382 552134
rect 154826 516218 155062 516454
rect 155146 516218 155382 516454
rect 154826 515898 155062 516134
rect 155146 515898 155382 516134
rect 154826 480218 155062 480454
rect 155146 480218 155382 480454
rect 154826 479898 155062 480134
rect 155146 479898 155382 480134
rect 154826 444218 155062 444454
rect 155146 444218 155382 444454
rect 154826 443898 155062 444134
rect 155146 443898 155382 444134
rect 154826 408218 155062 408454
rect 155146 408218 155382 408454
rect 154826 407898 155062 408134
rect 155146 407898 155382 408134
rect 154826 372218 155062 372454
rect 155146 372218 155382 372454
rect 154826 371898 155062 372134
rect 155146 371898 155382 372134
rect 154826 336218 155062 336454
rect 155146 336218 155382 336454
rect 154826 335898 155062 336134
rect 155146 335898 155382 336134
rect 154826 300218 155062 300454
rect 155146 300218 155382 300454
rect 154826 299898 155062 300134
rect 155146 299898 155382 300134
rect 154826 264218 155062 264454
rect 155146 264218 155382 264454
rect 154826 263898 155062 264134
rect 155146 263898 155382 264134
rect 159326 707482 159562 707718
rect 159646 707482 159882 707718
rect 159326 707162 159562 707398
rect 159646 707162 159882 707398
rect 159326 700718 159562 700954
rect 159646 700718 159882 700954
rect 159326 700398 159562 700634
rect 159646 700398 159882 700634
rect 159326 664718 159562 664954
rect 159646 664718 159882 664954
rect 159326 664398 159562 664634
rect 159646 664398 159882 664634
rect 159326 628718 159562 628954
rect 159646 628718 159882 628954
rect 159326 628398 159562 628634
rect 159646 628398 159882 628634
rect 159326 592718 159562 592954
rect 159646 592718 159882 592954
rect 159326 592398 159562 592634
rect 159646 592398 159882 592634
rect 159326 556718 159562 556954
rect 159646 556718 159882 556954
rect 159326 556398 159562 556634
rect 159646 556398 159882 556634
rect 159326 520718 159562 520954
rect 159646 520718 159882 520954
rect 159326 520398 159562 520634
rect 159646 520398 159882 520634
rect 159326 484718 159562 484954
rect 159646 484718 159882 484954
rect 159326 484398 159562 484634
rect 159646 484398 159882 484634
rect 159326 448718 159562 448954
rect 159646 448718 159882 448954
rect 159326 448398 159562 448634
rect 159646 448398 159882 448634
rect 159326 412718 159562 412954
rect 159646 412718 159882 412954
rect 159326 412398 159562 412634
rect 159646 412398 159882 412634
rect 159326 376718 159562 376954
rect 159646 376718 159882 376954
rect 159326 376398 159562 376634
rect 159646 376398 159882 376634
rect 159326 340718 159562 340954
rect 159646 340718 159882 340954
rect 159326 340398 159562 340634
rect 159646 340398 159882 340634
rect 159326 304718 159562 304954
rect 159646 304718 159882 304954
rect 159326 304398 159562 304634
rect 159646 304398 159882 304634
rect 159326 268718 159562 268954
rect 159646 268718 159882 268954
rect 159326 268398 159562 268634
rect 159646 268398 159882 268634
rect 163826 708442 164062 708678
rect 164146 708442 164382 708678
rect 163826 708122 164062 708358
rect 164146 708122 164382 708358
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 168326 709402 168562 709638
rect 168646 709402 168882 709638
rect 168326 709082 168562 709318
rect 168646 709082 168882 709318
rect 168326 673718 168562 673954
rect 168646 673718 168882 673954
rect 168326 673398 168562 673634
rect 168646 673398 168882 673634
rect 168326 637718 168562 637954
rect 168646 637718 168882 637954
rect 168326 637398 168562 637634
rect 168646 637398 168882 637634
rect 168326 601718 168562 601954
rect 168646 601718 168882 601954
rect 168326 601398 168562 601634
rect 168646 601398 168882 601634
rect 168326 565718 168562 565954
rect 168646 565718 168882 565954
rect 168326 565398 168562 565634
rect 168646 565398 168882 565634
rect 168326 529718 168562 529954
rect 168646 529718 168882 529954
rect 168326 529398 168562 529634
rect 168646 529398 168882 529634
rect 168326 493718 168562 493954
rect 168646 493718 168882 493954
rect 168326 493398 168562 493634
rect 168646 493398 168882 493634
rect 168326 457718 168562 457954
rect 168646 457718 168882 457954
rect 168326 457398 168562 457634
rect 168646 457398 168882 457634
rect 168326 421718 168562 421954
rect 168646 421718 168882 421954
rect 168326 421398 168562 421634
rect 168646 421398 168882 421634
rect 168326 385718 168562 385954
rect 168646 385718 168882 385954
rect 168326 385398 168562 385634
rect 168646 385398 168882 385634
rect 168326 349718 168562 349954
rect 168646 349718 168882 349954
rect 168326 349398 168562 349634
rect 168646 349398 168882 349634
rect 168326 313718 168562 313954
rect 168646 313718 168882 313954
rect 168326 313398 168562 313634
rect 168646 313398 168882 313634
rect 168326 277718 168562 277954
rect 168646 277718 168882 277954
rect 168326 277398 168562 277634
rect 168646 277398 168882 277634
rect 172826 710362 173062 710598
rect 173146 710362 173382 710598
rect 172826 710042 173062 710278
rect 173146 710042 173382 710278
rect 172826 678218 173062 678454
rect 173146 678218 173382 678454
rect 172826 677898 173062 678134
rect 173146 677898 173382 678134
rect 172826 642218 173062 642454
rect 173146 642218 173382 642454
rect 172826 641898 173062 642134
rect 173146 641898 173382 642134
rect 172826 606218 173062 606454
rect 173146 606218 173382 606454
rect 172826 605898 173062 606134
rect 173146 605898 173382 606134
rect 172826 570218 173062 570454
rect 173146 570218 173382 570454
rect 172826 569898 173062 570134
rect 173146 569898 173382 570134
rect 172826 534218 173062 534454
rect 173146 534218 173382 534454
rect 172826 533898 173062 534134
rect 173146 533898 173382 534134
rect 172826 498218 173062 498454
rect 173146 498218 173382 498454
rect 172826 497898 173062 498134
rect 173146 497898 173382 498134
rect 172826 462218 173062 462454
rect 173146 462218 173382 462454
rect 172826 461898 173062 462134
rect 173146 461898 173382 462134
rect 172826 426218 173062 426454
rect 173146 426218 173382 426454
rect 172826 425898 173062 426134
rect 173146 425898 173382 426134
rect 172826 390218 173062 390454
rect 173146 390218 173382 390454
rect 172826 389898 173062 390134
rect 173146 389898 173382 390134
rect 172826 354218 173062 354454
rect 173146 354218 173382 354454
rect 172826 353898 173062 354134
rect 173146 353898 173382 354134
rect 172826 318218 173062 318454
rect 173146 318218 173382 318454
rect 172826 317898 173062 318134
rect 173146 317898 173382 318134
rect 172826 282218 173062 282454
rect 173146 282218 173382 282454
rect 172826 281898 173062 282134
rect 173146 281898 173382 282134
rect 177326 711322 177562 711558
rect 177646 711322 177882 711558
rect 177326 711002 177562 711238
rect 177646 711002 177882 711238
rect 177326 682718 177562 682954
rect 177646 682718 177882 682954
rect 177326 682398 177562 682634
rect 177646 682398 177882 682634
rect 177326 646718 177562 646954
rect 177646 646718 177882 646954
rect 177326 646398 177562 646634
rect 177646 646398 177882 646634
rect 177326 610718 177562 610954
rect 177646 610718 177882 610954
rect 177326 610398 177562 610634
rect 177646 610398 177882 610634
rect 177326 574718 177562 574954
rect 177646 574718 177882 574954
rect 177326 574398 177562 574634
rect 177646 574398 177882 574634
rect 177326 538718 177562 538954
rect 177646 538718 177882 538954
rect 177326 538398 177562 538634
rect 177646 538398 177882 538634
rect 177326 502718 177562 502954
rect 177646 502718 177882 502954
rect 177326 502398 177562 502634
rect 177646 502398 177882 502634
rect 177326 466718 177562 466954
rect 177646 466718 177882 466954
rect 177326 466398 177562 466634
rect 177646 466398 177882 466634
rect 177326 430718 177562 430954
rect 177646 430718 177882 430954
rect 177326 430398 177562 430634
rect 177646 430398 177882 430634
rect 177326 394718 177562 394954
rect 177646 394718 177882 394954
rect 177326 394398 177562 394634
rect 177646 394398 177882 394634
rect 177326 358718 177562 358954
rect 177646 358718 177882 358954
rect 177326 358398 177562 358634
rect 177646 358398 177882 358634
rect 177326 322718 177562 322954
rect 177646 322718 177882 322954
rect 177326 322398 177562 322634
rect 177646 322398 177882 322634
rect 177326 286718 177562 286954
rect 177646 286718 177882 286954
rect 177326 286398 177562 286634
rect 177646 286398 177882 286634
rect 177326 250718 177562 250954
rect 177646 250718 177882 250954
rect 177326 250398 177562 250634
rect 177646 250398 177882 250634
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 186326 705562 186562 705798
rect 186646 705562 186882 705798
rect 186326 705242 186562 705478
rect 186646 705242 186882 705478
rect 186326 691718 186562 691954
rect 186646 691718 186882 691954
rect 186326 691398 186562 691634
rect 186646 691398 186882 691634
rect 186326 655718 186562 655954
rect 186646 655718 186882 655954
rect 186326 655398 186562 655634
rect 186646 655398 186882 655634
rect 186326 619718 186562 619954
rect 186646 619718 186882 619954
rect 186326 619398 186562 619634
rect 186646 619398 186882 619634
rect 186326 583718 186562 583954
rect 186646 583718 186882 583954
rect 186326 583398 186562 583634
rect 186646 583398 186882 583634
rect 186326 547718 186562 547954
rect 186646 547718 186882 547954
rect 186326 547398 186562 547634
rect 186646 547398 186882 547634
rect 186326 511718 186562 511954
rect 186646 511718 186882 511954
rect 186326 511398 186562 511634
rect 186646 511398 186882 511634
rect 186326 475718 186562 475954
rect 186646 475718 186882 475954
rect 186326 475398 186562 475634
rect 186646 475398 186882 475634
rect 186326 439718 186562 439954
rect 186646 439718 186882 439954
rect 186326 439398 186562 439634
rect 186646 439398 186882 439634
rect 186326 403718 186562 403954
rect 186646 403718 186882 403954
rect 186326 403398 186562 403634
rect 186646 403398 186882 403634
rect 186326 367718 186562 367954
rect 186646 367718 186882 367954
rect 186326 367398 186562 367634
rect 186646 367398 186882 367634
rect 186326 331718 186562 331954
rect 186646 331718 186882 331954
rect 186326 331398 186562 331634
rect 186646 331398 186882 331634
rect 186326 295718 186562 295954
rect 186646 295718 186882 295954
rect 186326 295398 186562 295634
rect 186646 295398 186882 295634
rect 186326 259718 186562 259954
rect 186646 259718 186882 259954
rect 186326 259398 186562 259634
rect 186646 259398 186882 259634
rect 190826 706522 191062 706758
rect 191146 706522 191382 706758
rect 190826 706202 191062 706438
rect 191146 706202 191382 706438
rect 190826 696218 191062 696454
rect 191146 696218 191382 696454
rect 190826 695898 191062 696134
rect 191146 695898 191382 696134
rect 190826 660218 191062 660454
rect 191146 660218 191382 660454
rect 190826 659898 191062 660134
rect 191146 659898 191382 660134
rect 190826 624218 191062 624454
rect 191146 624218 191382 624454
rect 190826 623898 191062 624134
rect 191146 623898 191382 624134
rect 190826 588218 191062 588454
rect 191146 588218 191382 588454
rect 190826 587898 191062 588134
rect 191146 587898 191382 588134
rect 190826 552218 191062 552454
rect 191146 552218 191382 552454
rect 190826 551898 191062 552134
rect 191146 551898 191382 552134
rect 190826 516218 191062 516454
rect 191146 516218 191382 516454
rect 190826 515898 191062 516134
rect 191146 515898 191382 516134
rect 190826 480218 191062 480454
rect 191146 480218 191382 480454
rect 190826 479898 191062 480134
rect 191146 479898 191382 480134
rect 190826 444218 191062 444454
rect 191146 444218 191382 444454
rect 190826 443898 191062 444134
rect 191146 443898 191382 444134
rect 190826 408218 191062 408454
rect 191146 408218 191382 408454
rect 190826 407898 191062 408134
rect 191146 407898 191382 408134
rect 190826 372218 191062 372454
rect 191146 372218 191382 372454
rect 190826 371898 191062 372134
rect 191146 371898 191382 372134
rect 190826 336218 191062 336454
rect 191146 336218 191382 336454
rect 190826 335898 191062 336134
rect 191146 335898 191382 336134
rect 190826 300218 191062 300454
rect 191146 300218 191382 300454
rect 190826 299898 191062 300134
rect 191146 299898 191382 300134
rect 190826 264218 191062 264454
rect 191146 264218 191382 264454
rect 190826 263898 191062 264134
rect 191146 263898 191382 264134
rect 195326 707482 195562 707718
rect 195646 707482 195882 707718
rect 195326 707162 195562 707398
rect 195646 707162 195882 707398
rect 195326 700718 195562 700954
rect 195646 700718 195882 700954
rect 195326 700398 195562 700634
rect 195646 700398 195882 700634
rect 195326 664718 195562 664954
rect 195646 664718 195882 664954
rect 195326 664398 195562 664634
rect 195646 664398 195882 664634
rect 195326 628718 195562 628954
rect 195646 628718 195882 628954
rect 195326 628398 195562 628634
rect 195646 628398 195882 628634
rect 195326 592718 195562 592954
rect 195646 592718 195882 592954
rect 195326 592398 195562 592634
rect 195646 592398 195882 592634
rect 195326 556718 195562 556954
rect 195646 556718 195882 556954
rect 195326 556398 195562 556634
rect 195646 556398 195882 556634
rect 195326 520718 195562 520954
rect 195646 520718 195882 520954
rect 195326 520398 195562 520634
rect 195646 520398 195882 520634
rect 195326 484718 195562 484954
rect 195646 484718 195882 484954
rect 195326 484398 195562 484634
rect 195646 484398 195882 484634
rect 195326 448718 195562 448954
rect 195646 448718 195882 448954
rect 195326 448398 195562 448634
rect 195646 448398 195882 448634
rect 195326 412718 195562 412954
rect 195646 412718 195882 412954
rect 195326 412398 195562 412634
rect 195646 412398 195882 412634
rect 195326 376718 195562 376954
rect 195646 376718 195882 376954
rect 195326 376398 195562 376634
rect 195646 376398 195882 376634
rect 195326 340718 195562 340954
rect 195646 340718 195882 340954
rect 195326 340398 195562 340634
rect 195646 340398 195882 340634
rect 195326 304718 195562 304954
rect 195646 304718 195882 304954
rect 195326 304398 195562 304634
rect 195646 304398 195882 304634
rect 195326 268718 195562 268954
rect 195646 268718 195882 268954
rect 195326 268398 195562 268634
rect 195646 268398 195882 268634
rect 199826 708442 200062 708678
rect 200146 708442 200382 708678
rect 199826 708122 200062 708358
rect 200146 708122 200382 708358
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 204326 709402 204562 709638
rect 204646 709402 204882 709638
rect 204326 709082 204562 709318
rect 204646 709082 204882 709318
rect 204326 673718 204562 673954
rect 204646 673718 204882 673954
rect 204326 673398 204562 673634
rect 204646 673398 204882 673634
rect 204326 637718 204562 637954
rect 204646 637718 204882 637954
rect 204326 637398 204562 637634
rect 204646 637398 204882 637634
rect 204326 601718 204562 601954
rect 204646 601718 204882 601954
rect 204326 601398 204562 601634
rect 204646 601398 204882 601634
rect 204326 565718 204562 565954
rect 204646 565718 204882 565954
rect 204326 565398 204562 565634
rect 204646 565398 204882 565634
rect 204326 529718 204562 529954
rect 204646 529718 204882 529954
rect 204326 529398 204562 529634
rect 204646 529398 204882 529634
rect 204326 493718 204562 493954
rect 204646 493718 204882 493954
rect 204326 493398 204562 493634
rect 204646 493398 204882 493634
rect 204326 457718 204562 457954
rect 204646 457718 204882 457954
rect 204326 457398 204562 457634
rect 204646 457398 204882 457634
rect 204326 421718 204562 421954
rect 204646 421718 204882 421954
rect 204326 421398 204562 421634
rect 204646 421398 204882 421634
rect 204326 385718 204562 385954
rect 204646 385718 204882 385954
rect 204326 385398 204562 385634
rect 204646 385398 204882 385634
rect 204326 349718 204562 349954
rect 204646 349718 204882 349954
rect 204326 349398 204562 349634
rect 204646 349398 204882 349634
rect 204326 313718 204562 313954
rect 204646 313718 204882 313954
rect 204326 313398 204562 313634
rect 204646 313398 204882 313634
rect 204326 277718 204562 277954
rect 204646 277718 204882 277954
rect 204326 277398 204562 277634
rect 204646 277398 204882 277634
rect 208826 710362 209062 710598
rect 209146 710362 209382 710598
rect 208826 710042 209062 710278
rect 209146 710042 209382 710278
rect 208826 678218 209062 678454
rect 209146 678218 209382 678454
rect 208826 677898 209062 678134
rect 209146 677898 209382 678134
rect 208826 642218 209062 642454
rect 209146 642218 209382 642454
rect 208826 641898 209062 642134
rect 209146 641898 209382 642134
rect 208826 606218 209062 606454
rect 209146 606218 209382 606454
rect 208826 605898 209062 606134
rect 209146 605898 209382 606134
rect 208826 570218 209062 570454
rect 209146 570218 209382 570454
rect 208826 569898 209062 570134
rect 209146 569898 209382 570134
rect 208826 534218 209062 534454
rect 209146 534218 209382 534454
rect 208826 533898 209062 534134
rect 209146 533898 209382 534134
rect 208826 498218 209062 498454
rect 209146 498218 209382 498454
rect 208826 497898 209062 498134
rect 209146 497898 209382 498134
rect 208826 462218 209062 462454
rect 209146 462218 209382 462454
rect 208826 461898 209062 462134
rect 209146 461898 209382 462134
rect 208826 426218 209062 426454
rect 209146 426218 209382 426454
rect 208826 425898 209062 426134
rect 209146 425898 209382 426134
rect 208826 390218 209062 390454
rect 209146 390218 209382 390454
rect 208826 389898 209062 390134
rect 209146 389898 209382 390134
rect 208826 354218 209062 354454
rect 209146 354218 209382 354454
rect 208826 353898 209062 354134
rect 209146 353898 209382 354134
rect 208826 318218 209062 318454
rect 209146 318218 209382 318454
rect 208826 317898 209062 318134
rect 209146 317898 209382 318134
rect 208826 282218 209062 282454
rect 209146 282218 209382 282454
rect 208826 281898 209062 282134
rect 209146 281898 209382 282134
rect 213326 711322 213562 711558
rect 213646 711322 213882 711558
rect 213326 711002 213562 711238
rect 213646 711002 213882 711238
rect 213326 682718 213562 682954
rect 213646 682718 213882 682954
rect 213326 682398 213562 682634
rect 213646 682398 213882 682634
rect 213326 646718 213562 646954
rect 213646 646718 213882 646954
rect 213326 646398 213562 646634
rect 213646 646398 213882 646634
rect 213326 610718 213562 610954
rect 213646 610718 213882 610954
rect 213326 610398 213562 610634
rect 213646 610398 213882 610634
rect 213326 574718 213562 574954
rect 213646 574718 213882 574954
rect 213326 574398 213562 574634
rect 213646 574398 213882 574634
rect 213326 538718 213562 538954
rect 213646 538718 213882 538954
rect 213326 538398 213562 538634
rect 213646 538398 213882 538634
rect 213326 502718 213562 502954
rect 213646 502718 213882 502954
rect 213326 502398 213562 502634
rect 213646 502398 213882 502634
rect 213326 466718 213562 466954
rect 213646 466718 213882 466954
rect 213326 466398 213562 466634
rect 213646 466398 213882 466634
rect 213326 430718 213562 430954
rect 213646 430718 213882 430954
rect 213326 430398 213562 430634
rect 213646 430398 213882 430634
rect 213326 394718 213562 394954
rect 213646 394718 213882 394954
rect 213326 394398 213562 394634
rect 213646 394398 213882 394634
rect 213326 358718 213562 358954
rect 213646 358718 213882 358954
rect 213326 358398 213562 358634
rect 213646 358398 213882 358634
rect 213326 322718 213562 322954
rect 213646 322718 213882 322954
rect 213326 322398 213562 322634
rect 213646 322398 213882 322634
rect 213326 286718 213562 286954
rect 213646 286718 213882 286954
rect 213326 286398 213562 286634
rect 213646 286398 213882 286634
rect 213326 250718 213562 250954
rect 213646 250718 213882 250954
rect 213326 250398 213562 250634
rect 213646 250398 213882 250634
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 222326 705562 222562 705798
rect 222646 705562 222882 705798
rect 222326 705242 222562 705478
rect 222646 705242 222882 705478
rect 222326 691718 222562 691954
rect 222646 691718 222882 691954
rect 222326 691398 222562 691634
rect 222646 691398 222882 691634
rect 222326 655718 222562 655954
rect 222646 655718 222882 655954
rect 222326 655398 222562 655634
rect 222646 655398 222882 655634
rect 222326 619718 222562 619954
rect 222646 619718 222882 619954
rect 222326 619398 222562 619634
rect 222646 619398 222882 619634
rect 222326 583718 222562 583954
rect 222646 583718 222882 583954
rect 222326 583398 222562 583634
rect 222646 583398 222882 583634
rect 222326 547718 222562 547954
rect 222646 547718 222882 547954
rect 222326 547398 222562 547634
rect 222646 547398 222882 547634
rect 222326 511718 222562 511954
rect 222646 511718 222882 511954
rect 222326 511398 222562 511634
rect 222646 511398 222882 511634
rect 222326 475718 222562 475954
rect 222646 475718 222882 475954
rect 222326 475398 222562 475634
rect 222646 475398 222882 475634
rect 222326 439718 222562 439954
rect 222646 439718 222882 439954
rect 222326 439398 222562 439634
rect 222646 439398 222882 439634
rect 222326 403718 222562 403954
rect 222646 403718 222882 403954
rect 222326 403398 222562 403634
rect 222646 403398 222882 403634
rect 222326 367718 222562 367954
rect 222646 367718 222882 367954
rect 222326 367398 222562 367634
rect 222646 367398 222882 367634
rect 222326 331718 222562 331954
rect 222646 331718 222882 331954
rect 222326 331398 222562 331634
rect 222646 331398 222882 331634
rect 222326 295718 222562 295954
rect 222646 295718 222882 295954
rect 222326 295398 222562 295634
rect 222646 295398 222882 295634
rect 222326 259718 222562 259954
rect 222646 259718 222882 259954
rect 222326 259398 222562 259634
rect 222646 259398 222882 259634
rect 226826 706522 227062 706758
rect 227146 706522 227382 706758
rect 226826 706202 227062 706438
rect 227146 706202 227382 706438
rect 226826 696218 227062 696454
rect 227146 696218 227382 696454
rect 226826 695898 227062 696134
rect 227146 695898 227382 696134
rect 226826 660218 227062 660454
rect 227146 660218 227382 660454
rect 226826 659898 227062 660134
rect 227146 659898 227382 660134
rect 226826 624218 227062 624454
rect 227146 624218 227382 624454
rect 226826 623898 227062 624134
rect 227146 623898 227382 624134
rect 226826 588218 227062 588454
rect 227146 588218 227382 588454
rect 226826 587898 227062 588134
rect 227146 587898 227382 588134
rect 226826 552218 227062 552454
rect 227146 552218 227382 552454
rect 226826 551898 227062 552134
rect 227146 551898 227382 552134
rect 226826 516218 227062 516454
rect 227146 516218 227382 516454
rect 226826 515898 227062 516134
rect 227146 515898 227382 516134
rect 226826 480218 227062 480454
rect 227146 480218 227382 480454
rect 226826 479898 227062 480134
rect 227146 479898 227382 480134
rect 226826 444218 227062 444454
rect 227146 444218 227382 444454
rect 226826 443898 227062 444134
rect 227146 443898 227382 444134
rect 226826 408218 227062 408454
rect 227146 408218 227382 408454
rect 226826 407898 227062 408134
rect 227146 407898 227382 408134
rect 226826 372218 227062 372454
rect 227146 372218 227382 372454
rect 226826 371898 227062 372134
rect 227146 371898 227382 372134
rect 226826 336218 227062 336454
rect 227146 336218 227382 336454
rect 226826 335898 227062 336134
rect 227146 335898 227382 336134
rect 226826 300218 227062 300454
rect 227146 300218 227382 300454
rect 226826 299898 227062 300134
rect 227146 299898 227382 300134
rect 226826 264218 227062 264454
rect 227146 264218 227382 264454
rect 226826 263898 227062 264134
rect 227146 263898 227382 264134
rect 231326 707482 231562 707718
rect 231646 707482 231882 707718
rect 231326 707162 231562 707398
rect 231646 707162 231882 707398
rect 231326 700718 231562 700954
rect 231646 700718 231882 700954
rect 231326 700398 231562 700634
rect 231646 700398 231882 700634
rect 231326 664718 231562 664954
rect 231646 664718 231882 664954
rect 231326 664398 231562 664634
rect 231646 664398 231882 664634
rect 231326 628718 231562 628954
rect 231646 628718 231882 628954
rect 231326 628398 231562 628634
rect 231646 628398 231882 628634
rect 231326 592718 231562 592954
rect 231646 592718 231882 592954
rect 231326 592398 231562 592634
rect 231646 592398 231882 592634
rect 231326 556718 231562 556954
rect 231646 556718 231882 556954
rect 231326 556398 231562 556634
rect 231646 556398 231882 556634
rect 231326 520718 231562 520954
rect 231646 520718 231882 520954
rect 231326 520398 231562 520634
rect 231646 520398 231882 520634
rect 231326 484718 231562 484954
rect 231646 484718 231882 484954
rect 231326 484398 231562 484634
rect 231646 484398 231882 484634
rect 231326 448718 231562 448954
rect 231646 448718 231882 448954
rect 231326 448398 231562 448634
rect 231646 448398 231882 448634
rect 231326 412718 231562 412954
rect 231646 412718 231882 412954
rect 231326 412398 231562 412634
rect 231646 412398 231882 412634
rect 231326 376718 231562 376954
rect 231646 376718 231882 376954
rect 231326 376398 231562 376634
rect 231646 376398 231882 376634
rect 231326 340718 231562 340954
rect 231646 340718 231882 340954
rect 231326 340398 231562 340634
rect 231646 340398 231882 340634
rect 231326 304718 231562 304954
rect 231646 304718 231882 304954
rect 231326 304398 231562 304634
rect 231646 304398 231882 304634
rect 231326 268718 231562 268954
rect 231646 268718 231882 268954
rect 231326 268398 231562 268634
rect 231646 268398 231882 268634
rect 235826 708442 236062 708678
rect 236146 708442 236382 708678
rect 235826 708122 236062 708358
rect 236146 708122 236382 708358
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 235826 273218 236062 273454
rect 236146 273218 236382 273454
rect 235826 272898 236062 273134
rect 236146 272898 236382 273134
rect 240326 709402 240562 709638
rect 240646 709402 240882 709638
rect 240326 709082 240562 709318
rect 240646 709082 240882 709318
rect 240326 673718 240562 673954
rect 240646 673718 240882 673954
rect 240326 673398 240562 673634
rect 240646 673398 240882 673634
rect 240326 637718 240562 637954
rect 240646 637718 240882 637954
rect 240326 637398 240562 637634
rect 240646 637398 240882 637634
rect 240326 601718 240562 601954
rect 240646 601718 240882 601954
rect 240326 601398 240562 601634
rect 240646 601398 240882 601634
rect 240326 565718 240562 565954
rect 240646 565718 240882 565954
rect 240326 565398 240562 565634
rect 240646 565398 240882 565634
rect 240326 529718 240562 529954
rect 240646 529718 240882 529954
rect 240326 529398 240562 529634
rect 240646 529398 240882 529634
rect 240326 493718 240562 493954
rect 240646 493718 240882 493954
rect 240326 493398 240562 493634
rect 240646 493398 240882 493634
rect 240326 457718 240562 457954
rect 240646 457718 240882 457954
rect 240326 457398 240562 457634
rect 240646 457398 240882 457634
rect 240326 421718 240562 421954
rect 240646 421718 240882 421954
rect 240326 421398 240562 421634
rect 240646 421398 240882 421634
rect 240326 385718 240562 385954
rect 240646 385718 240882 385954
rect 240326 385398 240562 385634
rect 240646 385398 240882 385634
rect 240326 349718 240562 349954
rect 240646 349718 240882 349954
rect 240326 349398 240562 349634
rect 240646 349398 240882 349634
rect 240326 313718 240562 313954
rect 240646 313718 240882 313954
rect 240326 313398 240562 313634
rect 240646 313398 240882 313634
rect 240326 277718 240562 277954
rect 240646 277718 240882 277954
rect 240326 277398 240562 277634
rect 240646 277398 240882 277634
rect 244826 710362 245062 710598
rect 245146 710362 245382 710598
rect 244826 710042 245062 710278
rect 245146 710042 245382 710278
rect 244826 678218 245062 678454
rect 245146 678218 245382 678454
rect 244826 677898 245062 678134
rect 245146 677898 245382 678134
rect 244826 642218 245062 642454
rect 245146 642218 245382 642454
rect 244826 641898 245062 642134
rect 245146 641898 245382 642134
rect 244826 606218 245062 606454
rect 245146 606218 245382 606454
rect 244826 605898 245062 606134
rect 245146 605898 245382 606134
rect 244826 570218 245062 570454
rect 245146 570218 245382 570454
rect 244826 569898 245062 570134
rect 245146 569898 245382 570134
rect 244826 534218 245062 534454
rect 245146 534218 245382 534454
rect 244826 533898 245062 534134
rect 245146 533898 245382 534134
rect 244826 498218 245062 498454
rect 245146 498218 245382 498454
rect 244826 497898 245062 498134
rect 245146 497898 245382 498134
rect 244826 462218 245062 462454
rect 245146 462218 245382 462454
rect 244826 461898 245062 462134
rect 245146 461898 245382 462134
rect 244826 426218 245062 426454
rect 245146 426218 245382 426454
rect 244826 425898 245062 426134
rect 245146 425898 245382 426134
rect 244826 390218 245062 390454
rect 245146 390218 245382 390454
rect 244826 389898 245062 390134
rect 245146 389898 245382 390134
rect 244826 354218 245062 354454
rect 245146 354218 245382 354454
rect 244826 353898 245062 354134
rect 245146 353898 245382 354134
rect 244826 318218 245062 318454
rect 245146 318218 245382 318454
rect 244826 317898 245062 318134
rect 245146 317898 245382 318134
rect 244826 282218 245062 282454
rect 245146 282218 245382 282454
rect 244826 281898 245062 282134
rect 245146 281898 245382 282134
rect 249326 711322 249562 711558
rect 249646 711322 249882 711558
rect 249326 711002 249562 711238
rect 249646 711002 249882 711238
rect 249326 682718 249562 682954
rect 249646 682718 249882 682954
rect 249326 682398 249562 682634
rect 249646 682398 249882 682634
rect 249326 646718 249562 646954
rect 249646 646718 249882 646954
rect 249326 646398 249562 646634
rect 249646 646398 249882 646634
rect 249326 610718 249562 610954
rect 249646 610718 249882 610954
rect 249326 610398 249562 610634
rect 249646 610398 249882 610634
rect 249326 574718 249562 574954
rect 249646 574718 249882 574954
rect 249326 574398 249562 574634
rect 249646 574398 249882 574634
rect 249326 538718 249562 538954
rect 249646 538718 249882 538954
rect 249326 538398 249562 538634
rect 249646 538398 249882 538634
rect 249326 502718 249562 502954
rect 249646 502718 249882 502954
rect 249326 502398 249562 502634
rect 249646 502398 249882 502634
rect 249326 466718 249562 466954
rect 249646 466718 249882 466954
rect 249326 466398 249562 466634
rect 249646 466398 249882 466634
rect 249326 430718 249562 430954
rect 249646 430718 249882 430954
rect 249326 430398 249562 430634
rect 249646 430398 249882 430634
rect 249326 394718 249562 394954
rect 249646 394718 249882 394954
rect 249326 394398 249562 394634
rect 249646 394398 249882 394634
rect 249326 358718 249562 358954
rect 249646 358718 249882 358954
rect 249326 358398 249562 358634
rect 249646 358398 249882 358634
rect 249326 322718 249562 322954
rect 249646 322718 249882 322954
rect 249326 322398 249562 322634
rect 249646 322398 249882 322634
rect 249326 286718 249562 286954
rect 249646 286718 249882 286954
rect 249326 286398 249562 286634
rect 249646 286398 249882 286634
rect 249326 250718 249562 250954
rect 249646 250718 249882 250954
rect 249326 250398 249562 250634
rect 249646 250398 249882 250634
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 258326 705562 258562 705798
rect 258646 705562 258882 705798
rect 258326 705242 258562 705478
rect 258646 705242 258882 705478
rect 258326 691718 258562 691954
rect 258646 691718 258882 691954
rect 258326 691398 258562 691634
rect 258646 691398 258882 691634
rect 258326 655718 258562 655954
rect 258646 655718 258882 655954
rect 258326 655398 258562 655634
rect 258646 655398 258882 655634
rect 258326 619718 258562 619954
rect 258646 619718 258882 619954
rect 258326 619398 258562 619634
rect 258646 619398 258882 619634
rect 258326 583718 258562 583954
rect 258646 583718 258882 583954
rect 258326 583398 258562 583634
rect 258646 583398 258882 583634
rect 258326 547718 258562 547954
rect 258646 547718 258882 547954
rect 258326 547398 258562 547634
rect 258646 547398 258882 547634
rect 258326 511718 258562 511954
rect 258646 511718 258882 511954
rect 258326 511398 258562 511634
rect 258646 511398 258882 511634
rect 258326 475718 258562 475954
rect 258646 475718 258882 475954
rect 258326 475398 258562 475634
rect 258646 475398 258882 475634
rect 258326 439718 258562 439954
rect 258646 439718 258882 439954
rect 258326 439398 258562 439634
rect 258646 439398 258882 439634
rect 258326 403718 258562 403954
rect 258646 403718 258882 403954
rect 258326 403398 258562 403634
rect 258646 403398 258882 403634
rect 258326 367718 258562 367954
rect 258646 367718 258882 367954
rect 258326 367398 258562 367634
rect 258646 367398 258882 367634
rect 258326 331718 258562 331954
rect 258646 331718 258882 331954
rect 258326 331398 258562 331634
rect 258646 331398 258882 331634
rect 258326 295718 258562 295954
rect 258646 295718 258882 295954
rect 258326 295398 258562 295634
rect 258646 295398 258882 295634
rect 258326 259718 258562 259954
rect 258646 259718 258882 259954
rect 258326 259398 258562 259634
rect 258646 259398 258882 259634
rect 262826 706522 263062 706758
rect 263146 706522 263382 706758
rect 262826 706202 263062 706438
rect 263146 706202 263382 706438
rect 262826 696218 263062 696454
rect 263146 696218 263382 696454
rect 262826 695898 263062 696134
rect 263146 695898 263382 696134
rect 262826 660218 263062 660454
rect 263146 660218 263382 660454
rect 262826 659898 263062 660134
rect 263146 659898 263382 660134
rect 262826 624218 263062 624454
rect 263146 624218 263382 624454
rect 262826 623898 263062 624134
rect 263146 623898 263382 624134
rect 262826 588218 263062 588454
rect 263146 588218 263382 588454
rect 262826 587898 263062 588134
rect 263146 587898 263382 588134
rect 262826 552218 263062 552454
rect 263146 552218 263382 552454
rect 262826 551898 263062 552134
rect 263146 551898 263382 552134
rect 262826 516218 263062 516454
rect 263146 516218 263382 516454
rect 262826 515898 263062 516134
rect 263146 515898 263382 516134
rect 262826 480218 263062 480454
rect 263146 480218 263382 480454
rect 262826 479898 263062 480134
rect 263146 479898 263382 480134
rect 262826 444218 263062 444454
rect 263146 444218 263382 444454
rect 262826 443898 263062 444134
rect 263146 443898 263382 444134
rect 262826 408218 263062 408454
rect 263146 408218 263382 408454
rect 262826 407898 263062 408134
rect 263146 407898 263382 408134
rect 262826 372218 263062 372454
rect 263146 372218 263382 372454
rect 262826 371898 263062 372134
rect 263146 371898 263382 372134
rect 262826 336218 263062 336454
rect 263146 336218 263382 336454
rect 262826 335898 263062 336134
rect 263146 335898 263382 336134
rect 262826 300218 263062 300454
rect 263146 300218 263382 300454
rect 262826 299898 263062 300134
rect 263146 299898 263382 300134
rect 262826 264218 263062 264454
rect 263146 264218 263382 264454
rect 262826 263898 263062 264134
rect 263146 263898 263382 264134
rect 267326 707482 267562 707718
rect 267646 707482 267882 707718
rect 267326 707162 267562 707398
rect 267646 707162 267882 707398
rect 267326 700718 267562 700954
rect 267646 700718 267882 700954
rect 267326 700398 267562 700634
rect 267646 700398 267882 700634
rect 267326 664718 267562 664954
rect 267646 664718 267882 664954
rect 267326 664398 267562 664634
rect 267646 664398 267882 664634
rect 267326 628718 267562 628954
rect 267646 628718 267882 628954
rect 267326 628398 267562 628634
rect 267646 628398 267882 628634
rect 267326 592718 267562 592954
rect 267646 592718 267882 592954
rect 267326 592398 267562 592634
rect 267646 592398 267882 592634
rect 267326 556718 267562 556954
rect 267646 556718 267882 556954
rect 267326 556398 267562 556634
rect 267646 556398 267882 556634
rect 267326 520718 267562 520954
rect 267646 520718 267882 520954
rect 267326 520398 267562 520634
rect 267646 520398 267882 520634
rect 267326 484718 267562 484954
rect 267646 484718 267882 484954
rect 267326 484398 267562 484634
rect 267646 484398 267882 484634
rect 267326 448718 267562 448954
rect 267646 448718 267882 448954
rect 267326 448398 267562 448634
rect 267646 448398 267882 448634
rect 267326 412718 267562 412954
rect 267646 412718 267882 412954
rect 267326 412398 267562 412634
rect 267646 412398 267882 412634
rect 267326 376718 267562 376954
rect 267646 376718 267882 376954
rect 267326 376398 267562 376634
rect 267646 376398 267882 376634
rect 267326 340718 267562 340954
rect 267646 340718 267882 340954
rect 267326 340398 267562 340634
rect 267646 340398 267882 340634
rect 267326 304718 267562 304954
rect 267646 304718 267882 304954
rect 267326 304398 267562 304634
rect 267646 304398 267882 304634
rect 267326 268718 267562 268954
rect 267646 268718 267882 268954
rect 267326 268398 267562 268634
rect 267646 268398 267882 268634
rect 271826 708442 272062 708678
rect 272146 708442 272382 708678
rect 271826 708122 272062 708358
rect 272146 708122 272382 708358
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 276326 709402 276562 709638
rect 276646 709402 276882 709638
rect 276326 709082 276562 709318
rect 276646 709082 276882 709318
rect 276326 673718 276562 673954
rect 276646 673718 276882 673954
rect 276326 673398 276562 673634
rect 276646 673398 276882 673634
rect 276326 637718 276562 637954
rect 276646 637718 276882 637954
rect 276326 637398 276562 637634
rect 276646 637398 276882 637634
rect 276326 601718 276562 601954
rect 276646 601718 276882 601954
rect 276326 601398 276562 601634
rect 276646 601398 276882 601634
rect 276326 565718 276562 565954
rect 276646 565718 276882 565954
rect 276326 565398 276562 565634
rect 276646 565398 276882 565634
rect 276326 529718 276562 529954
rect 276646 529718 276882 529954
rect 276326 529398 276562 529634
rect 276646 529398 276882 529634
rect 276326 493718 276562 493954
rect 276646 493718 276882 493954
rect 276326 493398 276562 493634
rect 276646 493398 276882 493634
rect 276326 457718 276562 457954
rect 276646 457718 276882 457954
rect 276326 457398 276562 457634
rect 276646 457398 276882 457634
rect 276326 421718 276562 421954
rect 276646 421718 276882 421954
rect 276326 421398 276562 421634
rect 276646 421398 276882 421634
rect 276326 385718 276562 385954
rect 276646 385718 276882 385954
rect 276326 385398 276562 385634
rect 276646 385398 276882 385634
rect 276326 349718 276562 349954
rect 276646 349718 276882 349954
rect 276326 349398 276562 349634
rect 276646 349398 276882 349634
rect 276326 313718 276562 313954
rect 276646 313718 276882 313954
rect 276326 313398 276562 313634
rect 276646 313398 276882 313634
rect 276326 277718 276562 277954
rect 276646 277718 276882 277954
rect 276326 277398 276562 277634
rect 276646 277398 276882 277634
rect 280826 710362 281062 710598
rect 281146 710362 281382 710598
rect 280826 710042 281062 710278
rect 281146 710042 281382 710278
rect 280826 678218 281062 678454
rect 281146 678218 281382 678454
rect 280826 677898 281062 678134
rect 281146 677898 281382 678134
rect 280826 642218 281062 642454
rect 281146 642218 281382 642454
rect 280826 641898 281062 642134
rect 281146 641898 281382 642134
rect 280826 606218 281062 606454
rect 281146 606218 281382 606454
rect 280826 605898 281062 606134
rect 281146 605898 281382 606134
rect 280826 570218 281062 570454
rect 281146 570218 281382 570454
rect 280826 569898 281062 570134
rect 281146 569898 281382 570134
rect 280826 534218 281062 534454
rect 281146 534218 281382 534454
rect 280826 533898 281062 534134
rect 281146 533898 281382 534134
rect 280826 498218 281062 498454
rect 281146 498218 281382 498454
rect 280826 497898 281062 498134
rect 281146 497898 281382 498134
rect 280826 462218 281062 462454
rect 281146 462218 281382 462454
rect 280826 461898 281062 462134
rect 281146 461898 281382 462134
rect 280826 426218 281062 426454
rect 281146 426218 281382 426454
rect 280826 425898 281062 426134
rect 281146 425898 281382 426134
rect 280826 390218 281062 390454
rect 281146 390218 281382 390454
rect 280826 389898 281062 390134
rect 281146 389898 281382 390134
rect 280826 354218 281062 354454
rect 281146 354218 281382 354454
rect 280826 353898 281062 354134
rect 281146 353898 281382 354134
rect 280826 318218 281062 318454
rect 281146 318218 281382 318454
rect 280826 317898 281062 318134
rect 281146 317898 281382 318134
rect 280826 282218 281062 282454
rect 281146 282218 281382 282454
rect 280826 281898 281062 282134
rect 281146 281898 281382 282134
rect 285326 711322 285562 711558
rect 285646 711322 285882 711558
rect 285326 711002 285562 711238
rect 285646 711002 285882 711238
rect 285326 682718 285562 682954
rect 285646 682718 285882 682954
rect 285326 682398 285562 682634
rect 285646 682398 285882 682634
rect 285326 646718 285562 646954
rect 285646 646718 285882 646954
rect 285326 646398 285562 646634
rect 285646 646398 285882 646634
rect 285326 610718 285562 610954
rect 285646 610718 285882 610954
rect 285326 610398 285562 610634
rect 285646 610398 285882 610634
rect 285326 574718 285562 574954
rect 285646 574718 285882 574954
rect 285326 574398 285562 574634
rect 285646 574398 285882 574634
rect 285326 538718 285562 538954
rect 285646 538718 285882 538954
rect 285326 538398 285562 538634
rect 285646 538398 285882 538634
rect 285326 502718 285562 502954
rect 285646 502718 285882 502954
rect 285326 502398 285562 502634
rect 285646 502398 285882 502634
rect 285326 466718 285562 466954
rect 285646 466718 285882 466954
rect 285326 466398 285562 466634
rect 285646 466398 285882 466634
rect 285326 430718 285562 430954
rect 285646 430718 285882 430954
rect 285326 430398 285562 430634
rect 285646 430398 285882 430634
rect 285326 394718 285562 394954
rect 285646 394718 285882 394954
rect 285326 394398 285562 394634
rect 285646 394398 285882 394634
rect 285326 358718 285562 358954
rect 285646 358718 285882 358954
rect 285326 358398 285562 358634
rect 285646 358398 285882 358634
rect 285326 322718 285562 322954
rect 285646 322718 285882 322954
rect 285326 322398 285562 322634
rect 285646 322398 285882 322634
rect 285326 286718 285562 286954
rect 285646 286718 285882 286954
rect 285326 286398 285562 286634
rect 285646 286398 285882 286634
rect 285326 250718 285562 250954
rect 285646 250718 285882 250954
rect 285326 250398 285562 250634
rect 285646 250398 285882 250634
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 294326 705562 294562 705798
rect 294646 705562 294882 705798
rect 294326 705242 294562 705478
rect 294646 705242 294882 705478
rect 294326 691718 294562 691954
rect 294646 691718 294882 691954
rect 294326 691398 294562 691634
rect 294646 691398 294882 691634
rect 294326 655718 294562 655954
rect 294646 655718 294882 655954
rect 294326 655398 294562 655634
rect 294646 655398 294882 655634
rect 294326 619718 294562 619954
rect 294646 619718 294882 619954
rect 294326 619398 294562 619634
rect 294646 619398 294882 619634
rect 294326 583718 294562 583954
rect 294646 583718 294882 583954
rect 294326 583398 294562 583634
rect 294646 583398 294882 583634
rect 294326 547718 294562 547954
rect 294646 547718 294882 547954
rect 294326 547398 294562 547634
rect 294646 547398 294882 547634
rect 294326 511718 294562 511954
rect 294646 511718 294882 511954
rect 294326 511398 294562 511634
rect 294646 511398 294882 511634
rect 294326 475718 294562 475954
rect 294646 475718 294882 475954
rect 294326 475398 294562 475634
rect 294646 475398 294882 475634
rect 294326 439718 294562 439954
rect 294646 439718 294882 439954
rect 294326 439398 294562 439634
rect 294646 439398 294882 439634
rect 294326 403718 294562 403954
rect 294646 403718 294882 403954
rect 294326 403398 294562 403634
rect 294646 403398 294882 403634
rect 294326 367718 294562 367954
rect 294646 367718 294882 367954
rect 294326 367398 294562 367634
rect 294646 367398 294882 367634
rect 294326 331718 294562 331954
rect 294646 331718 294882 331954
rect 294326 331398 294562 331634
rect 294646 331398 294882 331634
rect 294326 295718 294562 295954
rect 294646 295718 294882 295954
rect 294326 295398 294562 295634
rect 294646 295398 294882 295634
rect 294326 259718 294562 259954
rect 294646 259718 294882 259954
rect 294326 259398 294562 259634
rect 294646 259398 294882 259634
rect 298826 706522 299062 706758
rect 299146 706522 299382 706758
rect 298826 706202 299062 706438
rect 299146 706202 299382 706438
rect 298826 696218 299062 696454
rect 299146 696218 299382 696454
rect 298826 695898 299062 696134
rect 299146 695898 299382 696134
rect 298826 660218 299062 660454
rect 299146 660218 299382 660454
rect 298826 659898 299062 660134
rect 299146 659898 299382 660134
rect 298826 624218 299062 624454
rect 299146 624218 299382 624454
rect 298826 623898 299062 624134
rect 299146 623898 299382 624134
rect 298826 588218 299062 588454
rect 299146 588218 299382 588454
rect 298826 587898 299062 588134
rect 299146 587898 299382 588134
rect 298826 552218 299062 552454
rect 299146 552218 299382 552454
rect 298826 551898 299062 552134
rect 299146 551898 299382 552134
rect 298826 516218 299062 516454
rect 299146 516218 299382 516454
rect 298826 515898 299062 516134
rect 299146 515898 299382 516134
rect 298826 480218 299062 480454
rect 299146 480218 299382 480454
rect 298826 479898 299062 480134
rect 299146 479898 299382 480134
rect 298826 444218 299062 444454
rect 299146 444218 299382 444454
rect 298826 443898 299062 444134
rect 299146 443898 299382 444134
rect 298826 408218 299062 408454
rect 299146 408218 299382 408454
rect 298826 407898 299062 408134
rect 299146 407898 299382 408134
rect 298826 372218 299062 372454
rect 299146 372218 299382 372454
rect 298826 371898 299062 372134
rect 299146 371898 299382 372134
rect 298826 336218 299062 336454
rect 299146 336218 299382 336454
rect 298826 335898 299062 336134
rect 299146 335898 299382 336134
rect 298826 300218 299062 300454
rect 299146 300218 299382 300454
rect 298826 299898 299062 300134
rect 299146 299898 299382 300134
rect 298826 264218 299062 264454
rect 299146 264218 299382 264454
rect 298826 263898 299062 264134
rect 299146 263898 299382 264134
rect 303326 707482 303562 707718
rect 303646 707482 303882 707718
rect 303326 707162 303562 707398
rect 303646 707162 303882 707398
rect 303326 700718 303562 700954
rect 303646 700718 303882 700954
rect 303326 700398 303562 700634
rect 303646 700398 303882 700634
rect 303326 664718 303562 664954
rect 303646 664718 303882 664954
rect 303326 664398 303562 664634
rect 303646 664398 303882 664634
rect 303326 628718 303562 628954
rect 303646 628718 303882 628954
rect 303326 628398 303562 628634
rect 303646 628398 303882 628634
rect 303326 592718 303562 592954
rect 303646 592718 303882 592954
rect 303326 592398 303562 592634
rect 303646 592398 303882 592634
rect 303326 556718 303562 556954
rect 303646 556718 303882 556954
rect 303326 556398 303562 556634
rect 303646 556398 303882 556634
rect 303326 520718 303562 520954
rect 303646 520718 303882 520954
rect 303326 520398 303562 520634
rect 303646 520398 303882 520634
rect 303326 484718 303562 484954
rect 303646 484718 303882 484954
rect 303326 484398 303562 484634
rect 303646 484398 303882 484634
rect 303326 448718 303562 448954
rect 303646 448718 303882 448954
rect 303326 448398 303562 448634
rect 303646 448398 303882 448634
rect 303326 412718 303562 412954
rect 303646 412718 303882 412954
rect 303326 412398 303562 412634
rect 303646 412398 303882 412634
rect 303326 376718 303562 376954
rect 303646 376718 303882 376954
rect 303326 376398 303562 376634
rect 303646 376398 303882 376634
rect 303326 340718 303562 340954
rect 303646 340718 303882 340954
rect 303326 340398 303562 340634
rect 303646 340398 303882 340634
rect 303326 304718 303562 304954
rect 303646 304718 303882 304954
rect 303326 304398 303562 304634
rect 303646 304398 303882 304634
rect 303326 268718 303562 268954
rect 303646 268718 303882 268954
rect 303326 268398 303562 268634
rect 303646 268398 303882 268634
rect 307826 708442 308062 708678
rect 308146 708442 308382 708678
rect 307826 708122 308062 708358
rect 308146 708122 308382 708358
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 312326 709402 312562 709638
rect 312646 709402 312882 709638
rect 312326 709082 312562 709318
rect 312646 709082 312882 709318
rect 312326 673718 312562 673954
rect 312646 673718 312882 673954
rect 312326 673398 312562 673634
rect 312646 673398 312882 673634
rect 312326 637718 312562 637954
rect 312646 637718 312882 637954
rect 312326 637398 312562 637634
rect 312646 637398 312882 637634
rect 312326 601718 312562 601954
rect 312646 601718 312882 601954
rect 312326 601398 312562 601634
rect 312646 601398 312882 601634
rect 312326 565718 312562 565954
rect 312646 565718 312882 565954
rect 312326 565398 312562 565634
rect 312646 565398 312882 565634
rect 312326 529718 312562 529954
rect 312646 529718 312882 529954
rect 312326 529398 312562 529634
rect 312646 529398 312882 529634
rect 312326 493718 312562 493954
rect 312646 493718 312882 493954
rect 312326 493398 312562 493634
rect 312646 493398 312882 493634
rect 312326 457718 312562 457954
rect 312646 457718 312882 457954
rect 312326 457398 312562 457634
rect 312646 457398 312882 457634
rect 312326 421718 312562 421954
rect 312646 421718 312882 421954
rect 312326 421398 312562 421634
rect 312646 421398 312882 421634
rect 312326 385718 312562 385954
rect 312646 385718 312882 385954
rect 312326 385398 312562 385634
rect 312646 385398 312882 385634
rect 312326 349718 312562 349954
rect 312646 349718 312882 349954
rect 312326 349398 312562 349634
rect 312646 349398 312882 349634
rect 312326 313718 312562 313954
rect 312646 313718 312882 313954
rect 312326 313398 312562 313634
rect 312646 313398 312882 313634
rect 312326 277718 312562 277954
rect 312646 277718 312882 277954
rect 312326 277398 312562 277634
rect 312646 277398 312882 277634
rect 316826 710362 317062 710598
rect 317146 710362 317382 710598
rect 316826 710042 317062 710278
rect 317146 710042 317382 710278
rect 316826 678218 317062 678454
rect 317146 678218 317382 678454
rect 316826 677898 317062 678134
rect 317146 677898 317382 678134
rect 316826 642218 317062 642454
rect 317146 642218 317382 642454
rect 316826 641898 317062 642134
rect 317146 641898 317382 642134
rect 316826 606218 317062 606454
rect 317146 606218 317382 606454
rect 316826 605898 317062 606134
rect 317146 605898 317382 606134
rect 316826 570218 317062 570454
rect 317146 570218 317382 570454
rect 316826 569898 317062 570134
rect 317146 569898 317382 570134
rect 316826 534218 317062 534454
rect 317146 534218 317382 534454
rect 316826 533898 317062 534134
rect 317146 533898 317382 534134
rect 316826 498218 317062 498454
rect 317146 498218 317382 498454
rect 316826 497898 317062 498134
rect 317146 497898 317382 498134
rect 316826 462218 317062 462454
rect 317146 462218 317382 462454
rect 316826 461898 317062 462134
rect 317146 461898 317382 462134
rect 316826 426218 317062 426454
rect 317146 426218 317382 426454
rect 316826 425898 317062 426134
rect 317146 425898 317382 426134
rect 316826 390218 317062 390454
rect 317146 390218 317382 390454
rect 316826 389898 317062 390134
rect 317146 389898 317382 390134
rect 316826 354218 317062 354454
rect 317146 354218 317382 354454
rect 316826 353898 317062 354134
rect 317146 353898 317382 354134
rect 316826 318218 317062 318454
rect 317146 318218 317382 318454
rect 316826 317898 317062 318134
rect 317146 317898 317382 318134
rect 316826 282218 317062 282454
rect 317146 282218 317382 282454
rect 316826 281898 317062 282134
rect 317146 281898 317382 282134
rect 321326 711322 321562 711558
rect 321646 711322 321882 711558
rect 321326 711002 321562 711238
rect 321646 711002 321882 711238
rect 321326 682718 321562 682954
rect 321646 682718 321882 682954
rect 321326 682398 321562 682634
rect 321646 682398 321882 682634
rect 321326 646718 321562 646954
rect 321646 646718 321882 646954
rect 321326 646398 321562 646634
rect 321646 646398 321882 646634
rect 321326 610718 321562 610954
rect 321646 610718 321882 610954
rect 321326 610398 321562 610634
rect 321646 610398 321882 610634
rect 321326 574718 321562 574954
rect 321646 574718 321882 574954
rect 321326 574398 321562 574634
rect 321646 574398 321882 574634
rect 321326 538718 321562 538954
rect 321646 538718 321882 538954
rect 321326 538398 321562 538634
rect 321646 538398 321882 538634
rect 321326 502718 321562 502954
rect 321646 502718 321882 502954
rect 321326 502398 321562 502634
rect 321646 502398 321882 502634
rect 321326 466718 321562 466954
rect 321646 466718 321882 466954
rect 321326 466398 321562 466634
rect 321646 466398 321882 466634
rect 321326 430718 321562 430954
rect 321646 430718 321882 430954
rect 321326 430398 321562 430634
rect 321646 430398 321882 430634
rect 321326 394718 321562 394954
rect 321646 394718 321882 394954
rect 321326 394398 321562 394634
rect 321646 394398 321882 394634
rect 321326 358718 321562 358954
rect 321646 358718 321882 358954
rect 321326 358398 321562 358634
rect 321646 358398 321882 358634
rect 321326 322718 321562 322954
rect 321646 322718 321882 322954
rect 321326 322398 321562 322634
rect 321646 322398 321882 322634
rect 321326 286718 321562 286954
rect 321646 286718 321882 286954
rect 321326 286398 321562 286634
rect 321646 286398 321882 286634
rect 321326 250718 321562 250954
rect 321646 250718 321882 250954
rect 321326 250398 321562 250634
rect 321646 250398 321882 250634
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 330326 705562 330562 705798
rect 330646 705562 330882 705798
rect 330326 705242 330562 705478
rect 330646 705242 330882 705478
rect 330326 691718 330562 691954
rect 330646 691718 330882 691954
rect 330326 691398 330562 691634
rect 330646 691398 330882 691634
rect 330326 655718 330562 655954
rect 330646 655718 330882 655954
rect 330326 655398 330562 655634
rect 330646 655398 330882 655634
rect 330326 619718 330562 619954
rect 330646 619718 330882 619954
rect 330326 619398 330562 619634
rect 330646 619398 330882 619634
rect 330326 583718 330562 583954
rect 330646 583718 330882 583954
rect 330326 583398 330562 583634
rect 330646 583398 330882 583634
rect 330326 547718 330562 547954
rect 330646 547718 330882 547954
rect 330326 547398 330562 547634
rect 330646 547398 330882 547634
rect 330326 511718 330562 511954
rect 330646 511718 330882 511954
rect 330326 511398 330562 511634
rect 330646 511398 330882 511634
rect 330326 475718 330562 475954
rect 330646 475718 330882 475954
rect 330326 475398 330562 475634
rect 330646 475398 330882 475634
rect 330326 439718 330562 439954
rect 330646 439718 330882 439954
rect 330326 439398 330562 439634
rect 330646 439398 330882 439634
rect 330326 403718 330562 403954
rect 330646 403718 330882 403954
rect 330326 403398 330562 403634
rect 330646 403398 330882 403634
rect 330326 367718 330562 367954
rect 330646 367718 330882 367954
rect 330326 367398 330562 367634
rect 330646 367398 330882 367634
rect 330326 331718 330562 331954
rect 330646 331718 330882 331954
rect 330326 331398 330562 331634
rect 330646 331398 330882 331634
rect 330326 295718 330562 295954
rect 330646 295718 330882 295954
rect 330326 295398 330562 295634
rect 330646 295398 330882 295634
rect 330326 259718 330562 259954
rect 330646 259718 330882 259954
rect 330326 259398 330562 259634
rect 330646 259398 330882 259634
rect 334826 706522 335062 706758
rect 335146 706522 335382 706758
rect 334826 706202 335062 706438
rect 335146 706202 335382 706438
rect 334826 696218 335062 696454
rect 335146 696218 335382 696454
rect 334826 695898 335062 696134
rect 335146 695898 335382 696134
rect 334826 660218 335062 660454
rect 335146 660218 335382 660454
rect 334826 659898 335062 660134
rect 335146 659898 335382 660134
rect 334826 624218 335062 624454
rect 335146 624218 335382 624454
rect 334826 623898 335062 624134
rect 335146 623898 335382 624134
rect 334826 588218 335062 588454
rect 335146 588218 335382 588454
rect 334826 587898 335062 588134
rect 335146 587898 335382 588134
rect 334826 552218 335062 552454
rect 335146 552218 335382 552454
rect 334826 551898 335062 552134
rect 335146 551898 335382 552134
rect 334826 516218 335062 516454
rect 335146 516218 335382 516454
rect 334826 515898 335062 516134
rect 335146 515898 335382 516134
rect 334826 480218 335062 480454
rect 335146 480218 335382 480454
rect 334826 479898 335062 480134
rect 335146 479898 335382 480134
rect 334826 444218 335062 444454
rect 335146 444218 335382 444454
rect 334826 443898 335062 444134
rect 335146 443898 335382 444134
rect 334826 408218 335062 408454
rect 335146 408218 335382 408454
rect 334826 407898 335062 408134
rect 335146 407898 335382 408134
rect 334826 372218 335062 372454
rect 335146 372218 335382 372454
rect 334826 371898 335062 372134
rect 335146 371898 335382 372134
rect 334826 336218 335062 336454
rect 335146 336218 335382 336454
rect 334826 335898 335062 336134
rect 335146 335898 335382 336134
rect 334826 300218 335062 300454
rect 335146 300218 335382 300454
rect 334826 299898 335062 300134
rect 335146 299898 335382 300134
rect 334826 264218 335062 264454
rect 335146 264218 335382 264454
rect 334826 263898 335062 264134
rect 335146 263898 335382 264134
rect 339326 707482 339562 707718
rect 339646 707482 339882 707718
rect 339326 707162 339562 707398
rect 339646 707162 339882 707398
rect 339326 700718 339562 700954
rect 339646 700718 339882 700954
rect 339326 700398 339562 700634
rect 339646 700398 339882 700634
rect 339326 664718 339562 664954
rect 339646 664718 339882 664954
rect 339326 664398 339562 664634
rect 339646 664398 339882 664634
rect 339326 628718 339562 628954
rect 339646 628718 339882 628954
rect 339326 628398 339562 628634
rect 339646 628398 339882 628634
rect 339326 592718 339562 592954
rect 339646 592718 339882 592954
rect 339326 592398 339562 592634
rect 339646 592398 339882 592634
rect 339326 556718 339562 556954
rect 339646 556718 339882 556954
rect 339326 556398 339562 556634
rect 339646 556398 339882 556634
rect 339326 520718 339562 520954
rect 339646 520718 339882 520954
rect 339326 520398 339562 520634
rect 339646 520398 339882 520634
rect 339326 484718 339562 484954
rect 339646 484718 339882 484954
rect 339326 484398 339562 484634
rect 339646 484398 339882 484634
rect 339326 448718 339562 448954
rect 339646 448718 339882 448954
rect 339326 448398 339562 448634
rect 339646 448398 339882 448634
rect 339326 412718 339562 412954
rect 339646 412718 339882 412954
rect 339326 412398 339562 412634
rect 339646 412398 339882 412634
rect 339326 376718 339562 376954
rect 339646 376718 339882 376954
rect 339326 376398 339562 376634
rect 339646 376398 339882 376634
rect 339326 340718 339562 340954
rect 339646 340718 339882 340954
rect 339326 340398 339562 340634
rect 339646 340398 339882 340634
rect 339326 304718 339562 304954
rect 339646 304718 339882 304954
rect 339326 304398 339562 304634
rect 339646 304398 339882 304634
rect 339326 268718 339562 268954
rect 339646 268718 339882 268954
rect 339326 268398 339562 268634
rect 339646 268398 339882 268634
rect 343826 708442 344062 708678
rect 344146 708442 344382 708678
rect 343826 708122 344062 708358
rect 344146 708122 344382 708358
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 348326 709402 348562 709638
rect 348646 709402 348882 709638
rect 348326 709082 348562 709318
rect 348646 709082 348882 709318
rect 348326 673718 348562 673954
rect 348646 673718 348882 673954
rect 348326 673398 348562 673634
rect 348646 673398 348882 673634
rect 348326 637718 348562 637954
rect 348646 637718 348882 637954
rect 348326 637398 348562 637634
rect 348646 637398 348882 637634
rect 348326 601718 348562 601954
rect 348646 601718 348882 601954
rect 348326 601398 348562 601634
rect 348646 601398 348882 601634
rect 348326 565718 348562 565954
rect 348646 565718 348882 565954
rect 348326 565398 348562 565634
rect 348646 565398 348882 565634
rect 348326 529718 348562 529954
rect 348646 529718 348882 529954
rect 348326 529398 348562 529634
rect 348646 529398 348882 529634
rect 348326 493718 348562 493954
rect 348646 493718 348882 493954
rect 348326 493398 348562 493634
rect 348646 493398 348882 493634
rect 348326 457718 348562 457954
rect 348646 457718 348882 457954
rect 348326 457398 348562 457634
rect 348646 457398 348882 457634
rect 348326 421718 348562 421954
rect 348646 421718 348882 421954
rect 348326 421398 348562 421634
rect 348646 421398 348882 421634
rect 348326 385718 348562 385954
rect 348646 385718 348882 385954
rect 348326 385398 348562 385634
rect 348646 385398 348882 385634
rect 348326 349718 348562 349954
rect 348646 349718 348882 349954
rect 348326 349398 348562 349634
rect 348646 349398 348882 349634
rect 348326 313718 348562 313954
rect 348646 313718 348882 313954
rect 348326 313398 348562 313634
rect 348646 313398 348882 313634
rect 348326 277718 348562 277954
rect 348646 277718 348882 277954
rect 348326 277398 348562 277634
rect 348646 277398 348882 277634
rect 352826 710362 353062 710598
rect 353146 710362 353382 710598
rect 352826 710042 353062 710278
rect 353146 710042 353382 710278
rect 352826 678218 353062 678454
rect 353146 678218 353382 678454
rect 352826 677898 353062 678134
rect 353146 677898 353382 678134
rect 352826 642218 353062 642454
rect 353146 642218 353382 642454
rect 352826 641898 353062 642134
rect 353146 641898 353382 642134
rect 352826 606218 353062 606454
rect 353146 606218 353382 606454
rect 352826 605898 353062 606134
rect 353146 605898 353382 606134
rect 352826 570218 353062 570454
rect 353146 570218 353382 570454
rect 352826 569898 353062 570134
rect 353146 569898 353382 570134
rect 352826 534218 353062 534454
rect 353146 534218 353382 534454
rect 352826 533898 353062 534134
rect 353146 533898 353382 534134
rect 352826 498218 353062 498454
rect 353146 498218 353382 498454
rect 352826 497898 353062 498134
rect 353146 497898 353382 498134
rect 352826 462218 353062 462454
rect 353146 462218 353382 462454
rect 352826 461898 353062 462134
rect 353146 461898 353382 462134
rect 352826 426218 353062 426454
rect 353146 426218 353382 426454
rect 352826 425898 353062 426134
rect 353146 425898 353382 426134
rect 352826 390218 353062 390454
rect 353146 390218 353382 390454
rect 352826 389898 353062 390134
rect 353146 389898 353382 390134
rect 352826 354218 353062 354454
rect 353146 354218 353382 354454
rect 352826 353898 353062 354134
rect 353146 353898 353382 354134
rect 352826 318218 353062 318454
rect 353146 318218 353382 318454
rect 352826 317898 353062 318134
rect 353146 317898 353382 318134
rect 352826 282218 353062 282454
rect 353146 282218 353382 282454
rect 352826 281898 353062 282134
rect 353146 281898 353382 282134
rect 357326 711322 357562 711558
rect 357646 711322 357882 711558
rect 357326 711002 357562 711238
rect 357646 711002 357882 711238
rect 357326 682718 357562 682954
rect 357646 682718 357882 682954
rect 357326 682398 357562 682634
rect 357646 682398 357882 682634
rect 357326 646718 357562 646954
rect 357646 646718 357882 646954
rect 357326 646398 357562 646634
rect 357646 646398 357882 646634
rect 357326 610718 357562 610954
rect 357646 610718 357882 610954
rect 357326 610398 357562 610634
rect 357646 610398 357882 610634
rect 357326 574718 357562 574954
rect 357646 574718 357882 574954
rect 357326 574398 357562 574634
rect 357646 574398 357882 574634
rect 357326 538718 357562 538954
rect 357646 538718 357882 538954
rect 357326 538398 357562 538634
rect 357646 538398 357882 538634
rect 357326 502718 357562 502954
rect 357646 502718 357882 502954
rect 357326 502398 357562 502634
rect 357646 502398 357882 502634
rect 357326 466718 357562 466954
rect 357646 466718 357882 466954
rect 357326 466398 357562 466634
rect 357646 466398 357882 466634
rect 357326 430718 357562 430954
rect 357646 430718 357882 430954
rect 357326 430398 357562 430634
rect 357646 430398 357882 430634
rect 357326 394718 357562 394954
rect 357646 394718 357882 394954
rect 357326 394398 357562 394634
rect 357646 394398 357882 394634
rect 357326 358718 357562 358954
rect 357646 358718 357882 358954
rect 357326 358398 357562 358634
rect 357646 358398 357882 358634
rect 357326 322718 357562 322954
rect 357646 322718 357882 322954
rect 357326 322398 357562 322634
rect 357646 322398 357882 322634
rect 357326 286718 357562 286954
rect 357646 286718 357882 286954
rect 357326 286398 357562 286634
rect 357646 286398 357882 286634
rect 357326 250718 357562 250954
rect 357646 250718 357882 250954
rect 357326 250398 357562 250634
rect 357646 250398 357882 250634
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 366326 705562 366562 705798
rect 366646 705562 366882 705798
rect 366326 705242 366562 705478
rect 366646 705242 366882 705478
rect 366326 691718 366562 691954
rect 366646 691718 366882 691954
rect 366326 691398 366562 691634
rect 366646 691398 366882 691634
rect 366326 655718 366562 655954
rect 366646 655718 366882 655954
rect 366326 655398 366562 655634
rect 366646 655398 366882 655634
rect 366326 619718 366562 619954
rect 366646 619718 366882 619954
rect 366326 619398 366562 619634
rect 366646 619398 366882 619634
rect 366326 583718 366562 583954
rect 366646 583718 366882 583954
rect 366326 583398 366562 583634
rect 366646 583398 366882 583634
rect 366326 547718 366562 547954
rect 366646 547718 366882 547954
rect 366326 547398 366562 547634
rect 366646 547398 366882 547634
rect 366326 511718 366562 511954
rect 366646 511718 366882 511954
rect 366326 511398 366562 511634
rect 366646 511398 366882 511634
rect 366326 475718 366562 475954
rect 366646 475718 366882 475954
rect 366326 475398 366562 475634
rect 366646 475398 366882 475634
rect 366326 439718 366562 439954
rect 366646 439718 366882 439954
rect 366326 439398 366562 439634
rect 366646 439398 366882 439634
rect 366326 403718 366562 403954
rect 366646 403718 366882 403954
rect 366326 403398 366562 403634
rect 366646 403398 366882 403634
rect 366326 367718 366562 367954
rect 366646 367718 366882 367954
rect 366326 367398 366562 367634
rect 366646 367398 366882 367634
rect 366326 331718 366562 331954
rect 366646 331718 366882 331954
rect 366326 331398 366562 331634
rect 366646 331398 366882 331634
rect 366326 295718 366562 295954
rect 366646 295718 366882 295954
rect 366326 295398 366562 295634
rect 366646 295398 366882 295634
rect 366326 259718 366562 259954
rect 366646 259718 366882 259954
rect 366326 259398 366562 259634
rect 366646 259398 366882 259634
rect 370826 706522 371062 706758
rect 371146 706522 371382 706758
rect 370826 706202 371062 706438
rect 371146 706202 371382 706438
rect 370826 696218 371062 696454
rect 371146 696218 371382 696454
rect 370826 695898 371062 696134
rect 371146 695898 371382 696134
rect 370826 660218 371062 660454
rect 371146 660218 371382 660454
rect 370826 659898 371062 660134
rect 371146 659898 371382 660134
rect 370826 624218 371062 624454
rect 371146 624218 371382 624454
rect 370826 623898 371062 624134
rect 371146 623898 371382 624134
rect 370826 588218 371062 588454
rect 371146 588218 371382 588454
rect 370826 587898 371062 588134
rect 371146 587898 371382 588134
rect 370826 552218 371062 552454
rect 371146 552218 371382 552454
rect 370826 551898 371062 552134
rect 371146 551898 371382 552134
rect 370826 516218 371062 516454
rect 371146 516218 371382 516454
rect 370826 515898 371062 516134
rect 371146 515898 371382 516134
rect 370826 480218 371062 480454
rect 371146 480218 371382 480454
rect 370826 479898 371062 480134
rect 371146 479898 371382 480134
rect 370826 444218 371062 444454
rect 371146 444218 371382 444454
rect 370826 443898 371062 444134
rect 371146 443898 371382 444134
rect 370826 408218 371062 408454
rect 371146 408218 371382 408454
rect 370826 407898 371062 408134
rect 371146 407898 371382 408134
rect 370826 372218 371062 372454
rect 371146 372218 371382 372454
rect 370826 371898 371062 372134
rect 371146 371898 371382 372134
rect 370826 336218 371062 336454
rect 371146 336218 371382 336454
rect 370826 335898 371062 336134
rect 371146 335898 371382 336134
rect 370826 300218 371062 300454
rect 371146 300218 371382 300454
rect 370826 299898 371062 300134
rect 371146 299898 371382 300134
rect 370826 264218 371062 264454
rect 371146 264218 371382 264454
rect 370826 263898 371062 264134
rect 371146 263898 371382 264134
rect 375326 707482 375562 707718
rect 375646 707482 375882 707718
rect 375326 707162 375562 707398
rect 375646 707162 375882 707398
rect 375326 700718 375562 700954
rect 375646 700718 375882 700954
rect 375326 700398 375562 700634
rect 375646 700398 375882 700634
rect 375326 664718 375562 664954
rect 375646 664718 375882 664954
rect 375326 664398 375562 664634
rect 375646 664398 375882 664634
rect 375326 628718 375562 628954
rect 375646 628718 375882 628954
rect 375326 628398 375562 628634
rect 375646 628398 375882 628634
rect 375326 592718 375562 592954
rect 375646 592718 375882 592954
rect 375326 592398 375562 592634
rect 375646 592398 375882 592634
rect 375326 556718 375562 556954
rect 375646 556718 375882 556954
rect 375326 556398 375562 556634
rect 375646 556398 375882 556634
rect 375326 520718 375562 520954
rect 375646 520718 375882 520954
rect 375326 520398 375562 520634
rect 375646 520398 375882 520634
rect 375326 484718 375562 484954
rect 375646 484718 375882 484954
rect 375326 484398 375562 484634
rect 375646 484398 375882 484634
rect 375326 448718 375562 448954
rect 375646 448718 375882 448954
rect 375326 448398 375562 448634
rect 375646 448398 375882 448634
rect 375326 412718 375562 412954
rect 375646 412718 375882 412954
rect 375326 412398 375562 412634
rect 375646 412398 375882 412634
rect 375326 376718 375562 376954
rect 375646 376718 375882 376954
rect 375326 376398 375562 376634
rect 375646 376398 375882 376634
rect 375326 340718 375562 340954
rect 375646 340718 375882 340954
rect 375326 340398 375562 340634
rect 375646 340398 375882 340634
rect 375326 304718 375562 304954
rect 375646 304718 375882 304954
rect 375326 304398 375562 304634
rect 375646 304398 375882 304634
rect 375326 268718 375562 268954
rect 375646 268718 375882 268954
rect 375326 268398 375562 268634
rect 375646 268398 375882 268634
rect 379826 708442 380062 708678
rect 380146 708442 380382 708678
rect 379826 708122 380062 708358
rect 380146 708122 380382 708358
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 384326 709402 384562 709638
rect 384646 709402 384882 709638
rect 384326 709082 384562 709318
rect 384646 709082 384882 709318
rect 384326 673718 384562 673954
rect 384646 673718 384882 673954
rect 384326 673398 384562 673634
rect 384646 673398 384882 673634
rect 384326 637718 384562 637954
rect 384646 637718 384882 637954
rect 384326 637398 384562 637634
rect 384646 637398 384882 637634
rect 384326 601718 384562 601954
rect 384646 601718 384882 601954
rect 384326 601398 384562 601634
rect 384646 601398 384882 601634
rect 384326 565718 384562 565954
rect 384646 565718 384882 565954
rect 384326 565398 384562 565634
rect 384646 565398 384882 565634
rect 384326 529718 384562 529954
rect 384646 529718 384882 529954
rect 384326 529398 384562 529634
rect 384646 529398 384882 529634
rect 384326 493718 384562 493954
rect 384646 493718 384882 493954
rect 384326 493398 384562 493634
rect 384646 493398 384882 493634
rect 384326 457718 384562 457954
rect 384646 457718 384882 457954
rect 384326 457398 384562 457634
rect 384646 457398 384882 457634
rect 384326 421718 384562 421954
rect 384646 421718 384882 421954
rect 384326 421398 384562 421634
rect 384646 421398 384882 421634
rect 384326 385718 384562 385954
rect 384646 385718 384882 385954
rect 384326 385398 384562 385634
rect 384646 385398 384882 385634
rect 384326 349718 384562 349954
rect 384646 349718 384882 349954
rect 384326 349398 384562 349634
rect 384646 349398 384882 349634
rect 384326 313718 384562 313954
rect 384646 313718 384882 313954
rect 384326 313398 384562 313634
rect 384646 313398 384882 313634
rect 384326 277718 384562 277954
rect 384646 277718 384882 277954
rect 384326 277398 384562 277634
rect 384646 277398 384882 277634
rect 388826 710362 389062 710598
rect 389146 710362 389382 710598
rect 388826 710042 389062 710278
rect 389146 710042 389382 710278
rect 388826 678218 389062 678454
rect 389146 678218 389382 678454
rect 388826 677898 389062 678134
rect 389146 677898 389382 678134
rect 388826 642218 389062 642454
rect 389146 642218 389382 642454
rect 388826 641898 389062 642134
rect 389146 641898 389382 642134
rect 388826 606218 389062 606454
rect 389146 606218 389382 606454
rect 388826 605898 389062 606134
rect 389146 605898 389382 606134
rect 388826 570218 389062 570454
rect 389146 570218 389382 570454
rect 388826 569898 389062 570134
rect 389146 569898 389382 570134
rect 388826 534218 389062 534454
rect 389146 534218 389382 534454
rect 388826 533898 389062 534134
rect 389146 533898 389382 534134
rect 388826 498218 389062 498454
rect 389146 498218 389382 498454
rect 388826 497898 389062 498134
rect 389146 497898 389382 498134
rect 388826 462218 389062 462454
rect 389146 462218 389382 462454
rect 388826 461898 389062 462134
rect 389146 461898 389382 462134
rect 388826 426218 389062 426454
rect 389146 426218 389382 426454
rect 388826 425898 389062 426134
rect 389146 425898 389382 426134
rect 388826 390218 389062 390454
rect 389146 390218 389382 390454
rect 388826 389898 389062 390134
rect 389146 389898 389382 390134
rect 388826 354218 389062 354454
rect 389146 354218 389382 354454
rect 388826 353898 389062 354134
rect 389146 353898 389382 354134
rect 388826 318218 389062 318454
rect 389146 318218 389382 318454
rect 388826 317898 389062 318134
rect 389146 317898 389382 318134
rect 388826 282218 389062 282454
rect 389146 282218 389382 282454
rect 388826 281898 389062 282134
rect 389146 281898 389382 282134
rect 393326 711322 393562 711558
rect 393646 711322 393882 711558
rect 393326 711002 393562 711238
rect 393646 711002 393882 711238
rect 393326 682718 393562 682954
rect 393646 682718 393882 682954
rect 393326 682398 393562 682634
rect 393646 682398 393882 682634
rect 393326 646718 393562 646954
rect 393646 646718 393882 646954
rect 393326 646398 393562 646634
rect 393646 646398 393882 646634
rect 393326 610718 393562 610954
rect 393646 610718 393882 610954
rect 393326 610398 393562 610634
rect 393646 610398 393882 610634
rect 393326 574718 393562 574954
rect 393646 574718 393882 574954
rect 393326 574398 393562 574634
rect 393646 574398 393882 574634
rect 393326 538718 393562 538954
rect 393646 538718 393882 538954
rect 393326 538398 393562 538634
rect 393646 538398 393882 538634
rect 393326 502718 393562 502954
rect 393646 502718 393882 502954
rect 393326 502398 393562 502634
rect 393646 502398 393882 502634
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 393326 466718 393562 466954
rect 393646 466718 393882 466954
rect 393326 466398 393562 466634
rect 393646 466398 393882 466634
rect 393326 430718 393562 430954
rect 393646 430718 393882 430954
rect 393326 430398 393562 430634
rect 393646 430398 393882 430634
rect 393326 394718 393562 394954
rect 393646 394718 393882 394954
rect 393326 394398 393562 394634
rect 393646 394398 393882 394634
rect 393326 358718 393562 358954
rect 393646 358718 393882 358954
rect 393326 358398 393562 358634
rect 393646 358398 393882 358634
rect 393326 322718 393562 322954
rect 393646 322718 393882 322954
rect 393326 322398 393562 322634
rect 393646 322398 393882 322634
rect 393326 286718 393562 286954
rect 393646 286718 393882 286954
rect 393326 286398 393562 286634
rect 393646 286398 393882 286634
rect 393326 250718 393562 250954
rect 393646 250718 393882 250954
rect 393326 250398 393562 250634
rect 393646 250398 393882 250634
rect 65342 246067 65578 246303
rect 65662 246067 65898 246303
rect 65982 246067 66218 246303
rect 66302 246067 66538 246303
rect 66622 246067 66858 246303
rect 66942 246067 67178 246303
rect 67262 246067 67498 246303
rect 67582 246067 67818 246303
rect 67902 246067 68138 246303
rect 68222 246067 68458 246303
rect 68542 246067 68778 246303
rect 68862 246067 69098 246303
rect 69182 246067 69418 246303
rect 69502 246067 69738 246303
rect 69822 246067 70058 246303
rect 65462 241717 65698 241953
rect 65782 241717 66018 241953
rect 66102 241717 66338 241953
rect 66422 241717 66658 241953
rect 66742 241717 66978 241953
rect 67062 241717 67298 241953
rect 67382 241717 67618 241953
rect 67702 241717 67938 241953
rect 68022 241717 68258 241953
rect 68342 241717 68578 241953
rect 68662 241717 68898 241953
rect 68982 241717 69218 241953
rect 69302 241717 69538 241953
rect 69622 241717 69858 241953
rect 69942 241717 70178 241953
rect 70262 241717 70498 241953
rect 70582 241717 70818 241953
rect 70902 241717 71138 241953
rect 65462 241397 65698 241633
rect 65782 241397 66018 241633
rect 66102 241397 66338 241633
rect 66422 241397 66658 241633
rect 66742 241397 66978 241633
rect 67062 241397 67298 241633
rect 67382 241397 67618 241633
rect 67702 241397 67938 241633
rect 68022 241397 68258 241633
rect 68342 241397 68578 241633
rect 68662 241397 68898 241633
rect 68982 241397 69218 241633
rect 69302 241397 69538 241633
rect 69622 241397 69858 241633
rect 69942 241397 70178 241633
rect 70262 241397 70498 241633
rect 70582 241397 70818 241633
rect 70902 241397 71138 241633
rect 42326 223718 42562 223954
rect 42646 223718 42882 223954
rect 42326 223398 42562 223634
rect 42646 223398 42882 223634
rect 42326 187718 42562 187954
rect 42646 187718 42882 187954
rect 42326 187398 42562 187634
rect 42646 187398 42882 187634
rect 42326 151718 42562 151954
rect 42646 151718 42882 151954
rect 42326 151398 42562 151634
rect 42646 151398 42882 151634
rect 42326 115718 42562 115954
rect 42646 115718 42882 115954
rect 42326 115398 42562 115634
rect 42646 115398 42882 115634
rect 42326 79718 42562 79954
rect 42646 79718 42882 79954
rect 42326 79398 42562 79634
rect 42646 79398 42882 79634
rect 42326 43718 42562 43954
rect 42646 43718 42882 43954
rect 42326 43398 42562 43634
rect 42646 43398 42882 43634
rect 42326 7718 42562 7954
rect 42646 7718 42882 7954
rect 42326 7398 42562 7634
rect 42646 7398 42882 7634
rect 42326 -1542 42562 -1306
rect 42646 -1542 42882 -1306
rect 42326 -1862 42562 -1626
rect 42646 -1862 42882 -1626
rect 46826 228217 47062 228453
rect 47146 228217 47382 228453
rect 46826 227897 47062 228133
rect 47146 227897 47382 228133
rect 46826 192218 47062 192454
rect 47146 192218 47382 192454
rect 46826 191898 47062 192134
rect 47146 191898 47382 192134
rect 46826 156218 47062 156454
rect 47146 156218 47382 156454
rect 46826 155898 47062 156134
rect 47146 155898 47382 156134
rect 46826 120218 47062 120454
rect 47146 120218 47382 120454
rect 46826 119898 47062 120134
rect 47146 119898 47382 120134
rect 46826 84218 47062 84454
rect 47146 84218 47382 84454
rect 46826 83898 47062 84134
rect 47146 83898 47382 84134
rect 46826 48218 47062 48454
rect 47146 48218 47382 48454
rect 46826 47898 47062 48134
rect 47146 47898 47382 48134
rect 46826 12218 47062 12454
rect 47146 12218 47382 12454
rect 46826 11898 47062 12134
rect 47146 11898 47382 12134
rect 46826 -2502 47062 -2266
rect 47146 -2502 47382 -2266
rect 46826 -2822 47062 -2586
rect 47146 -2822 47382 -2586
rect 51326 196718 51562 196954
rect 51646 196718 51882 196954
rect 51326 196398 51562 196634
rect 51646 196398 51882 196634
rect 51326 160718 51562 160954
rect 51646 160718 51882 160954
rect 51326 160398 51562 160634
rect 51646 160398 51882 160634
rect 51326 124718 51562 124954
rect 51646 124718 51882 124954
rect 51326 124398 51562 124634
rect 51646 124398 51882 124634
rect 51326 88718 51562 88954
rect 51646 88718 51882 88954
rect 51326 88398 51562 88634
rect 51646 88398 51882 88634
rect 51326 52718 51562 52954
rect 51646 52718 51882 52954
rect 51326 52398 51562 52634
rect 51646 52398 51882 52634
rect 51326 16718 51562 16954
rect 51646 16718 51882 16954
rect 51326 16398 51562 16634
rect 51646 16398 51882 16634
rect 51326 -3462 51562 -3226
rect 51646 -3462 51882 -3226
rect 51326 -3782 51562 -3546
rect 51646 -3782 51882 -3546
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -4422 56062 -4186
rect 56146 -4422 56382 -4186
rect 55826 -4742 56062 -4506
rect 56146 -4742 56382 -4506
rect 60326 205718 60562 205954
rect 60646 205718 60882 205954
rect 60326 205398 60562 205634
rect 60646 205398 60882 205634
rect 60326 169718 60562 169954
rect 60646 169718 60882 169954
rect 60326 169398 60562 169634
rect 60646 169398 60882 169634
rect 60326 133718 60562 133954
rect 60646 133718 60882 133954
rect 60326 133398 60562 133634
rect 60646 133398 60882 133634
rect 60326 97718 60562 97954
rect 60646 97718 60882 97954
rect 60326 97398 60562 97634
rect 60646 97398 60882 97634
rect 60326 61718 60562 61954
rect 60646 61718 60882 61954
rect 60326 61398 60562 61634
rect 60646 61398 60882 61634
rect 60326 25718 60562 25954
rect 60646 25718 60882 25954
rect 60326 25398 60562 25634
rect 60646 25398 60882 25634
rect 60326 -5382 60562 -5146
rect 60646 -5382 60882 -5146
rect 60326 -5702 60562 -5466
rect 60646 -5702 60882 -5466
rect 64826 210218 65062 210454
rect 65146 210218 65382 210454
rect 64826 209898 65062 210134
rect 65146 209898 65382 210134
rect 64826 174218 65062 174454
rect 65146 174218 65382 174454
rect 64826 173898 65062 174134
rect 65146 173898 65382 174134
rect 64826 138218 65062 138454
rect 65146 138218 65382 138454
rect 64826 137898 65062 138134
rect 65146 137898 65382 138134
rect 64826 102218 65062 102454
rect 65146 102218 65382 102454
rect 64826 101898 65062 102134
rect 65146 101898 65382 102134
rect 64826 66218 65062 66454
rect 65146 66218 65382 66454
rect 64826 65898 65062 66134
rect 65146 65898 65382 66134
rect 64826 30218 65062 30454
rect 65146 30218 65382 30454
rect 64826 29898 65062 30134
rect 65146 29898 65382 30134
rect 64826 -6342 65062 -6106
rect 65146 -6342 65382 -6106
rect 64826 -6662 65062 -6426
rect 65146 -6662 65382 -6426
rect 69326 214718 69562 214954
rect 69646 214718 69882 214954
rect 69326 214398 69562 214634
rect 69646 214398 69882 214634
rect 69326 178718 69562 178954
rect 69646 178718 69882 178954
rect 69326 178398 69562 178634
rect 69646 178398 69882 178634
rect 69326 142718 69562 142954
rect 69646 142718 69882 142954
rect 69326 142398 69562 142634
rect 69646 142398 69882 142634
rect 69326 106718 69562 106954
rect 69646 106718 69882 106954
rect 69326 106398 69562 106634
rect 69646 106398 69882 106634
rect 69326 70718 69562 70954
rect 69646 70718 69882 70954
rect 69326 70398 69562 70634
rect 69646 70398 69882 70634
rect 69326 34718 69562 34954
rect 69646 34718 69882 34954
rect 69326 34398 69562 34634
rect 69646 34398 69882 34634
rect 69326 -7302 69562 -7066
rect 69646 -7302 69882 -7066
rect 69326 -7622 69562 -7386
rect 69646 -7622 69882 -7386
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 78326 223718 78562 223954
rect 78646 223718 78882 223954
rect 78326 223398 78562 223634
rect 78646 223398 78882 223634
rect 78326 187718 78562 187954
rect 78646 187718 78882 187954
rect 78326 187398 78562 187634
rect 78646 187398 78882 187634
rect 78326 151718 78562 151954
rect 78646 151718 78882 151954
rect 78326 151398 78562 151634
rect 78646 151398 78882 151634
rect 78326 115718 78562 115954
rect 78646 115718 78882 115954
rect 78326 115398 78562 115634
rect 78646 115398 78882 115634
rect 78326 79718 78562 79954
rect 78646 79718 78882 79954
rect 78326 79398 78562 79634
rect 78646 79398 78882 79634
rect 78326 43718 78562 43954
rect 78646 43718 78882 43954
rect 78326 43398 78562 43634
rect 78646 43398 78882 43634
rect 78326 7718 78562 7954
rect 78646 7718 78882 7954
rect 78326 7398 78562 7634
rect 78646 7398 78882 7634
rect 78326 -1542 78562 -1306
rect 78646 -1542 78882 -1306
rect 78326 -1862 78562 -1626
rect 78646 -1862 78882 -1626
rect 82826 228217 83062 228453
rect 83146 228217 83382 228453
rect 82826 227897 83062 228133
rect 83146 227897 83382 228133
rect 82826 192218 83062 192454
rect 83146 192218 83382 192454
rect 82826 191898 83062 192134
rect 83146 191898 83382 192134
rect 82826 156218 83062 156454
rect 83146 156218 83382 156454
rect 82826 155898 83062 156134
rect 83146 155898 83382 156134
rect 82826 120218 83062 120454
rect 83146 120218 83382 120454
rect 82826 119898 83062 120134
rect 83146 119898 83382 120134
rect 82826 84218 83062 84454
rect 83146 84218 83382 84454
rect 82826 83898 83062 84134
rect 83146 83898 83382 84134
rect 82826 48218 83062 48454
rect 83146 48218 83382 48454
rect 82826 47898 83062 48134
rect 83146 47898 83382 48134
rect 82826 12218 83062 12454
rect 83146 12218 83382 12454
rect 82826 11898 83062 12134
rect 83146 11898 83382 12134
rect 82826 -2502 83062 -2266
rect 83146 -2502 83382 -2266
rect 82826 -2822 83062 -2586
rect 83146 -2822 83382 -2586
rect 87326 196718 87562 196954
rect 87646 196718 87882 196954
rect 87326 196398 87562 196634
rect 87646 196398 87882 196634
rect 87326 160718 87562 160954
rect 87646 160718 87882 160954
rect 87326 160398 87562 160634
rect 87646 160398 87882 160634
rect 87326 124718 87562 124954
rect 87646 124718 87882 124954
rect 87326 124398 87562 124634
rect 87646 124398 87882 124634
rect 87326 88718 87562 88954
rect 87646 88718 87882 88954
rect 87326 88398 87562 88634
rect 87646 88398 87882 88634
rect 87326 52718 87562 52954
rect 87646 52718 87882 52954
rect 87326 52398 87562 52634
rect 87646 52398 87882 52634
rect 87326 16718 87562 16954
rect 87646 16718 87882 16954
rect 87326 16398 87562 16634
rect 87646 16398 87882 16634
rect 87326 -3462 87562 -3226
rect 87646 -3462 87882 -3226
rect 87326 -3782 87562 -3546
rect 87646 -3782 87882 -3546
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 91826 129218 92062 129454
rect 92146 129218 92382 129454
rect 91826 128898 92062 129134
rect 92146 128898 92382 129134
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -4422 92062 -4186
rect 92146 -4422 92382 -4186
rect 91826 -4742 92062 -4506
rect 92146 -4742 92382 -4506
rect 96326 205718 96562 205954
rect 96646 205718 96882 205954
rect 96326 205398 96562 205634
rect 96646 205398 96882 205634
rect 96326 169718 96562 169954
rect 96646 169718 96882 169954
rect 96326 169398 96562 169634
rect 96646 169398 96882 169634
rect 96326 133718 96562 133954
rect 96646 133718 96882 133954
rect 96326 133398 96562 133634
rect 96646 133398 96882 133634
rect 96326 97718 96562 97954
rect 96646 97718 96882 97954
rect 96326 97398 96562 97634
rect 96646 97398 96882 97634
rect 96326 61718 96562 61954
rect 96646 61718 96882 61954
rect 96326 61398 96562 61634
rect 96646 61398 96882 61634
rect 96326 25718 96562 25954
rect 96646 25718 96882 25954
rect 96326 25398 96562 25634
rect 96646 25398 96882 25634
rect 96326 -5382 96562 -5146
rect 96646 -5382 96882 -5146
rect 96326 -5702 96562 -5466
rect 96646 -5702 96882 -5466
rect 100826 210218 101062 210454
rect 101146 210218 101382 210454
rect 100826 209898 101062 210134
rect 101146 209898 101382 210134
rect 100826 174218 101062 174454
rect 101146 174218 101382 174454
rect 100826 173898 101062 174134
rect 101146 173898 101382 174134
rect 100826 138218 101062 138454
rect 101146 138218 101382 138454
rect 100826 137898 101062 138134
rect 101146 137898 101382 138134
rect 100826 102218 101062 102454
rect 101146 102218 101382 102454
rect 100826 101898 101062 102134
rect 101146 101898 101382 102134
rect 100826 66218 101062 66454
rect 101146 66218 101382 66454
rect 100826 65898 101062 66134
rect 101146 65898 101382 66134
rect 100826 30218 101062 30454
rect 101146 30218 101382 30454
rect 100826 29898 101062 30134
rect 101146 29898 101382 30134
rect 100826 -6342 101062 -6106
rect 101146 -6342 101382 -6106
rect 100826 -6662 101062 -6426
rect 101146 -6662 101382 -6426
rect 105326 214718 105562 214954
rect 105646 214718 105882 214954
rect 105326 214398 105562 214634
rect 105646 214398 105882 214634
rect 105326 178718 105562 178954
rect 105646 178718 105882 178954
rect 105326 178398 105562 178634
rect 105646 178398 105882 178634
rect 105326 142718 105562 142954
rect 105646 142718 105882 142954
rect 105326 142398 105562 142634
rect 105646 142398 105882 142634
rect 105326 106718 105562 106954
rect 105646 106718 105882 106954
rect 105326 106398 105562 106634
rect 105646 106398 105882 106634
rect 105326 70718 105562 70954
rect 105646 70718 105882 70954
rect 105326 70398 105562 70634
rect 105646 70398 105882 70634
rect 105326 34718 105562 34954
rect 105646 34718 105882 34954
rect 105326 34398 105562 34634
rect 105646 34398 105882 34634
rect 105326 -7302 105562 -7066
rect 105646 -7302 105882 -7066
rect 105326 -7622 105562 -7386
rect 105646 -7622 105882 -7386
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 114326 223718 114562 223954
rect 114646 223718 114882 223954
rect 114326 223398 114562 223634
rect 114646 223398 114882 223634
rect 114326 187718 114562 187954
rect 114646 187718 114882 187954
rect 114326 187398 114562 187634
rect 114646 187398 114882 187634
rect 114326 151718 114562 151954
rect 114646 151718 114882 151954
rect 114326 151398 114562 151634
rect 114646 151398 114882 151634
rect 118826 228217 119062 228453
rect 119146 228217 119382 228453
rect 118826 227897 119062 228133
rect 119146 227897 119382 228133
rect 118826 192218 119062 192454
rect 119146 192218 119382 192454
rect 118826 191898 119062 192134
rect 119146 191898 119382 192134
rect 118826 156218 119062 156454
rect 119146 156218 119382 156454
rect 118826 155898 119062 156134
rect 119146 155898 119382 156134
rect 123326 196718 123562 196954
rect 123646 196718 123882 196954
rect 123326 196398 123562 196634
rect 123646 196398 123882 196634
rect 123326 160718 123562 160954
rect 123646 160718 123882 160954
rect 123326 160398 123562 160634
rect 123646 160398 123882 160634
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 127826 165218 128062 165454
rect 128146 165218 128382 165454
rect 127826 164898 128062 165134
rect 128146 164898 128382 165134
rect 172826 210218 173062 210454
rect 173146 210218 173382 210454
rect 172826 209898 173062 210134
rect 173146 209898 173382 210134
rect 132326 205718 132562 205954
rect 132646 205718 132882 205954
rect 132326 205398 132562 205634
rect 132646 205398 132882 205634
rect 136036 205625 136272 205861
rect 136356 205625 136592 205861
rect 136676 205625 136912 205861
rect 136996 205625 137232 205861
rect 137316 205625 137552 205861
rect 137636 205625 137872 205861
rect 137956 205625 138192 205861
rect 138276 205625 138512 205861
rect 138596 205625 138832 205861
rect 138916 205625 139152 205861
rect 139236 205625 139472 205861
rect 139556 205625 139792 205861
rect 139876 205625 140112 205861
rect 140196 205625 140432 205861
rect 140516 205625 140752 205861
rect 140836 205625 141072 205861
rect 141156 205625 141392 205861
rect 141476 205625 141712 205861
rect 141796 205625 142032 205861
rect 142116 205625 142352 205861
rect 142436 205625 142672 205861
rect 142756 205625 142992 205861
rect 143076 205625 143312 205861
rect 143396 205625 143632 205861
rect 143716 205625 143952 205861
rect 144036 205625 144272 205861
rect 144356 205625 144592 205861
rect 144676 205625 144912 205861
rect 144996 205625 145232 205861
rect 145316 205625 145552 205861
rect 145636 205625 145872 205861
rect 145956 205625 146192 205861
rect 146276 205625 146512 205861
rect 146596 205625 146832 205861
rect 146916 205625 147152 205861
rect 147236 205625 147472 205861
rect 147556 205625 147792 205861
rect 147876 205625 148112 205861
rect 148196 205625 148432 205861
rect 148516 205625 148752 205861
rect 148836 205625 149072 205861
rect 149156 205625 149392 205861
rect 149476 205625 149712 205861
rect 149796 205625 150032 205861
rect 150116 205625 150352 205861
rect 150436 205625 150672 205861
rect 150756 205625 150992 205861
rect 151076 205625 151312 205861
rect 151396 205625 151632 205861
rect 151716 205625 151952 205861
rect 152036 205625 152272 205861
rect 152356 205625 152592 205861
rect 152676 205625 152912 205861
rect 152996 205625 153232 205861
rect 153316 205625 153552 205861
rect 153636 205625 153872 205861
rect 153956 205625 154192 205861
rect 154276 205625 154512 205861
rect 154596 205625 154832 205861
rect 154916 205625 155152 205861
rect 155236 205625 155472 205861
rect 155556 205625 155792 205861
rect 155876 205625 156112 205861
rect 156196 205625 156432 205861
rect 156516 205625 156752 205861
rect 156836 205625 157072 205861
rect 157156 205625 157392 205861
rect 157476 205625 157712 205861
rect 157796 205625 158032 205861
rect 158116 205625 158352 205861
rect 158436 205625 158672 205861
rect 158756 205625 158992 205861
rect 159076 205625 159312 205861
rect 159396 205625 159632 205861
rect 159716 205625 159952 205861
rect 160036 205625 160272 205861
rect 160356 205625 160592 205861
rect 160676 205625 160912 205861
rect 160996 205625 161232 205861
rect 161316 205625 161552 205861
rect 161636 205625 161872 205861
rect 161956 205625 162192 205861
rect 162276 205625 162512 205861
rect 162596 205625 162832 205861
rect 162916 205625 163152 205861
rect 163236 205625 163472 205861
rect 163556 205625 163792 205861
rect 163876 205625 164112 205861
rect 164196 205625 164432 205861
rect 164516 205625 164752 205861
rect 164836 205625 165072 205861
rect 165156 205625 165392 205861
rect 137376 201175 137612 201411
rect 137696 201175 137932 201411
rect 138016 201175 138252 201411
rect 138336 201175 138572 201411
rect 138656 201175 138892 201411
rect 138976 201175 139212 201411
rect 139296 201175 139532 201411
rect 139616 201175 139852 201411
rect 139936 201175 140172 201411
rect 140256 201175 140492 201411
rect 140576 201175 140812 201411
rect 140896 201175 141132 201411
rect 141216 201175 141452 201411
rect 141536 201175 141772 201411
rect 141856 201175 142092 201411
rect 142176 201175 142412 201411
rect 142496 201175 142732 201411
rect 142816 201175 143052 201411
rect 143136 201175 143372 201411
rect 143456 201175 143692 201411
rect 143776 201175 144012 201411
rect 144096 201175 144332 201411
rect 144416 201175 144652 201411
rect 144736 201175 144972 201411
rect 145056 201175 145292 201411
rect 145376 201175 145612 201411
rect 145696 201175 145932 201411
rect 146016 201175 146252 201411
rect 146336 201175 146572 201411
rect 146656 201175 146892 201411
rect 146976 201175 147212 201411
rect 147296 201175 147532 201411
rect 147616 201175 147852 201411
rect 147936 201175 148172 201411
rect 148256 201175 148492 201411
rect 148576 201175 148812 201411
rect 148896 201175 149132 201411
rect 149216 201175 149452 201411
rect 149536 201175 149772 201411
rect 149856 201175 150092 201411
rect 150176 201175 150412 201411
rect 150496 201175 150732 201411
rect 150816 201175 151052 201411
rect 151136 201175 151372 201411
rect 151456 201175 151692 201411
rect 151776 201175 152012 201411
rect 152096 201175 152332 201411
rect 152416 201175 152652 201411
rect 152736 201175 152972 201411
rect 153056 201175 153292 201411
rect 153376 201175 153612 201411
rect 153696 201175 153932 201411
rect 154016 201175 154252 201411
rect 154336 201175 154572 201411
rect 154656 201175 154892 201411
rect 154976 201175 155212 201411
rect 155296 201175 155532 201411
rect 155616 201175 155852 201411
rect 155936 201175 156172 201411
rect 156256 201175 156492 201411
rect 156576 201175 156812 201411
rect 156896 201175 157132 201411
rect 157216 201175 157452 201411
rect 157536 201175 157772 201411
rect 157856 201175 158092 201411
rect 158176 201175 158412 201411
rect 158496 201175 158732 201411
rect 158816 201175 159052 201411
rect 159136 201175 159372 201411
rect 159456 201175 159692 201411
rect 159776 201175 160012 201411
rect 160096 201175 160332 201411
rect 160416 201175 160652 201411
rect 160736 201175 160972 201411
rect 161056 201175 161292 201411
rect 161376 201175 161612 201411
rect 161696 201175 161932 201411
rect 162016 201175 162252 201411
rect 162336 201175 162572 201411
rect 162656 201175 162892 201411
rect 162976 201175 163212 201411
rect 163296 201175 163532 201411
rect 163616 201175 163852 201411
rect 163936 201175 164172 201411
rect 164256 201175 164492 201411
rect 164576 201175 164812 201411
rect 164896 201175 165132 201411
rect 165216 201175 165452 201411
rect 137066 174218 137302 174454
rect 137386 174218 137622 174454
rect 137706 174218 137942 174454
rect 138026 174218 138262 174454
rect 138346 174218 138582 174454
rect 138666 174218 138902 174454
rect 138986 174218 139222 174454
rect 139306 174218 139542 174454
rect 139626 174218 139862 174454
rect 139946 174218 140182 174454
rect 140266 174218 140502 174454
rect 140586 174218 140822 174454
rect 140906 174218 141142 174454
rect 141226 174218 141462 174454
rect 137066 173898 137302 174134
rect 137386 173898 137622 174134
rect 137706 173898 137942 174134
rect 138026 173898 138262 174134
rect 138346 173898 138582 174134
rect 138666 173898 138902 174134
rect 138986 173898 139222 174134
rect 139306 173898 139542 174134
rect 139626 173898 139862 174134
rect 139946 173898 140182 174134
rect 140266 173898 140502 174134
rect 140586 173898 140822 174134
rect 140906 173898 141142 174134
rect 141226 173898 141462 174134
rect 132326 169718 132562 169954
rect 132646 169718 132882 169954
rect 132326 169398 132562 169634
rect 132646 169398 132882 169634
rect 172826 174218 173062 174454
rect 173146 174218 173382 174454
rect 172826 173898 173062 174134
rect 173146 173898 173382 174134
rect 172826 138218 173062 138454
rect 173146 138218 173382 138454
rect 172826 137898 173062 138134
rect 173146 137898 173382 138134
rect 177326 214718 177562 214954
rect 177646 214718 177882 214954
rect 177326 214398 177562 214634
rect 177646 214398 177882 214634
rect 177326 178718 177562 178954
rect 177646 178718 177882 178954
rect 177326 178398 177562 178634
rect 177646 178398 177882 178634
rect 177326 142718 177562 142954
rect 177646 142718 177882 142954
rect 177326 142398 177562 142634
rect 177646 142398 177882 142634
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 135610 115718 135846 115954
rect 135610 115398 135846 115634
rect 166330 115718 166566 115954
rect 166330 115398 166566 115634
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 120250 111218 120486 111454
rect 120250 110898 120486 111134
rect 150970 111218 151206 111454
rect 150970 110898 151206 111134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 135610 79718 135846 79954
rect 135610 79398 135846 79634
rect 166330 79718 166566 79954
rect 166330 79398 166566 79634
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 114326 43718 114562 43954
rect 114646 43718 114882 43954
rect 114326 43398 114562 43634
rect 114646 43398 114882 43634
rect 114326 7718 114562 7954
rect 114646 7718 114882 7954
rect 114326 7398 114562 7634
rect 114646 7398 114882 7634
rect 114326 -1542 114562 -1306
rect 114646 -1542 114882 -1306
rect 114326 -1862 114562 -1626
rect 114646 -1862 114882 -1626
rect 118826 48218 119062 48454
rect 119146 48218 119382 48454
rect 118826 47898 119062 48134
rect 119146 47898 119382 48134
rect 118826 12218 119062 12454
rect 119146 12218 119382 12454
rect 118826 11898 119062 12134
rect 119146 11898 119382 12134
rect 123326 52718 123562 52954
rect 123646 52718 123882 52954
rect 123326 52398 123562 52634
rect 123646 52398 123882 52634
rect 123326 16718 123562 16954
rect 123646 16718 123882 16954
rect 123326 16398 123562 16634
rect 123646 16398 123882 16634
rect 118826 -2502 119062 -2266
rect 119146 -2502 119382 -2266
rect 118826 -2822 119062 -2586
rect 119146 -2822 119382 -2586
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 123326 -3462 123562 -3226
rect 123646 -3462 123882 -3226
rect 123326 -3782 123562 -3546
rect 123646 -3782 123882 -3546
rect 132326 61718 132562 61954
rect 132646 61718 132882 61954
rect 132326 61398 132562 61634
rect 132646 61398 132882 61634
rect 132326 25718 132562 25954
rect 132646 25718 132882 25954
rect 132326 25398 132562 25634
rect 132646 25398 132882 25634
rect 127826 -4422 128062 -4186
rect 128146 -4422 128382 -4186
rect 127826 -4742 128062 -4506
rect 128146 -4742 128382 -4506
rect 136826 66218 137062 66454
rect 137146 66218 137382 66454
rect 136826 65898 137062 66134
rect 137146 65898 137382 66134
rect 136826 30218 137062 30454
rect 137146 30218 137382 30454
rect 136826 29898 137062 30134
rect 137146 29898 137382 30134
rect 132326 -5382 132562 -5146
rect 132646 -5382 132882 -5146
rect 132326 -5702 132562 -5466
rect 132646 -5702 132882 -5466
rect 141326 70718 141562 70954
rect 141646 70718 141882 70954
rect 141326 70398 141562 70634
rect 141646 70398 141882 70634
rect 141326 34718 141562 34954
rect 141646 34718 141882 34954
rect 141326 34398 141562 34634
rect 141646 34398 141882 34634
rect 136826 -6342 137062 -6106
rect 137146 -6342 137382 -6106
rect 136826 -6662 137062 -6426
rect 137146 -6662 137382 -6426
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 141326 -7302 141562 -7066
rect 141646 -7302 141882 -7066
rect 141326 -7622 141562 -7386
rect 141646 -7622 141882 -7386
rect 150326 43718 150562 43954
rect 150646 43718 150882 43954
rect 150326 43398 150562 43634
rect 150646 43398 150882 43634
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 150326 7718 150562 7954
rect 150646 7718 150882 7954
rect 150326 7398 150562 7634
rect 150646 7398 150882 7634
rect 154826 48218 155062 48454
rect 155146 48218 155382 48454
rect 154826 47898 155062 48134
rect 155146 47898 155382 48134
rect 154826 12218 155062 12454
rect 155146 12218 155382 12454
rect 154826 11898 155062 12134
rect 155146 11898 155382 12134
rect 150326 -1542 150562 -1306
rect 150646 -1542 150882 -1306
rect 150326 -1862 150562 -1626
rect 150646 -1862 150882 -1626
rect 159326 52718 159562 52954
rect 159646 52718 159882 52954
rect 159326 52398 159562 52634
rect 159646 52398 159882 52634
rect 159326 16718 159562 16954
rect 159646 16718 159882 16954
rect 159326 16398 159562 16634
rect 159646 16398 159882 16634
rect 154826 -2502 155062 -2266
rect 155146 -2502 155382 -2266
rect 154826 -2822 155062 -2586
rect 155146 -2822 155382 -2586
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 159326 -3462 159562 -3226
rect 159646 -3462 159882 -3226
rect 159326 -3782 159562 -3546
rect 159646 -3782 159882 -3546
rect 168326 61718 168562 61954
rect 168646 61718 168882 61954
rect 168326 61398 168562 61634
rect 168646 61398 168882 61634
rect 168326 25718 168562 25954
rect 168646 25718 168882 25954
rect 168326 25398 168562 25634
rect 168646 25398 168882 25634
rect 163826 -4422 164062 -4186
rect 164146 -4422 164382 -4186
rect 163826 -4742 164062 -4506
rect 164146 -4742 164382 -4506
rect 168326 -5382 168562 -5146
rect 168646 -5382 168882 -5146
rect 168326 -5702 168562 -5466
rect 168646 -5702 168882 -5466
rect 172826 66218 173062 66454
rect 173146 66218 173382 66454
rect 172826 65898 173062 66134
rect 173146 65898 173382 66134
rect 172826 30218 173062 30454
rect 173146 30218 173382 30454
rect 172826 29898 173062 30134
rect 173146 29898 173382 30134
rect 172826 -6342 173062 -6106
rect 173146 -6342 173382 -6106
rect 172826 -6662 173062 -6426
rect 173146 -6662 173382 -6426
rect 177326 70718 177562 70954
rect 177646 70718 177882 70954
rect 177326 70398 177562 70634
rect 177646 70398 177882 70634
rect 177326 34718 177562 34954
rect 177646 34718 177882 34954
rect 177326 34398 177562 34634
rect 177646 34398 177882 34634
rect 177326 -7302 177562 -7066
rect 177646 -7302 177882 -7066
rect 177326 -7622 177562 -7386
rect 177646 -7622 177882 -7386
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 186326 223718 186562 223954
rect 186646 223718 186882 223954
rect 186326 223398 186562 223634
rect 186646 223398 186882 223634
rect 186326 187718 186562 187954
rect 186646 187718 186882 187954
rect 186326 187398 186562 187634
rect 186646 187398 186882 187634
rect 186326 151718 186562 151954
rect 186646 151718 186882 151954
rect 186326 151398 186562 151634
rect 186646 151398 186882 151634
rect 186326 115718 186562 115954
rect 186646 115718 186882 115954
rect 186326 115398 186562 115634
rect 186646 115398 186882 115634
rect 186326 79718 186562 79954
rect 186646 79718 186882 79954
rect 186326 79398 186562 79634
rect 186646 79398 186882 79634
rect 186326 43718 186562 43954
rect 186646 43718 186882 43954
rect 186326 43398 186562 43634
rect 186646 43398 186882 43634
rect 186326 7718 186562 7954
rect 186646 7718 186882 7954
rect 186326 7398 186562 7634
rect 186646 7398 186882 7634
rect 186326 -1542 186562 -1306
rect 186646 -1542 186882 -1306
rect 186326 -1862 186562 -1626
rect 186646 -1862 186882 -1626
rect 190826 228217 191062 228453
rect 191146 228217 191382 228453
rect 190826 227897 191062 228133
rect 191146 227897 191382 228133
rect 190826 192218 191062 192454
rect 191146 192218 191382 192454
rect 190826 191898 191062 192134
rect 191146 191898 191382 192134
rect 190826 156218 191062 156454
rect 191146 156218 191382 156454
rect 190826 155898 191062 156134
rect 191146 155898 191382 156134
rect 190826 120218 191062 120454
rect 191146 120218 191382 120454
rect 190826 119898 191062 120134
rect 191146 119898 191382 120134
rect 190826 84218 191062 84454
rect 191146 84218 191382 84454
rect 190826 83898 191062 84134
rect 191146 83898 191382 84134
rect 190826 48218 191062 48454
rect 191146 48218 191382 48454
rect 190826 47898 191062 48134
rect 191146 47898 191382 48134
rect 190826 12218 191062 12454
rect 191146 12218 191382 12454
rect 190826 11898 191062 12134
rect 191146 11898 191382 12134
rect 190826 -2502 191062 -2266
rect 191146 -2502 191382 -2266
rect 190826 -2822 191062 -2586
rect 191146 -2822 191382 -2586
rect 195326 196718 195562 196954
rect 195646 196718 195882 196954
rect 195326 196398 195562 196634
rect 195646 196398 195882 196634
rect 195326 160718 195562 160954
rect 195646 160718 195882 160954
rect 195326 160398 195562 160634
rect 195646 160398 195882 160634
rect 195326 124718 195562 124954
rect 195646 124718 195882 124954
rect 195326 124398 195562 124634
rect 195646 124398 195882 124634
rect 195326 88718 195562 88954
rect 195646 88718 195882 88954
rect 195326 88398 195562 88634
rect 195646 88398 195882 88634
rect 195326 52718 195562 52954
rect 195646 52718 195882 52954
rect 195326 52398 195562 52634
rect 195646 52398 195882 52634
rect 195326 16718 195562 16954
rect 195646 16718 195882 16954
rect 195326 16398 195562 16634
rect 195646 16398 195882 16634
rect 195326 -3462 195562 -3226
rect 195646 -3462 195882 -3226
rect 195326 -3782 195562 -3546
rect 195646 -3782 195882 -3546
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -4422 200062 -4186
rect 200146 -4422 200382 -4186
rect 199826 -4742 200062 -4506
rect 200146 -4742 200382 -4506
rect 204326 205718 204562 205954
rect 204646 205718 204882 205954
rect 204326 205398 204562 205634
rect 204646 205398 204882 205634
rect 204326 169718 204562 169954
rect 204646 169718 204882 169954
rect 204326 169398 204562 169634
rect 204646 169398 204882 169634
rect 204326 133718 204562 133954
rect 204646 133718 204882 133954
rect 204326 133398 204562 133634
rect 204646 133398 204882 133634
rect 204326 97718 204562 97954
rect 204646 97718 204882 97954
rect 204326 97398 204562 97634
rect 204646 97398 204882 97634
rect 204326 61718 204562 61954
rect 204646 61718 204882 61954
rect 204326 61398 204562 61634
rect 204646 61398 204882 61634
rect 204326 25718 204562 25954
rect 204646 25718 204882 25954
rect 204326 25398 204562 25634
rect 204646 25398 204882 25634
rect 204326 -5382 204562 -5146
rect 204646 -5382 204882 -5146
rect 204326 -5702 204562 -5466
rect 204646 -5702 204882 -5466
rect 208826 210218 209062 210454
rect 209146 210218 209382 210454
rect 208826 209898 209062 210134
rect 209146 209898 209382 210134
rect 208826 174218 209062 174454
rect 209146 174218 209382 174454
rect 208826 173898 209062 174134
rect 209146 173898 209382 174134
rect 208826 138218 209062 138454
rect 209146 138218 209382 138454
rect 208826 137898 209062 138134
rect 209146 137898 209382 138134
rect 208826 102218 209062 102454
rect 209146 102218 209382 102454
rect 208826 101898 209062 102134
rect 209146 101898 209382 102134
rect 208826 66218 209062 66454
rect 209146 66218 209382 66454
rect 208826 65898 209062 66134
rect 209146 65898 209382 66134
rect 208826 30218 209062 30454
rect 209146 30218 209382 30454
rect 208826 29898 209062 30134
rect 209146 29898 209382 30134
rect 208826 -6342 209062 -6106
rect 209146 -6342 209382 -6106
rect 208826 -6662 209062 -6426
rect 209146 -6662 209382 -6426
rect 213326 214718 213562 214954
rect 213646 214718 213882 214954
rect 213326 214398 213562 214634
rect 213646 214398 213882 214634
rect 213326 178718 213562 178954
rect 213646 178718 213882 178954
rect 213326 178398 213562 178634
rect 213646 178398 213882 178634
rect 213326 142718 213562 142954
rect 213646 142718 213882 142954
rect 213326 142398 213562 142634
rect 213646 142398 213882 142634
rect 213326 106718 213562 106954
rect 213646 106718 213882 106954
rect 213326 106398 213562 106634
rect 213646 106398 213882 106634
rect 213326 70718 213562 70954
rect 213646 70718 213882 70954
rect 213326 70398 213562 70634
rect 213646 70398 213882 70634
rect 213326 34718 213562 34954
rect 213646 34718 213882 34954
rect 213326 34398 213562 34634
rect 213646 34398 213882 34634
rect 213326 -7302 213562 -7066
rect 213646 -7302 213882 -7066
rect 213326 -7622 213562 -7386
rect 213646 -7622 213882 -7386
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 222326 223718 222562 223954
rect 222646 223718 222882 223954
rect 222326 223398 222562 223634
rect 222646 223398 222882 223634
rect 222326 187718 222562 187954
rect 222646 187718 222882 187954
rect 222326 187398 222562 187634
rect 222646 187398 222882 187634
rect 222326 151718 222562 151954
rect 222646 151718 222882 151954
rect 222326 151398 222562 151634
rect 222646 151398 222882 151634
rect 222326 115718 222562 115954
rect 222646 115718 222882 115954
rect 222326 115398 222562 115634
rect 222646 115398 222882 115634
rect 222326 79718 222562 79954
rect 222646 79718 222882 79954
rect 222326 79398 222562 79634
rect 222646 79398 222882 79634
rect 222326 43718 222562 43954
rect 222646 43718 222882 43954
rect 222326 43398 222562 43634
rect 222646 43398 222882 43634
rect 222326 7718 222562 7954
rect 222646 7718 222882 7954
rect 222326 7398 222562 7634
rect 222646 7398 222882 7634
rect 222326 -1542 222562 -1306
rect 222646 -1542 222882 -1306
rect 222326 -1862 222562 -1626
rect 222646 -1862 222882 -1626
rect 226826 228217 227062 228453
rect 227146 228217 227382 228453
rect 226826 227897 227062 228133
rect 227146 227897 227382 228133
rect 226826 192218 227062 192454
rect 227146 192218 227382 192454
rect 226826 191898 227062 192134
rect 227146 191898 227382 192134
rect 226826 156218 227062 156454
rect 227146 156218 227382 156454
rect 226826 155898 227062 156134
rect 227146 155898 227382 156134
rect 226826 120218 227062 120454
rect 227146 120218 227382 120454
rect 226826 119898 227062 120134
rect 227146 119898 227382 120134
rect 226826 84218 227062 84454
rect 227146 84218 227382 84454
rect 226826 83898 227062 84134
rect 227146 83898 227382 84134
rect 226826 48218 227062 48454
rect 227146 48218 227382 48454
rect 226826 47898 227062 48134
rect 227146 47898 227382 48134
rect 226826 12218 227062 12454
rect 227146 12218 227382 12454
rect 226826 11898 227062 12134
rect 227146 11898 227382 12134
rect 226826 -2502 227062 -2266
rect 227146 -2502 227382 -2266
rect 226826 -2822 227062 -2586
rect 227146 -2822 227382 -2586
rect 231326 196718 231562 196954
rect 231646 196718 231882 196954
rect 231326 196398 231562 196634
rect 231646 196398 231882 196634
rect 231326 160718 231562 160954
rect 231646 160718 231882 160954
rect 231326 160398 231562 160634
rect 231646 160398 231882 160634
rect 231326 124718 231562 124954
rect 231646 124718 231882 124954
rect 231326 124398 231562 124634
rect 231646 124398 231882 124634
rect 231326 88718 231562 88954
rect 231646 88718 231882 88954
rect 231326 88398 231562 88634
rect 231646 88398 231882 88634
rect 231326 52718 231562 52954
rect 231646 52718 231882 52954
rect 231326 52398 231562 52634
rect 231646 52398 231882 52634
rect 231326 16718 231562 16954
rect 231646 16718 231882 16954
rect 231326 16398 231562 16634
rect 231646 16398 231882 16634
rect 231326 -3462 231562 -3226
rect 231646 -3462 231882 -3226
rect 231326 -3782 231562 -3546
rect 231646 -3782 231882 -3546
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -4422 236062 -4186
rect 236146 -4422 236382 -4186
rect 235826 -4742 236062 -4506
rect 236146 -4742 236382 -4506
rect 240326 205718 240562 205954
rect 240646 205718 240882 205954
rect 240326 205398 240562 205634
rect 240646 205398 240882 205634
rect 240326 169718 240562 169954
rect 240646 169718 240882 169954
rect 240326 169398 240562 169634
rect 240646 169398 240882 169634
rect 240326 133718 240562 133954
rect 240646 133718 240882 133954
rect 240326 133398 240562 133634
rect 240646 133398 240882 133634
rect 240326 97718 240562 97954
rect 240646 97718 240882 97954
rect 240326 97398 240562 97634
rect 240646 97398 240882 97634
rect 240326 61718 240562 61954
rect 240646 61718 240882 61954
rect 240326 61398 240562 61634
rect 240646 61398 240882 61634
rect 240326 25718 240562 25954
rect 240646 25718 240882 25954
rect 240326 25398 240562 25634
rect 240646 25398 240882 25634
rect 240326 -5382 240562 -5146
rect 240646 -5382 240882 -5146
rect 240326 -5702 240562 -5466
rect 240646 -5702 240882 -5466
rect 244826 210218 245062 210454
rect 245146 210218 245382 210454
rect 244826 209898 245062 210134
rect 245146 209898 245382 210134
rect 244826 174218 245062 174454
rect 245146 174218 245382 174454
rect 244826 173898 245062 174134
rect 245146 173898 245382 174134
rect 244826 138218 245062 138454
rect 245146 138218 245382 138454
rect 244826 137898 245062 138134
rect 245146 137898 245382 138134
rect 244826 102218 245062 102454
rect 245146 102218 245382 102454
rect 244826 101898 245062 102134
rect 245146 101898 245382 102134
rect 244826 66218 245062 66454
rect 245146 66218 245382 66454
rect 244826 65898 245062 66134
rect 245146 65898 245382 66134
rect 244826 30218 245062 30454
rect 245146 30218 245382 30454
rect 244826 29898 245062 30134
rect 245146 29898 245382 30134
rect 244826 -6342 245062 -6106
rect 245146 -6342 245382 -6106
rect 244826 -6662 245062 -6426
rect 245146 -6662 245382 -6426
rect 249326 214718 249562 214954
rect 249646 214718 249882 214954
rect 249326 214398 249562 214634
rect 249646 214398 249882 214634
rect 249326 178718 249562 178954
rect 249646 178718 249882 178954
rect 249326 178398 249562 178634
rect 249646 178398 249882 178634
rect 249326 142718 249562 142954
rect 249646 142718 249882 142954
rect 249326 142398 249562 142634
rect 249646 142398 249882 142634
rect 249326 106718 249562 106954
rect 249646 106718 249882 106954
rect 249326 106398 249562 106634
rect 249646 106398 249882 106634
rect 249326 70718 249562 70954
rect 249646 70718 249882 70954
rect 249326 70398 249562 70634
rect 249646 70398 249882 70634
rect 249326 34718 249562 34954
rect 249646 34718 249882 34954
rect 249326 34398 249562 34634
rect 249646 34398 249882 34634
rect 249326 -7302 249562 -7066
rect 249646 -7302 249882 -7066
rect 249326 -7622 249562 -7386
rect 249646 -7622 249882 -7386
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 258326 223718 258562 223954
rect 258646 223718 258882 223954
rect 258326 223398 258562 223634
rect 258646 223398 258882 223634
rect 258326 187718 258562 187954
rect 258646 187718 258882 187954
rect 258326 187398 258562 187634
rect 258646 187398 258882 187634
rect 258326 151718 258562 151954
rect 258646 151718 258882 151954
rect 258326 151398 258562 151634
rect 258646 151398 258882 151634
rect 258326 115718 258562 115954
rect 258646 115718 258882 115954
rect 258326 115398 258562 115634
rect 258646 115398 258882 115634
rect 258326 79718 258562 79954
rect 258646 79718 258882 79954
rect 258326 79398 258562 79634
rect 258646 79398 258882 79634
rect 258326 43718 258562 43954
rect 258646 43718 258882 43954
rect 258326 43398 258562 43634
rect 258646 43398 258882 43634
rect 258326 7718 258562 7954
rect 258646 7718 258882 7954
rect 258326 7398 258562 7634
rect 258646 7398 258882 7634
rect 258326 -1542 258562 -1306
rect 258646 -1542 258882 -1306
rect 258326 -1862 258562 -1626
rect 258646 -1862 258882 -1626
rect 262826 228217 263062 228453
rect 263146 228217 263382 228453
rect 262826 227897 263062 228133
rect 263146 227897 263382 228133
rect 262826 192218 263062 192454
rect 263146 192218 263382 192454
rect 262826 191898 263062 192134
rect 263146 191898 263382 192134
rect 262826 156218 263062 156454
rect 263146 156218 263382 156454
rect 262826 155898 263062 156134
rect 263146 155898 263382 156134
rect 262826 120218 263062 120454
rect 263146 120218 263382 120454
rect 262826 119898 263062 120134
rect 263146 119898 263382 120134
rect 262826 84218 263062 84454
rect 263146 84218 263382 84454
rect 262826 83898 263062 84134
rect 263146 83898 263382 84134
rect 262826 48218 263062 48454
rect 263146 48218 263382 48454
rect 262826 47898 263062 48134
rect 263146 47898 263382 48134
rect 262826 12218 263062 12454
rect 263146 12218 263382 12454
rect 262826 11898 263062 12134
rect 263146 11898 263382 12134
rect 262826 -2502 263062 -2266
rect 263146 -2502 263382 -2266
rect 262826 -2822 263062 -2586
rect 263146 -2822 263382 -2586
rect 267326 196718 267562 196954
rect 267646 196718 267882 196954
rect 267326 196398 267562 196634
rect 267646 196398 267882 196634
rect 267326 160718 267562 160954
rect 267646 160718 267882 160954
rect 267326 160398 267562 160634
rect 267646 160398 267882 160634
rect 267326 124718 267562 124954
rect 267646 124718 267882 124954
rect 267326 124398 267562 124634
rect 267646 124398 267882 124634
rect 267326 88718 267562 88954
rect 267646 88718 267882 88954
rect 267326 88398 267562 88634
rect 267646 88398 267882 88634
rect 267326 52718 267562 52954
rect 267646 52718 267882 52954
rect 267326 52398 267562 52634
rect 267646 52398 267882 52634
rect 267326 16718 267562 16954
rect 267646 16718 267882 16954
rect 267326 16398 267562 16634
rect 267646 16398 267882 16634
rect 267326 -3462 267562 -3226
rect 267646 -3462 267882 -3226
rect 267326 -3782 267562 -3546
rect 267646 -3782 267882 -3546
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -4422 272062 -4186
rect 272146 -4422 272382 -4186
rect 271826 -4742 272062 -4506
rect 272146 -4742 272382 -4506
rect 276326 205718 276562 205954
rect 276646 205718 276882 205954
rect 276326 205398 276562 205634
rect 276646 205398 276882 205634
rect 276326 169718 276562 169954
rect 276646 169718 276882 169954
rect 276326 169398 276562 169634
rect 276646 169398 276882 169634
rect 276326 133718 276562 133954
rect 276646 133718 276882 133954
rect 276326 133398 276562 133634
rect 276646 133398 276882 133634
rect 276326 97718 276562 97954
rect 276646 97718 276882 97954
rect 276326 97398 276562 97634
rect 276646 97398 276882 97634
rect 276326 61718 276562 61954
rect 276646 61718 276882 61954
rect 276326 61398 276562 61634
rect 276646 61398 276882 61634
rect 276326 25718 276562 25954
rect 276646 25718 276882 25954
rect 276326 25398 276562 25634
rect 276646 25398 276882 25634
rect 276326 -5382 276562 -5146
rect 276646 -5382 276882 -5146
rect 276326 -5702 276562 -5466
rect 276646 -5702 276882 -5466
rect 280826 210218 281062 210454
rect 281146 210218 281382 210454
rect 280826 209898 281062 210134
rect 281146 209898 281382 210134
rect 280826 174218 281062 174454
rect 281146 174218 281382 174454
rect 280826 173898 281062 174134
rect 281146 173898 281382 174134
rect 280826 138218 281062 138454
rect 281146 138218 281382 138454
rect 280826 137898 281062 138134
rect 281146 137898 281382 138134
rect 280826 102218 281062 102454
rect 281146 102218 281382 102454
rect 280826 101898 281062 102134
rect 281146 101898 281382 102134
rect 280826 66218 281062 66454
rect 281146 66218 281382 66454
rect 280826 65898 281062 66134
rect 281146 65898 281382 66134
rect 280826 30218 281062 30454
rect 281146 30218 281382 30454
rect 280826 29898 281062 30134
rect 281146 29898 281382 30134
rect 280826 -6342 281062 -6106
rect 281146 -6342 281382 -6106
rect 280826 -6662 281062 -6426
rect 281146 -6662 281382 -6426
rect 285326 214718 285562 214954
rect 285646 214718 285882 214954
rect 285326 214398 285562 214634
rect 285646 214398 285882 214634
rect 285326 178718 285562 178954
rect 285646 178718 285882 178954
rect 285326 178398 285562 178634
rect 285646 178398 285882 178634
rect 285326 142718 285562 142954
rect 285646 142718 285882 142954
rect 285326 142398 285562 142634
rect 285646 142398 285882 142634
rect 285326 106718 285562 106954
rect 285646 106718 285882 106954
rect 285326 106398 285562 106634
rect 285646 106398 285882 106634
rect 285326 70718 285562 70954
rect 285646 70718 285882 70954
rect 285326 70398 285562 70634
rect 285646 70398 285882 70634
rect 285326 34718 285562 34954
rect 285646 34718 285882 34954
rect 285326 34398 285562 34634
rect 285646 34398 285882 34634
rect 285326 -7302 285562 -7066
rect 285646 -7302 285882 -7066
rect 285326 -7622 285562 -7386
rect 285646 -7622 285882 -7386
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 294326 223718 294562 223954
rect 294646 223718 294882 223954
rect 294326 223398 294562 223634
rect 294646 223398 294882 223634
rect 294326 187718 294562 187954
rect 294646 187718 294882 187954
rect 294326 187398 294562 187634
rect 294646 187398 294882 187634
rect 294326 151718 294562 151954
rect 294646 151718 294882 151954
rect 294326 151398 294562 151634
rect 294646 151398 294882 151634
rect 294326 115718 294562 115954
rect 294646 115718 294882 115954
rect 294326 115398 294562 115634
rect 294646 115398 294882 115634
rect 294326 79718 294562 79954
rect 294646 79718 294882 79954
rect 294326 79398 294562 79634
rect 294646 79398 294882 79634
rect 294326 43718 294562 43954
rect 294646 43718 294882 43954
rect 294326 43398 294562 43634
rect 294646 43398 294882 43634
rect 294326 7718 294562 7954
rect 294646 7718 294882 7954
rect 294326 7398 294562 7634
rect 294646 7398 294882 7634
rect 294326 -1542 294562 -1306
rect 294646 -1542 294882 -1306
rect 294326 -1862 294562 -1626
rect 294646 -1862 294882 -1626
rect 298826 228217 299062 228453
rect 299146 228217 299382 228453
rect 298826 227897 299062 228133
rect 299146 227897 299382 228133
rect 298826 192218 299062 192454
rect 299146 192218 299382 192454
rect 298826 191898 299062 192134
rect 299146 191898 299382 192134
rect 298826 156218 299062 156454
rect 299146 156218 299382 156454
rect 298826 155898 299062 156134
rect 299146 155898 299382 156134
rect 298826 120218 299062 120454
rect 299146 120218 299382 120454
rect 298826 119898 299062 120134
rect 299146 119898 299382 120134
rect 298826 84218 299062 84454
rect 299146 84218 299382 84454
rect 298826 83898 299062 84134
rect 299146 83898 299382 84134
rect 298826 48218 299062 48454
rect 299146 48218 299382 48454
rect 298826 47898 299062 48134
rect 299146 47898 299382 48134
rect 298826 12218 299062 12454
rect 299146 12218 299382 12454
rect 298826 11898 299062 12134
rect 299146 11898 299382 12134
rect 298826 -2502 299062 -2266
rect 299146 -2502 299382 -2266
rect 298826 -2822 299062 -2586
rect 299146 -2822 299382 -2586
rect 303326 196718 303562 196954
rect 303646 196718 303882 196954
rect 303326 196398 303562 196634
rect 303646 196398 303882 196634
rect 303326 160718 303562 160954
rect 303646 160718 303882 160954
rect 303326 160398 303562 160634
rect 303646 160398 303882 160634
rect 303326 124718 303562 124954
rect 303646 124718 303882 124954
rect 303326 124398 303562 124634
rect 303646 124398 303882 124634
rect 303326 88718 303562 88954
rect 303646 88718 303882 88954
rect 303326 88398 303562 88634
rect 303646 88398 303882 88634
rect 303326 52718 303562 52954
rect 303646 52718 303882 52954
rect 303326 52398 303562 52634
rect 303646 52398 303882 52634
rect 303326 16718 303562 16954
rect 303646 16718 303882 16954
rect 303326 16398 303562 16634
rect 303646 16398 303882 16634
rect 303326 -3462 303562 -3226
rect 303646 -3462 303882 -3226
rect 303326 -3782 303562 -3546
rect 303646 -3782 303882 -3546
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -4422 308062 -4186
rect 308146 -4422 308382 -4186
rect 307826 -4742 308062 -4506
rect 308146 -4742 308382 -4506
rect 312326 205718 312562 205954
rect 312646 205718 312882 205954
rect 312326 205398 312562 205634
rect 312646 205398 312882 205634
rect 312326 169718 312562 169954
rect 312646 169718 312882 169954
rect 312326 169398 312562 169634
rect 312646 169398 312882 169634
rect 312326 133718 312562 133954
rect 312646 133718 312882 133954
rect 312326 133398 312562 133634
rect 312646 133398 312882 133634
rect 312326 97718 312562 97954
rect 312646 97718 312882 97954
rect 312326 97398 312562 97634
rect 312646 97398 312882 97634
rect 312326 61718 312562 61954
rect 312646 61718 312882 61954
rect 312326 61398 312562 61634
rect 312646 61398 312882 61634
rect 312326 25718 312562 25954
rect 312646 25718 312882 25954
rect 312326 25398 312562 25634
rect 312646 25398 312882 25634
rect 312326 -5382 312562 -5146
rect 312646 -5382 312882 -5146
rect 312326 -5702 312562 -5466
rect 312646 -5702 312882 -5466
rect 316826 210218 317062 210454
rect 317146 210218 317382 210454
rect 316826 209898 317062 210134
rect 317146 209898 317382 210134
rect 316826 174218 317062 174454
rect 317146 174218 317382 174454
rect 316826 173898 317062 174134
rect 317146 173898 317382 174134
rect 316826 138218 317062 138454
rect 317146 138218 317382 138454
rect 316826 137898 317062 138134
rect 317146 137898 317382 138134
rect 316826 102218 317062 102454
rect 317146 102218 317382 102454
rect 316826 101898 317062 102134
rect 317146 101898 317382 102134
rect 316826 66218 317062 66454
rect 317146 66218 317382 66454
rect 316826 65898 317062 66134
rect 317146 65898 317382 66134
rect 316826 30218 317062 30454
rect 317146 30218 317382 30454
rect 316826 29898 317062 30134
rect 317146 29898 317382 30134
rect 316826 -6342 317062 -6106
rect 317146 -6342 317382 -6106
rect 316826 -6662 317062 -6426
rect 317146 -6662 317382 -6426
rect 321326 214718 321562 214954
rect 321646 214718 321882 214954
rect 321326 214398 321562 214634
rect 321646 214398 321882 214634
rect 321326 178718 321562 178954
rect 321646 178718 321882 178954
rect 321326 178398 321562 178634
rect 321646 178398 321882 178634
rect 321326 142718 321562 142954
rect 321646 142718 321882 142954
rect 321326 142398 321562 142634
rect 321646 142398 321882 142634
rect 321326 106718 321562 106954
rect 321646 106718 321882 106954
rect 321326 106398 321562 106634
rect 321646 106398 321882 106634
rect 321326 70718 321562 70954
rect 321646 70718 321882 70954
rect 321326 70398 321562 70634
rect 321646 70398 321882 70634
rect 321326 34718 321562 34954
rect 321646 34718 321882 34954
rect 321326 34398 321562 34634
rect 321646 34398 321882 34634
rect 321326 -7302 321562 -7066
rect 321646 -7302 321882 -7066
rect 321326 -7622 321562 -7386
rect 321646 -7622 321882 -7386
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 330326 223718 330562 223954
rect 330646 223718 330882 223954
rect 330326 223398 330562 223634
rect 330646 223398 330882 223634
rect 330326 187718 330562 187954
rect 330646 187718 330882 187954
rect 330326 187398 330562 187634
rect 330646 187398 330882 187634
rect 330326 151718 330562 151954
rect 330646 151718 330882 151954
rect 330326 151398 330562 151634
rect 330646 151398 330882 151634
rect 330326 115718 330562 115954
rect 330646 115718 330882 115954
rect 330326 115398 330562 115634
rect 330646 115398 330882 115634
rect 330326 79718 330562 79954
rect 330646 79718 330882 79954
rect 330326 79398 330562 79634
rect 330646 79398 330882 79634
rect 330326 43718 330562 43954
rect 330646 43718 330882 43954
rect 330326 43398 330562 43634
rect 330646 43398 330882 43634
rect 330326 7718 330562 7954
rect 330646 7718 330882 7954
rect 330326 7398 330562 7634
rect 330646 7398 330882 7634
rect 330326 -1542 330562 -1306
rect 330646 -1542 330882 -1306
rect 330326 -1862 330562 -1626
rect 330646 -1862 330882 -1626
rect 334826 228217 335062 228453
rect 335146 228217 335382 228453
rect 334826 227897 335062 228133
rect 335146 227897 335382 228133
rect 334826 192218 335062 192454
rect 335146 192218 335382 192454
rect 334826 191898 335062 192134
rect 335146 191898 335382 192134
rect 334826 156218 335062 156454
rect 335146 156218 335382 156454
rect 334826 155898 335062 156134
rect 335146 155898 335382 156134
rect 334826 120218 335062 120454
rect 335146 120218 335382 120454
rect 334826 119898 335062 120134
rect 335146 119898 335382 120134
rect 334826 84218 335062 84454
rect 335146 84218 335382 84454
rect 334826 83898 335062 84134
rect 335146 83898 335382 84134
rect 334826 48218 335062 48454
rect 335146 48218 335382 48454
rect 334826 47898 335062 48134
rect 335146 47898 335382 48134
rect 334826 12218 335062 12454
rect 335146 12218 335382 12454
rect 334826 11898 335062 12134
rect 335146 11898 335382 12134
rect 334826 -2502 335062 -2266
rect 335146 -2502 335382 -2266
rect 334826 -2822 335062 -2586
rect 335146 -2822 335382 -2586
rect 339326 196718 339562 196954
rect 339646 196718 339882 196954
rect 339326 196398 339562 196634
rect 339646 196398 339882 196634
rect 339326 160718 339562 160954
rect 339646 160718 339882 160954
rect 339326 160398 339562 160634
rect 339646 160398 339882 160634
rect 339326 124718 339562 124954
rect 339646 124718 339882 124954
rect 339326 124398 339562 124634
rect 339646 124398 339882 124634
rect 339326 88718 339562 88954
rect 339646 88718 339882 88954
rect 339326 88398 339562 88634
rect 339646 88398 339882 88634
rect 339326 52718 339562 52954
rect 339646 52718 339882 52954
rect 339326 52398 339562 52634
rect 339646 52398 339882 52634
rect 339326 16718 339562 16954
rect 339646 16718 339882 16954
rect 339326 16398 339562 16634
rect 339646 16398 339882 16634
rect 339326 -3462 339562 -3226
rect 339646 -3462 339882 -3226
rect 339326 -3782 339562 -3546
rect 339646 -3782 339882 -3546
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -4422 344062 -4186
rect 344146 -4422 344382 -4186
rect 343826 -4742 344062 -4506
rect 344146 -4742 344382 -4506
rect 348326 205718 348562 205954
rect 348646 205718 348882 205954
rect 348326 205398 348562 205634
rect 348646 205398 348882 205634
rect 348326 169718 348562 169954
rect 348646 169718 348882 169954
rect 348326 169398 348562 169634
rect 348646 169398 348882 169634
rect 348326 133718 348562 133954
rect 348646 133718 348882 133954
rect 348326 133398 348562 133634
rect 348646 133398 348882 133634
rect 348326 97718 348562 97954
rect 348646 97718 348882 97954
rect 348326 97398 348562 97634
rect 348646 97398 348882 97634
rect 348326 61718 348562 61954
rect 348646 61718 348882 61954
rect 348326 61398 348562 61634
rect 348646 61398 348882 61634
rect 348326 25718 348562 25954
rect 348646 25718 348882 25954
rect 348326 25398 348562 25634
rect 348646 25398 348882 25634
rect 348326 -5382 348562 -5146
rect 348646 -5382 348882 -5146
rect 348326 -5702 348562 -5466
rect 348646 -5702 348882 -5466
rect 352826 210218 353062 210454
rect 353146 210218 353382 210454
rect 352826 209898 353062 210134
rect 353146 209898 353382 210134
rect 352826 174218 353062 174454
rect 353146 174218 353382 174454
rect 352826 173898 353062 174134
rect 353146 173898 353382 174134
rect 352826 138218 353062 138454
rect 353146 138218 353382 138454
rect 352826 137898 353062 138134
rect 353146 137898 353382 138134
rect 352826 102218 353062 102454
rect 353146 102218 353382 102454
rect 352826 101898 353062 102134
rect 353146 101898 353382 102134
rect 352826 66218 353062 66454
rect 353146 66218 353382 66454
rect 352826 65898 353062 66134
rect 353146 65898 353382 66134
rect 352826 30218 353062 30454
rect 353146 30218 353382 30454
rect 352826 29898 353062 30134
rect 353146 29898 353382 30134
rect 352826 -6342 353062 -6106
rect 353146 -6342 353382 -6106
rect 352826 -6662 353062 -6426
rect 353146 -6662 353382 -6426
rect 357326 214718 357562 214954
rect 357646 214718 357882 214954
rect 357326 214398 357562 214634
rect 357646 214398 357882 214634
rect 357326 178718 357562 178954
rect 357646 178718 357882 178954
rect 357326 178398 357562 178634
rect 357646 178398 357882 178634
rect 357326 142718 357562 142954
rect 357646 142718 357882 142954
rect 357326 142398 357562 142634
rect 357646 142398 357882 142634
rect 357326 106718 357562 106954
rect 357646 106718 357882 106954
rect 357326 106398 357562 106634
rect 357646 106398 357882 106634
rect 357326 70718 357562 70954
rect 357646 70718 357882 70954
rect 357326 70398 357562 70634
rect 357646 70398 357882 70634
rect 357326 34718 357562 34954
rect 357646 34718 357882 34954
rect 357326 34398 357562 34634
rect 357646 34398 357882 34634
rect 357326 -7302 357562 -7066
rect 357646 -7302 357882 -7066
rect 357326 -7622 357562 -7386
rect 357646 -7622 357882 -7386
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 366326 223718 366562 223954
rect 366646 223718 366882 223954
rect 366326 223398 366562 223634
rect 366646 223398 366882 223634
rect 366326 187718 366562 187954
rect 366646 187718 366882 187954
rect 366326 187398 366562 187634
rect 366646 187398 366882 187634
rect 366326 151718 366562 151954
rect 366646 151718 366882 151954
rect 366326 151398 366562 151634
rect 366646 151398 366882 151634
rect 366326 115718 366562 115954
rect 366646 115718 366882 115954
rect 366326 115398 366562 115634
rect 366646 115398 366882 115634
rect 366326 79718 366562 79954
rect 366646 79718 366882 79954
rect 366326 79398 366562 79634
rect 366646 79398 366882 79634
rect 366326 43718 366562 43954
rect 366646 43718 366882 43954
rect 366326 43398 366562 43634
rect 366646 43398 366882 43634
rect 366326 7718 366562 7954
rect 366646 7718 366882 7954
rect 366326 7398 366562 7634
rect 366646 7398 366882 7634
rect 366326 -1542 366562 -1306
rect 366646 -1542 366882 -1306
rect 366326 -1862 366562 -1626
rect 366646 -1862 366882 -1626
rect 370826 228217 371062 228453
rect 371146 228217 371382 228453
rect 370826 227897 371062 228133
rect 371146 227897 371382 228133
rect 370826 192218 371062 192454
rect 371146 192218 371382 192454
rect 370826 191898 371062 192134
rect 371146 191898 371382 192134
rect 370826 156218 371062 156454
rect 371146 156218 371382 156454
rect 370826 155898 371062 156134
rect 371146 155898 371382 156134
rect 370826 120218 371062 120454
rect 371146 120218 371382 120454
rect 370826 119898 371062 120134
rect 371146 119898 371382 120134
rect 370826 84218 371062 84454
rect 371146 84218 371382 84454
rect 370826 83898 371062 84134
rect 371146 83898 371382 84134
rect 370826 48218 371062 48454
rect 371146 48218 371382 48454
rect 370826 47898 371062 48134
rect 371146 47898 371382 48134
rect 370826 12218 371062 12454
rect 371146 12218 371382 12454
rect 370826 11898 371062 12134
rect 371146 11898 371382 12134
rect 370826 -2502 371062 -2266
rect 371146 -2502 371382 -2266
rect 370826 -2822 371062 -2586
rect 371146 -2822 371382 -2586
rect 375326 196718 375562 196954
rect 375646 196718 375882 196954
rect 375326 196398 375562 196634
rect 375646 196398 375882 196634
rect 375326 160718 375562 160954
rect 375646 160718 375882 160954
rect 375326 160398 375562 160634
rect 375646 160398 375882 160634
rect 375326 124718 375562 124954
rect 375646 124718 375882 124954
rect 375326 124398 375562 124634
rect 375646 124398 375882 124634
rect 375326 88718 375562 88954
rect 375646 88718 375882 88954
rect 375326 88398 375562 88634
rect 375646 88398 375882 88634
rect 375326 52718 375562 52954
rect 375646 52718 375882 52954
rect 375326 52398 375562 52634
rect 375646 52398 375882 52634
rect 375326 16718 375562 16954
rect 375646 16718 375882 16954
rect 375326 16398 375562 16634
rect 375646 16398 375882 16634
rect 375326 -3462 375562 -3226
rect 375646 -3462 375882 -3226
rect 375326 -3782 375562 -3546
rect 375646 -3782 375882 -3546
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -4422 380062 -4186
rect 380146 -4422 380382 -4186
rect 379826 -4742 380062 -4506
rect 380146 -4742 380382 -4506
rect 384326 205718 384562 205954
rect 384646 205718 384882 205954
rect 384326 205398 384562 205634
rect 384646 205398 384882 205634
rect 384326 169718 384562 169954
rect 384646 169718 384882 169954
rect 384326 169398 384562 169634
rect 384646 169398 384882 169634
rect 384326 133718 384562 133954
rect 384646 133718 384882 133954
rect 384326 133398 384562 133634
rect 384646 133398 384882 133634
rect 384326 97718 384562 97954
rect 384646 97718 384882 97954
rect 384326 97398 384562 97634
rect 384646 97398 384882 97634
rect 384326 61718 384562 61954
rect 384646 61718 384882 61954
rect 384326 61398 384562 61634
rect 384646 61398 384882 61634
rect 384326 25718 384562 25954
rect 384646 25718 384882 25954
rect 384326 25398 384562 25634
rect 384646 25398 384882 25634
rect 384326 -5382 384562 -5146
rect 384646 -5382 384882 -5146
rect 384326 -5702 384562 -5466
rect 384646 -5702 384882 -5466
rect 388826 210218 389062 210454
rect 389146 210218 389382 210454
rect 388826 209898 389062 210134
rect 389146 209898 389382 210134
rect 388826 174218 389062 174454
rect 389146 174218 389382 174454
rect 388826 173898 389062 174134
rect 389146 173898 389382 174134
rect 388826 138218 389062 138454
rect 389146 138218 389382 138454
rect 388826 137898 389062 138134
rect 389146 137898 389382 138134
rect 388826 102218 389062 102454
rect 389146 102218 389382 102454
rect 388826 101898 389062 102134
rect 389146 101898 389382 102134
rect 388826 66218 389062 66454
rect 389146 66218 389382 66454
rect 388826 65898 389062 66134
rect 389146 65898 389382 66134
rect 388826 30218 389062 30454
rect 389146 30218 389382 30454
rect 388826 29898 389062 30134
rect 389146 29898 389382 30134
rect 388826 -6342 389062 -6106
rect 389146 -6342 389382 -6106
rect 388826 -6662 389062 -6426
rect 389146 -6662 389382 -6426
rect 393326 214718 393562 214954
rect 393646 214718 393882 214954
rect 393326 214398 393562 214634
rect 393646 214398 393882 214634
rect 393326 178718 393562 178954
rect 393646 178718 393882 178954
rect 393326 178398 393562 178634
rect 393646 178398 393882 178634
rect 393326 142718 393562 142954
rect 393646 142718 393882 142954
rect 393326 142398 393562 142634
rect 393646 142398 393882 142634
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 402326 705562 402562 705798
rect 402646 705562 402882 705798
rect 402326 705242 402562 705478
rect 402646 705242 402882 705478
rect 402326 691718 402562 691954
rect 402646 691718 402882 691954
rect 402326 691398 402562 691634
rect 402646 691398 402882 691634
rect 402326 655718 402562 655954
rect 402646 655718 402882 655954
rect 402326 655398 402562 655634
rect 402646 655398 402882 655634
rect 402326 619718 402562 619954
rect 402646 619718 402882 619954
rect 402326 619398 402562 619634
rect 402646 619398 402882 619634
rect 402326 583718 402562 583954
rect 402646 583718 402882 583954
rect 402326 583398 402562 583634
rect 402646 583398 402882 583634
rect 402326 547718 402562 547954
rect 402646 547718 402882 547954
rect 402326 547398 402562 547634
rect 402646 547398 402882 547634
rect 402326 511718 402562 511954
rect 402646 511718 402882 511954
rect 402326 511398 402562 511634
rect 402646 511398 402882 511634
rect 402326 475718 402562 475954
rect 402646 475718 402882 475954
rect 402326 475398 402562 475634
rect 402646 475398 402882 475634
rect 402326 439718 402562 439954
rect 402646 439718 402882 439954
rect 402326 439398 402562 439634
rect 402646 439398 402882 439634
rect 402326 403718 402562 403954
rect 402646 403718 402882 403954
rect 402326 403398 402562 403634
rect 402646 403398 402882 403634
rect 402326 367718 402562 367954
rect 402646 367718 402882 367954
rect 402326 367398 402562 367634
rect 402646 367398 402882 367634
rect 402326 331718 402562 331954
rect 402646 331718 402882 331954
rect 402326 331398 402562 331634
rect 402646 331398 402882 331634
rect 402326 295718 402562 295954
rect 402646 295718 402882 295954
rect 402326 295398 402562 295634
rect 402646 295398 402882 295634
rect 402326 259718 402562 259954
rect 402646 259718 402882 259954
rect 402326 259398 402562 259634
rect 402646 259398 402882 259634
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 393326 106718 393562 106954
rect 393646 106718 393882 106954
rect 393326 106398 393562 106634
rect 393646 106398 393882 106634
rect 393326 70718 393562 70954
rect 393646 70718 393882 70954
rect 393326 70398 393562 70634
rect 393646 70398 393882 70634
rect 393326 34718 393562 34954
rect 393646 34718 393882 34954
rect 393326 34398 393562 34634
rect 393646 34398 393882 34634
rect 393326 -7302 393562 -7066
rect 393646 -7302 393882 -7066
rect 393326 -7622 393562 -7386
rect 393646 -7622 393882 -7386
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 402326 223718 402562 223954
rect 402646 223718 402882 223954
rect 402326 223398 402562 223634
rect 402646 223398 402882 223634
rect 402326 187718 402562 187954
rect 402646 187718 402882 187954
rect 402326 187398 402562 187634
rect 402646 187398 402882 187634
rect 402326 151718 402562 151954
rect 402646 151718 402882 151954
rect 402326 151398 402562 151634
rect 402646 151398 402882 151634
rect 402326 115718 402562 115954
rect 402646 115718 402882 115954
rect 402326 115398 402562 115634
rect 402646 115398 402882 115634
rect 402326 79718 402562 79954
rect 402646 79718 402882 79954
rect 402326 79398 402562 79634
rect 402646 79398 402882 79634
rect 402326 43718 402562 43954
rect 402646 43718 402882 43954
rect 402326 43398 402562 43634
rect 402646 43398 402882 43634
rect 402326 7718 402562 7954
rect 402646 7718 402882 7954
rect 402326 7398 402562 7634
rect 402646 7398 402882 7634
rect 402326 -1542 402562 -1306
rect 402646 -1542 402882 -1306
rect 402326 -1862 402562 -1626
rect 402646 -1862 402882 -1626
rect 406826 706522 407062 706758
rect 407146 706522 407382 706758
rect 406826 706202 407062 706438
rect 407146 706202 407382 706438
rect 406826 696218 407062 696454
rect 407146 696218 407382 696454
rect 406826 695898 407062 696134
rect 407146 695898 407382 696134
rect 406826 660218 407062 660454
rect 407146 660218 407382 660454
rect 406826 659898 407062 660134
rect 407146 659898 407382 660134
rect 406826 624218 407062 624454
rect 407146 624218 407382 624454
rect 406826 623898 407062 624134
rect 407146 623898 407382 624134
rect 406826 588218 407062 588454
rect 407146 588218 407382 588454
rect 406826 587898 407062 588134
rect 407146 587898 407382 588134
rect 406826 552218 407062 552454
rect 407146 552218 407382 552454
rect 406826 551898 407062 552134
rect 407146 551898 407382 552134
rect 406826 516218 407062 516454
rect 407146 516218 407382 516454
rect 406826 515898 407062 516134
rect 407146 515898 407382 516134
rect 406826 480218 407062 480454
rect 407146 480218 407382 480454
rect 406826 479898 407062 480134
rect 407146 479898 407382 480134
rect 406826 444218 407062 444454
rect 407146 444218 407382 444454
rect 406826 443898 407062 444134
rect 407146 443898 407382 444134
rect 406826 408218 407062 408454
rect 407146 408218 407382 408454
rect 406826 407898 407062 408134
rect 407146 407898 407382 408134
rect 406826 372218 407062 372454
rect 407146 372218 407382 372454
rect 406826 371898 407062 372134
rect 407146 371898 407382 372134
rect 406826 336218 407062 336454
rect 407146 336218 407382 336454
rect 406826 335898 407062 336134
rect 407146 335898 407382 336134
rect 406826 300218 407062 300454
rect 407146 300218 407382 300454
rect 406826 299898 407062 300134
rect 407146 299898 407382 300134
rect 406826 264218 407062 264454
rect 407146 264218 407382 264454
rect 406826 263898 407062 264134
rect 407146 263898 407382 264134
rect 406826 228218 407062 228454
rect 407146 228218 407382 228454
rect 406826 227898 407062 228134
rect 407146 227898 407382 228134
rect 406826 192218 407062 192454
rect 407146 192218 407382 192454
rect 406826 191898 407062 192134
rect 407146 191898 407382 192134
rect 406826 156218 407062 156454
rect 407146 156218 407382 156454
rect 406826 155898 407062 156134
rect 407146 155898 407382 156134
rect 406826 120218 407062 120454
rect 407146 120218 407382 120454
rect 406826 119898 407062 120134
rect 407146 119898 407382 120134
rect 406826 84218 407062 84454
rect 407146 84218 407382 84454
rect 406826 83898 407062 84134
rect 407146 83898 407382 84134
rect 406826 48218 407062 48454
rect 407146 48218 407382 48454
rect 406826 47898 407062 48134
rect 407146 47898 407382 48134
rect 406826 12218 407062 12454
rect 407146 12218 407382 12454
rect 406826 11898 407062 12134
rect 407146 11898 407382 12134
rect 406826 -2502 407062 -2266
rect 407146 -2502 407382 -2266
rect 406826 -2822 407062 -2586
rect 407146 -2822 407382 -2586
rect 411326 707482 411562 707718
rect 411646 707482 411882 707718
rect 411326 707162 411562 707398
rect 411646 707162 411882 707398
rect 411326 700718 411562 700954
rect 411646 700718 411882 700954
rect 411326 700398 411562 700634
rect 411646 700398 411882 700634
rect 411326 664718 411562 664954
rect 411646 664718 411882 664954
rect 411326 664398 411562 664634
rect 411646 664398 411882 664634
rect 411326 628718 411562 628954
rect 411646 628718 411882 628954
rect 411326 628398 411562 628634
rect 411646 628398 411882 628634
rect 411326 592718 411562 592954
rect 411646 592718 411882 592954
rect 411326 592398 411562 592634
rect 411646 592398 411882 592634
rect 411326 556718 411562 556954
rect 411646 556718 411882 556954
rect 411326 556398 411562 556634
rect 411646 556398 411882 556634
rect 411326 520718 411562 520954
rect 411646 520718 411882 520954
rect 411326 520398 411562 520634
rect 411646 520398 411882 520634
rect 411326 484718 411562 484954
rect 411646 484718 411882 484954
rect 411326 484398 411562 484634
rect 411646 484398 411882 484634
rect 411326 448718 411562 448954
rect 411646 448718 411882 448954
rect 411326 448398 411562 448634
rect 411646 448398 411882 448634
rect 411326 412718 411562 412954
rect 411646 412718 411882 412954
rect 411326 412398 411562 412634
rect 411646 412398 411882 412634
rect 411326 376718 411562 376954
rect 411646 376718 411882 376954
rect 411326 376398 411562 376634
rect 411646 376398 411882 376634
rect 411326 340718 411562 340954
rect 411646 340718 411882 340954
rect 411326 340398 411562 340634
rect 411646 340398 411882 340634
rect 411326 304718 411562 304954
rect 411646 304718 411882 304954
rect 411326 304398 411562 304634
rect 411646 304398 411882 304634
rect 411326 268718 411562 268954
rect 411646 268718 411882 268954
rect 411326 268398 411562 268634
rect 411646 268398 411882 268634
rect 411326 232718 411562 232954
rect 411646 232718 411882 232954
rect 411326 232398 411562 232634
rect 411646 232398 411882 232634
rect 411326 196718 411562 196954
rect 411646 196718 411882 196954
rect 411326 196398 411562 196634
rect 411646 196398 411882 196634
rect 411326 160718 411562 160954
rect 411646 160718 411882 160954
rect 411326 160398 411562 160634
rect 411646 160398 411882 160634
rect 411326 124718 411562 124954
rect 411646 124718 411882 124954
rect 411326 124398 411562 124634
rect 411646 124398 411882 124634
rect 411326 88718 411562 88954
rect 411646 88718 411882 88954
rect 411326 88398 411562 88634
rect 411646 88398 411882 88634
rect 411326 52718 411562 52954
rect 411646 52718 411882 52954
rect 411326 52398 411562 52634
rect 411646 52398 411882 52634
rect 411326 16718 411562 16954
rect 411646 16718 411882 16954
rect 411326 16398 411562 16634
rect 411646 16398 411882 16634
rect 411326 -3462 411562 -3226
rect 411646 -3462 411882 -3226
rect 411326 -3782 411562 -3546
rect 411646 -3782 411882 -3546
rect 415826 708442 416062 708678
rect 416146 708442 416382 708678
rect 415826 708122 416062 708358
rect 416146 708122 416382 708358
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -4422 416062 -4186
rect 416146 -4422 416382 -4186
rect 415826 -4742 416062 -4506
rect 416146 -4742 416382 -4506
rect 420326 709402 420562 709638
rect 420646 709402 420882 709638
rect 420326 709082 420562 709318
rect 420646 709082 420882 709318
rect 420326 673718 420562 673954
rect 420646 673718 420882 673954
rect 420326 673398 420562 673634
rect 420646 673398 420882 673634
rect 420326 637718 420562 637954
rect 420646 637718 420882 637954
rect 420326 637398 420562 637634
rect 420646 637398 420882 637634
rect 420326 601718 420562 601954
rect 420646 601718 420882 601954
rect 420326 601398 420562 601634
rect 420646 601398 420882 601634
rect 420326 565718 420562 565954
rect 420646 565718 420882 565954
rect 420326 565398 420562 565634
rect 420646 565398 420882 565634
rect 420326 529718 420562 529954
rect 420646 529718 420882 529954
rect 420326 529398 420562 529634
rect 420646 529398 420882 529634
rect 420326 493718 420562 493954
rect 420646 493718 420882 493954
rect 420326 493398 420562 493634
rect 420646 493398 420882 493634
rect 420326 457718 420562 457954
rect 420646 457718 420882 457954
rect 420326 457398 420562 457634
rect 420646 457398 420882 457634
rect 420326 421718 420562 421954
rect 420646 421718 420882 421954
rect 420326 421398 420562 421634
rect 420646 421398 420882 421634
rect 420326 385718 420562 385954
rect 420646 385718 420882 385954
rect 420326 385398 420562 385634
rect 420646 385398 420882 385634
rect 420326 349718 420562 349954
rect 420646 349718 420882 349954
rect 420326 349398 420562 349634
rect 420646 349398 420882 349634
rect 420326 313718 420562 313954
rect 420646 313718 420882 313954
rect 420326 313398 420562 313634
rect 420646 313398 420882 313634
rect 420326 277718 420562 277954
rect 420646 277718 420882 277954
rect 420326 277398 420562 277634
rect 420646 277398 420882 277634
rect 420326 241718 420562 241954
rect 420646 241718 420882 241954
rect 420326 241398 420562 241634
rect 420646 241398 420882 241634
rect 420326 205718 420562 205954
rect 420646 205718 420882 205954
rect 420326 205398 420562 205634
rect 420646 205398 420882 205634
rect 420326 169718 420562 169954
rect 420646 169718 420882 169954
rect 420326 169398 420562 169634
rect 420646 169398 420882 169634
rect 420326 133718 420562 133954
rect 420646 133718 420882 133954
rect 420326 133398 420562 133634
rect 420646 133398 420882 133634
rect 420326 97718 420562 97954
rect 420646 97718 420882 97954
rect 420326 97398 420562 97634
rect 420646 97398 420882 97634
rect 420326 61718 420562 61954
rect 420646 61718 420882 61954
rect 420326 61398 420562 61634
rect 420646 61398 420882 61634
rect 420326 25718 420562 25954
rect 420646 25718 420882 25954
rect 420326 25398 420562 25634
rect 420646 25398 420882 25634
rect 420326 -5382 420562 -5146
rect 420646 -5382 420882 -5146
rect 420326 -5702 420562 -5466
rect 420646 -5702 420882 -5466
rect 424826 710362 425062 710598
rect 425146 710362 425382 710598
rect 424826 710042 425062 710278
rect 425146 710042 425382 710278
rect 424826 678218 425062 678454
rect 425146 678218 425382 678454
rect 424826 677898 425062 678134
rect 425146 677898 425382 678134
rect 424826 642218 425062 642454
rect 425146 642218 425382 642454
rect 424826 641898 425062 642134
rect 425146 641898 425382 642134
rect 424826 606218 425062 606454
rect 425146 606218 425382 606454
rect 424826 605898 425062 606134
rect 425146 605898 425382 606134
rect 424826 570218 425062 570454
rect 425146 570218 425382 570454
rect 424826 569898 425062 570134
rect 425146 569898 425382 570134
rect 424826 534218 425062 534454
rect 425146 534218 425382 534454
rect 424826 533898 425062 534134
rect 425146 533898 425382 534134
rect 424826 498218 425062 498454
rect 425146 498218 425382 498454
rect 424826 497898 425062 498134
rect 425146 497898 425382 498134
rect 424826 462218 425062 462454
rect 425146 462218 425382 462454
rect 424826 461898 425062 462134
rect 425146 461898 425382 462134
rect 424826 426218 425062 426454
rect 425146 426218 425382 426454
rect 424826 425898 425062 426134
rect 425146 425898 425382 426134
rect 424826 390218 425062 390454
rect 425146 390218 425382 390454
rect 424826 389898 425062 390134
rect 425146 389898 425382 390134
rect 424826 354218 425062 354454
rect 425146 354218 425382 354454
rect 424826 353898 425062 354134
rect 425146 353898 425382 354134
rect 424826 318218 425062 318454
rect 425146 318218 425382 318454
rect 424826 317898 425062 318134
rect 425146 317898 425382 318134
rect 424826 282218 425062 282454
rect 425146 282218 425382 282454
rect 424826 281898 425062 282134
rect 425146 281898 425382 282134
rect 424826 246218 425062 246454
rect 425146 246218 425382 246454
rect 424826 245898 425062 246134
rect 425146 245898 425382 246134
rect 424826 210218 425062 210454
rect 425146 210218 425382 210454
rect 424826 209898 425062 210134
rect 425146 209898 425382 210134
rect 424826 174218 425062 174454
rect 425146 174218 425382 174454
rect 424826 173898 425062 174134
rect 425146 173898 425382 174134
rect 424826 138218 425062 138454
rect 425146 138218 425382 138454
rect 424826 137898 425062 138134
rect 425146 137898 425382 138134
rect 424826 102218 425062 102454
rect 425146 102218 425382 102454
rect 424826 101898 425062 102134
rect 425146 101898 425382 102134
rect 424826 66218 425062 66454
rect 425146 66218 425382 66454
rect 424826 65898 425062 66134
rect 425146 65898 425382 66134
rect 424826 30218 425062 30454
rect 425146 30218 425382 30454
rect 424826 29898 425062 30134
rect 425146 29898 425382 30134
rect 424826 -6342 425062 -6106
rect 425146 -6342 425382 -6106
rect 424826 -6662 425062 -6426
rect 425146 -6662 425382 -6426
rect 429326 711322 429562 711558
rect 429646 711322 429882 711558
rect 429326 711002 429562 711238
rect 429646 711002 429882 711238
rect 429326 682718 429562 682954
rect 429646 682718 429882 682954
rect 429326 682398 429562 682634
rect 429646 682398 429882 682634
rect 429326 646718 429562 646954
rect 429646 646718 429882 646954
rect 429326 646398 429562 646634
rect 429646 646398 429882 646634
rect 429326 610718 429562 610954
rect 429646 610718 429882 610954
rect 429326 610398 429562 610634
rect 429646 610398 429882 610634
rect 429326 574718 429562 574954
rect 429646 574718 429882 574954
rect 429326 574398 429562 574634
rect 429646 574398 429882 574634
rect 429326 538718 429562 538954
rect 429646 538718 429882 538954
rect 429326 538398 429562 538634
rect 429646 538398 429882 538634
rect 429326 502718 429562 502954
rect 429646 502718 429882 502954
rect 429326 502398 429562 502634
rect 429646 502398 429882 502634
rect 429326 466718 429562 466954
rect 429646 466718 429882 466954
rect 429326 466398 429562 466634
rect 429646 466398 429882 466634
rect 429326 430718 429562 430954
rect 429646 430718 429882 430954
rect 429326 430398 429562 430634
rect 429646 430398 429882 430634
rect 429326 394718 429562 394954
rect 429646 394718 429882 394954
rect 429326 394398 429562 394634
rect 429646 394398 429882 394634
rect 429326 358718 429562 358954
rect 429646 358718 429882 358954
rect 429326 358398 429562 358634
rect 429646 358398 429882 358634
rect 429326 322718 429562 322954
rect 429646 322718 429882 322954
rect 429326 322398 429562 322634
rect 429646 322398 429882 322634
rect 429326 286718 429562 286954
rect 429646 286718 429882 286954
rect 429326 286398 429562 286634
rect 429646 286398 429882 286634
rect 429326 250718 429562 250954
rect 429646 250718 429882 250954
rect 429326 250398 429562 250634
rect 429646 250398 429882 250634
rect 429326 214718 429562 214954
rect 429646 214718 429882 214954
rect 429326 214398 429562 214634
rect 429646 214398 429882 214634
rect 429326 178718 429562 178954
rect 429646 178718 429882 178954
rect 429326 178398 429562 178634
rect 429646 178398 429882 178634
rect 429326 142718 429562 142954
rect 429646 142718 429882 142954
rect 429326 142398 429562 142634
rect 429646 142398 429882 142634
rect 429326 106718 429562 106954
rect 429646 106718 429882 106954
rect 429326 106398 429562 106634
rect 429646 106398 429882 106634
rect 429326 70718 429562 70954
rect 429646 70718 429882 70954
rect 429326 70398 429562 70634
rect 429646 70398 429882 70634
rect 429326 34718 429562 34954
rect 429646 34718 429882 34954
rect 429326 34398 429562 34634
rect 429646 34398 429882 34634
rect 429326 -7302 429562 -7066
rect 429646 -7302 429882 -7066
rect 429326 -7622 429562 -7386
rect 429646 -7622 429882 -7386
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 438326 705562 438562 705798
rect 438646 705562 438882 705798
rect 438326 705242 438562 705478
rect 438646 705242 438882 705478
rect 438326 691718 438562 691954
rect 438646 691718 438882 691954
rect 438326 691398 438562 691634
rect 438646 691398 438882 691634
rect 438326 655718 438562 655954
rect 438646 655718 438882 655954
rect 438326 655398 438562 655634
rect 438646 655398 438882 655634
rect 438326 619718 438562 619954
rect 438646 619718 438882 619954
rect 438326 619398 438562 619634
rect 438646 619398 438882 619634
rect 438326 583718 438562 583954
rect 438646 583718 438882 583954
rect 438326 583398 438562 583634
rect 438646 583398 438882 583634
rect 438326 547718 438562 547954
rect 438646 547718 438882 547954
rect 438326 547398 438562 547634
rect 438646 547398 438882 547634
rect 438326 511718 438562 511954
rect 438646 511718 438882 511954
rect 438326 511398 438562 511634
rect 438646 511398 438882 511634
rect 438326 475718 438562 475954
rect 438646 475718 438882 475954
rect 438326 475398 438562 475634
rect 438646 475398 438882 475634
rect 438326 439718 438562 439954
rect 438646 439718 438882 439954
rect 438326 439398 438562 439634
rect 438646 439398 438882 439634
rect 438326 403718 438562 403954
rect 438646 403718 438882 403954
rect 438326 403398 438562 403634
rect 438646 403398 438882 403634
rect 438326 367718 438562 367954
rect 438646 367718 438882 367954
rect 438326 367398 438562 367634
rect 438646 367398 438882 367634
rect 438326 331718 438562 331954
rect 438646 331718 438882 331954
rect 438326 331398 438562 331634
rect 438646 331398 438882 331634
rect 438326 295718 438562 295954
rect 438646 295718 438882 295954
rect 438326 295398 438562 295634
rect 438646 295398 438882 295634
rect 438326 259718 438562 259954
rect 438646 259718 438882 259954
rect 438326 259398 438562 259634
rect 438646 259398 438882 259634
rect 438326 223718 438562 223954
rect 438646 223718 438882 223954
rect 438326 223398 438562 223634
rect 438646 223398 438882 223634
rect 438326 187718 438562 187954
rect 438646 187718 438882 187954
rect 438326 187398 438562 187634
rect 438646 187398 438882 187634
rect 438326 151718 438562 151954
rect 438646 151718 438882 151954
rect 438326 151398 438562 151634
rect 438646 151398 438882 151634
rect 438326 115718 438562 115954
rect 438646 115718 438882 115954
rect 438326 115398 438562 115634
rect 438646 115398 438882 115634
rect 438326 79718 438562 79954
rect 438646 79718 438882 79954
rect 438326 79398 438562 79634
rect 438646 79398 438882 79634
rect 438326 43718 438562 43954
rect 438646 43718 438882 43954
rect 438326 43398 438562 43634
rect 438646 43398 438882 43634
rect 438326 7718 438562 7954
rect 438646 7718 438882 7954
rect 438326 7398 438562 7634
rect 438646 7398 438882 7634
rect 438326 -1542 438562 -1306
rect 438646 -1542 438882 -1306
rect 438326 -1862 438562 -1626
rect 438646 -1862 438882 -1626
rect 442826 706522 443062 706758
rect 443146 706522 443382 706758
rect 442826 706202 443062 706438
rect 443146 706202 443382 706438
rect 442826 696218 443062 696454
rect 443146 696218 443382 696454
rect 442826 695898 443062 696134
rect 443146 695898 443382 696134
rect 442826 660218 443062 660454
rect 443146 660218 443382 660454
rect 442826 659898 443062 660134
rect 443146 659898 443382 660134
rect 442826 624218 443062 624454
rect 443146 624218 443382 624454
rect 442826 623898 443062 624134
rect 443146 623898 443382 624134
rect 442826 588218 443062 588454
rect 443146 588218 443382 588454
rect 442826 587898 443062 588134
rect 443146 587898 443382 588134
rect 442826 552218 443062 552454
rect 443146 552218 443382 552454
rect 442826 551898 443062 552134
rect 443146 551898 443382 552134
rect 442826 516218 443062 516454
rect 443146 516218 443382 516454
rect 442826 515898 443062 516134
rect 443146 515898 443382 516134
rect 442826 480218 443062 480454
rect 443146 480218 443382 480454
rect 442826 479898 443062 480134
rect 443146 479898 443382 480134
rect 442826 444218 443062 444454
rect 443146 444218 443382 444454
rect 442826 443898 443062 444134
rect 443146 443898 443382 444134
rect 442826 408218 443062 408454
rect 443146 408218 443382 408454
rect 442826 407898 443062 408134
rect 443146 407898 443382 408134
rect 442826 372218 443062 372454
rect 443146 372218 443382 372454
rect 442826 371898 443062 372134
rect 443146 371898 443382 372134
rect 442826 336218 443062 336454
rect 443146 336218 443382 336454
rect 442826 335898 443062 336134
rect 443146 335898 443382 336134
rect 442826 300218 443062 300454
rect 443146 300218 443382 300454
rect 442826 299898 443062 300134
rect 443146 299898 443382 300134
rect 442826 264218 443062 264454
rect 443146 264218 443382 264454
rect 442826 263898 443062 264134
rect 443146 263898 443382 264134
rect 442826 228218 443062 228454
rect 443146 228218 443382 228454
rect 442826 227898 443062 228134
rect 443146 227898 443382 228134
rect 442826 192218 443062 192454
rect 443146 192218 443382 192454
rect 442826 191898 443062 192134
rect 443146 191898 443382 192134
rect 442826 156218 443062 156454
rect 443146 156218 443382 156454
rect 442826 155898 443062 156134
rect 443146 155898 443382 156134
rect 442826 120218 443062 120454
rect 443146 120218 443382 120454
rect 442826 119898 443062 120134
rect 443146 119898 443382 120134
rect 442826 84218 443062 84454
rect 443146 84218 443382 84454
rect 442826 83898 443062 84134
rect 443146 83898 443382 84134
rect 442826 48218 443062 48454
rect 443146 48218 443382 48454
rect 442826 47898 443062 48134
rect 443146 47898 443382 48134
rect 442826 12218 443062 12454
rect 443146 12218 443382 12454
rect 442826 11898 443062 12134
rect 443146 11898 443382 12134
rect 442826 -2502 443062 -2266
rect 443146 -2502 443382 -2266
rect 442826 -2822 443062 -2586
rect 443146 -2822 443382 -2586
rect 447326 707482 447562 707718
rect 447646 707482 447882 707718
rect 447326 707162 447562 707398
rect 447646 707162 447882 707398
rect 447326 700718 447562 700954
rect 447646 700718 447882 700954
rect 447326 700398 447562 700634
rect 447646 700398 447882 700634
rect 447326 664718 447562 664954
rect 447646 664718 447882 664954
rect 447326 664398 447562 664634
rect 447646 664398 447882 664634
rect 447326 628718 447562 628954
rect 447646 628718 447882 628954
rect 447326 628398 447562 628634
rect 447646 628398 447882 628634
rect 447326 592718 447562 592954
rect 447646 592718 447882 592954
rect 447326 592398 447562 592634
rect 447646 592398 447882 592634
rect 447326 556718 447562 556954
rect 447646 556718 447882 556954
rect 447326 556398 447562 556634
rect 447646 556398 447882 556634
rect 447326 520718 447562 520954
rect 447646 520718 447882 520954
rect 447326 520398 447562 520634
rect 447646 520398 447882 520634
rect 447326 484718 447562 484954
rect 447646 484718 447882 484954
rect 447326 484398 447562 484634
rect 447646 484398 447882 484634
rect 447326 448718 447562 448954
rect 447646 448718 447882 448954
rect 447326 448398 447562 448634
rect 447646 448398 447882 448634
rect 447326 412718 447562 412954
rect 447646 412718 447882 412954
rect 447326 412398 447562 412634
rect 447646 412398 447882 412634
rect 447326 376718 447562 376954
rect 447646 376718 447882 376954
rect 447326 376398 447562 376634
rect 447646 376398 447882 376634
rect 447326 340718 447562 340954
rect 447646 340718 447882 340954
rect 447326 340398 447562 340634
rect 447646 340398 447882 340634
rect 447326 304718 447562 304954
rect 447646 304718 447882 304954
rect 447326 304398 447562 304634
rect 447646 304398 447882 304634
rect 447326 268718 447562 268954
rect 447646 268718 447882 268954
rect 447326 268398 447562 268634
rect 447646 268398 447882 268634
rect 447326 232718 447562 232954
rect 447646 232718 447882 232954
rect 447326 232398 447562 232634
rect 447646 232398 447882 232634
rect 447326 196718 447562 196954
rect 447646 196718 447882 196954
rect 447326 196398 447562 196634
rect 447646 196398 447882 196634
rect 447326 160718 447562 160954
rect 447646 160718 447882 160954
rect 447326 160398 447562 160634
rect 447646 160398 447882 160634
rect 447326 124718 447562 124954
rect 447646 124718 447882 124954
rect 447326 124398 447562 124634
rect 447646 124398 447882 124634
rect 447326 88718 447562 88954
rect 447646 88718 447882 88954
rect 447326 88398 447562 88634
rect 447646 88398 447882 88634
rect 447326 52718 447562 52954
rect 447646 52718 447882 52954
rect 447326 52398 447562 52634
rect 447646 52398 447882 52634
rect 447326 16718 447562 16954
rect 447646 16718 447882 16954
rect 447326 16398 447562 16634
rect 447646 16398 447882 16634
rect 447326 -3462 447562 -3226
rect 447646 -3462 447882 -3226
rect 447326 -3782 447562 -3546
rect 447646 -3782 447882 -3546
rect 451826 708442 452062 708678
rect 452146 708442 452382 708678
rect 451826 708122 452062 708358
rect 452146 708122 452382 708358
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -4422 452062 -4186
rect 452146 -4422 452382 -4186
rect 451826 -4742 452062 -4506
rect 452146 -4742 452382 -4506
rect 456326 709402 456562 709638
rect 456646 709402 456882 709638
rect 456326 709082 456562 709318
rect 456646 709082 456882 709318
rect 456326 673718 456562 673954
rect 456646 673718 456882 673954
rect 456326 673398 456562 673634
rect 456646 673398 456882 673634
rect 456326 637718 456562 637954
rect 456646 637718 456882 637954
rect 456326 637398 456562 637634
rect 456646 637398 456882 637634
rect 456326 601718 456562 601954
rect 456646 601718 456882 601954
rect 456326 601398 456562 601634
rect 456646 601398 456882 601634
rect 456326 565718 456562 565954
rect 456646 565718 456882 565954
rect 456326 565398 456562 565634
rect 456646 565398 456882 565634
rect 456326 529718 456562 529954
rect 456646 529718 456882 529954
rect 456326 529398 456562 529634
rect 456646 529398 456882 529634
rect 456326 493718 456562 493954
rect 456646 493718 456882 493954
rect 456326 493398 456562 493634
rect 456646 493398 456882 493634
rect 456326 457718 456562 457954
rect 456646 457718 456882 457954
rect 456326 457398 456562 457634
rect 456646 457398 456882 457634
rect 456326 421718 456562 421954
rect 456646 421718 456882 421954
rect 456326 421398 456562 421634
rect 456646 421398 456882 421634
rect 456326 385718 456562 385954
rect 456646 385718 456882 385954
rect 456326 385398 456562 385634
rect 456646 385398 456882 385634
rect 456326 349718 456562 349954
rect 456646 349718 456882 349954
rect 456326 349398 456562 349634
rect 456646 349398 456882 349634
rect 456326 313718 456562 313954
rect 456646 313718 456882 313954
rect 456326 313398 456562 313634
rect 456646 313398 456882 313634
rect 456326 277718 456562 277954
rect 456646 277718 456882 277954
rect 456326 277398 456562 277634
rect 456646 277398 456882 277634
rect 456326 241718 456562 241954
rect 456646 241718 456882 241954
rect 456326 241398 456562 241634
rect 456646 241398 456882 241634
rect 456326 205718 456562 205954
rect 456646 205718 456882 205954
rect 456326 205398 456562 205634
rect 456646 205398 456882 205634
rect 456326 169718 456562 169954
rect 456646 169718 456882 169954
rect 456326 169398 456562 169634
rect 456646 169398 456882 169634
rect 456326 133718 456562 133954
rect 456646 133718 456882 133954
rect 456326 133398 456562 133634
rect 456646 133398 456882 133634
rect 456326 97718 456562 97954
rect 456646 97718 456882 97954
rect 456326 97398 456562 97634
rect 456646 97398 456882 97634
rect 456326 61718 456562 61954
rect 456646 61718 456882 61954
rect 456326 61398 456562 61634
rect 456646 61398 456882 61634
rect 456326 25718 456562 25954
rect 456646 25718 456882 25954
rect 456326 25398 456562 25634
rect 456646 25398 456882 25634
rect 456326 -5382 456562 -5146
rect 456646 -5382 456882 -5146
rect 456326 -5702 456562 -5466
rect 456646 -5702 456882 -5466
rect 460826 710362 461062 710598
rect 461146 710362 461382 710598
rect 460826 710042 461062 710278
rect 461146 710042 461382 710278
rect 460826 678218 461062 678454
rect 461146 678218 461382 678454
rect 460826 677898 461062 678134
rect 461146 677898 461382 678134
rect 460826 642218 461062 642454
rect 461146 642218 461382 642454
rect 460826 641898 461062 642134
rect 461146 641898 461382 642134
rect 460826 606218 461062 606454
rect 461146 606218 461382 606454
rect 460826 605898 461062 606134
rect 461146 605898 461382 606134
rect 460826 570218 461062 570454
rect 461146 570218 461382 570454
rect 460826 569898 461062 570134
rect 461146 569898 461382 570134
rect 460826 534218 461062 534454
rect 461146 534218 461382 534454
rect 460826 533898 461062 534134
rect 461146 533898 461382 534134
rect 460826 498218 461062 498454
rect 461146 498218 461382 498454
rect 460826 497898 461062 498134
rect 461146 497898 461382 498134
rect 460826 462218 461062 462454
rect 461146 462218 461382 462454
rect 460826 461898 461062 462134
rect 461146 461898 461382 462134
rect 460826 426218 461062 426454
rect 461146 426218 461382 426454
rect 460826 425898 461062 426134
rect 461146 425898 461382 426134
rect 460826 390218 461062 390454
rect 461146 390218 461382 390454
rect 460826 389898 461062 390134
rect 461146 389898 461382 390134
rect 460826 354218 461062 354454
rect 461146 354218 461382 354454
rect 460826 353898 461062 354134
rect 461146 353898 461382 354134
rect 460826 318218 461062 318454
rect 461146 318218 461382 318454
rect 460826 317898 461062 318134
rect 461146 317898 461382 318134
rect 460826 282218 461062 282454
rect 461146 282218 461382 282454
rect 460826 281898 461062 282134
rect 461146 281898 461382 282134
rect 460826 246218 461062 246454
rect 461146 246218 461382 246454
rect 460826 245898 461062 246134
rect 461146 245898 461382 246134
rect 460826 210218 461062 210454
rect 461146 210218 461382 210454
rect 460826 209898 461062 210134
rect 461146 209898 461382 210134
rect 460826 174218 461062 174454
rect 461146 174218 461382 174454
rect 460826 173898 461062 174134
rect 461146 173898 461382 174134
rect 460826 138218 461062 138454
rect 461146 138218 461382 138454
rect 460826 137898 461062 138134
rect 461146 137898 461382 138134
rect 460826 102218 461062 102454
rect 461146 102218 461382 102454
rect 460826 101898 461062 102134
rect 461146 101898 461382 102134
rect 460826 66218 461062 66454
rect 461146 66218 461382 66454
rect 460826 65898 461062 66134
rect 461146 65898 461382 66134
rect 460826 30218 461062 30454
rect 461146 30218 461382 30454
rect 460826 29898 461062 30134
rect 461146 29898 461382 30134
rect 460826 -6342 461062 -6106
rect 461146 -6342 461382 -6106
rect 460826 -6662 461062 -6426
rect 461146 -6662 461382 -6426
rect 465326 711322 465562 711558
rect 465646 711322 465882 711558
rect 465326 711002 465562 711238
rect 465646 711002 465882 711238
rect 465326 682718 465562 682954
rect 465646 682718 465882 682954
rect 465326 682398 465562 682634
rect 465646 682398 465882 682634
rect 465326 646718 465562 646954
rect 465646 646718 465882 646954
rect 465326 646398 465562 646634
rect 465646 646398 465882 646634
rect 465326 610718 465562 610954
rect 465646 610718 465882 610954
rect 465326 610398 465562 610634
rect 465646 610398 465882 610634
rect 465326 574718 465562 574954
rect 465646 574718 465882 574954
rect 465326 574398 465562 574634
rect 465646 574398 465882 574634
rect 465326 538718 465562 538954
rect 465646 538718 465882 538954
rect 465326 538398 465562 538634
rect 465646 538398 465882 538634
rect 465326 502718 465562 502954
rect 465646 502718 465882 502954
rect 465326 502398 465562 502634
rect 465646 502398 465882 502634
rect 465326 466718 465562 466954
rect 465646 466718 465882 466954
rect 465326 466398 465562 466634
rect 465646 466398 465882 466634
rect 465326 430718 465562 430954
rect 465646 430718 465882 430954
rect 465326 430398 465562 430634
rect 465646 430398 465882 430634
rect 465326 394718 465562 394954
rect 465646 394718 465882 394954
rect 465326 394398 465562 394634
rect 465646 394398 465882 394634
rect 465326 358718 465562 358954
rect 465646 358718 465882 358954
rect 465326 358398 465562 358634
rect 465646 358398 465882 358634
rect 465326 322718 465562 322954
rect 465646 322718 465882 322954
rect 465326 322398 465562 322634
rect 465646 322398 465882 322634
rect 465326 286718 465562 286954
rect 465646 286718 465882 286954
rect 465326 286398 465562 286634
rect 465646 286398 465882 286634
rect 465326 250718 465562 250954
rect 465646 250718 465882 250954
rect 465326 250398 465562 250634
rect 465646 250398 465882 250634
rect 465326 214718 465562 214954
rect 465646 214718 465882 214954
rect 465326 214398 465562 214634
rect 465646 214398 465882 214634
rect 465326 178718 465562 178954
rect 465646 178718 465882 178954
rect 465326 178398 465562 178634
rect 465646 178398 465882 178634
rect 465326 142718 465562 142954
rect 465646 142718 465882 142954
rect 465326 142398 465562 142634
rect 465646 142398 465882 142634
rect 465326 106718 465562 106954
rect 465646 106718 465882 106954
rect 465326 106398 465562 106634
rect 465646 106398 465882 106634
rect 465326 70718 465562 70954
rect 465646 70718 465882 70954
rect 465326 70398 465562 70634
rect 465646 70398 465882 70634
rect 465326 34718 465562 34954
rect 465646 34718 465882 34954
rect 465326 34398 465562 34634
rect 465646 34398 465882 34634
rect 465326 -7302 465562 -7066
rect 465646 -7302 465882 -7066
rect 465326 -7622 465562 -7386
rect 465646 -7622 465882 -7386
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 474326 705562 474562 705798
rect 474646 705562 474882 705798
rect 474326 705242 474562 705478
rect 474646 705242 474882 705478
rect 474326 691718 474562 691954
rect 474646 691718 474882 691954
rect 474326 691398 474562 691634
rect 474646 691398 474882 691634
rect 474326 655718 474562 655954
rect 474646 655718 474882 655954
rect 474326 655398 474562 655634
rect 474646 655398 474882 655634
rect 474326 619718 474562 619954
rect 474646 619718 474882 619954
rect 474326 619398 474562 619634
rect 474646 619398 474882 619634
rect 474326 583718 474562 583954
rect 474646 583718 474882 583954
rect 474326 583398 474562 583634
rect 474646 583398 474882 583634
rect 474326 547718 474562 547954
rect 474646 547718 474882 547954
rect 474326 547398 474562 547634
rect 474646 547398 474882 547634
rect 474326 511718 474562 511954
rect 474646 511718 474882 511954
rect 474326 511398 474562 511634
rect 474646 511398 474882 511634
rect 474326 475718 474562 475954
rect 474646 475718 474882 475954
rect 474326 475398 474562 475634
rect 474646 475398 474882 475634
rect 474326 439718 474562 439954
rect 474646 439718 474882 439954
rect 474326 439398 474562 439634
rect 474646 439398 474882 439634
rect 474326 403718 474562 403954
rect 474646 403718 474882 403954
rect 474326 403398 474562 403634
rect 474646 403398 474882 403634
rect 474326 367718 474562 367954
rect 474646 367718 474882 367954
rect 474326 367398 474562 367634
rect 474646 367398 474882 367634
rect 474326 331718 474562 331954
rect 474646 331718 474882 331954
rect 474326 331398 474562 331634
rect 474646 331398 474882 331634
rect 474326 295718 474562 295954
rect 474646 295718 474882 295954
rect 474326 295398 474562 295634
rect 474646 295398 474882 295634
rect 474326 259718 474562 259954
rect 474646 259718 474882 259954
rect 474326 259398 474562 259634
rect 474646 259398 474882 259634
rect 474326 223718 474562 223954
rect 474646 223718 474882 223954
rect 474326 223398 474562 223634
rect 474646 223398 474882 223634
rect 474326 187718 474562 187954
rect 474646 187718 474882 187954
rect 474326 187398 474562 187634
rect 474646 187398 474882 187634
rect 474326 151718 474562 151954
rect 474646 151718 474882 151954
rect 474326 151398 474562 151634
rect 474646 151398 474882 151634
rect 474326 115718 474562 115954
rect 474646 115718 474882 115954
rect 474326 115398 474562 115634
rect 474646 115398 474882 115634
rect 474326 79718 474562 79954
rect 474646 79718 474882 79954
rect 474326 79398 474562 79634
rect 474646 79398 474882 79634
rect 474326 43718 474562 43954
rect 474646 43718 474882 43954
rect 474326 43398 474562 43634
rect 474646 43398 474882 43634
rect 474326 7718 474562 7954
rect 474646 7718 474882 7954
rect 474326 7398 474562 7634
rect 474646 7398 474882 7634
rect 474326 -1542 474562 -1306
rect 474646 -1542 474882 -1306
rect 474326 -1862 474562 -1626
rect 474646 -1862 474882 -1626
rect 478826 706522 479062 706758
rect 479146 706522 479382 706758
rect 478826 706202 479062 706438
rect 479146 706202 479382 706438
rect 478826 696218 479062 696454
rect 479146 696218 479382 696454
rect 478826 695898 479062 696134
rect 479146 695898 479382 696134
rect 478826 660218 479062 660454
rect 479146 660218 479382 660454
rect 478826 659898 479062 660134
rect 479146 659898 479382 660134
rect 478826 624218 479062 624454
rect 479146 624218 479382 624454
rect 478826 623898 479062 624134
rect 479146 623898 479382 624134
rect 478826 588218 479062 588454
rect 479146 588218 479382 588454
rect 478826 587898 479062 588134
rect 479146 587898 479382 588134
rect 478826 552218 479062 552454
rect 479146 552218 479382 552454
rect 478826 551898 479062 552134
rect 479146 551898 479382 552134
rect 478826 516218 479062 516454
rect 479146 516218 479382 516454
rect 478826 515898 479062 516134
rect 479146 515898 479382 516134
rect 478826 480218 479062 480454
rect 479146 480218 479382 480454
rect 478826 479898 479062 480134
rect 479146 479898 479382 480134
rect 478826 444218 479062 444454
rect 479146 444218 479382 444454
rect 478826 443898 479062 444134
rect 479146 443898 479382 444134
rect 478826 408218 479062 408454
rect 479146 408218 479382 408454
rect 478826 407898 479062 408134
rect 479146 407898 479382 408134
rect 478826 372218 479062 372454
rect 479146 372218 479382 372454
rect 478826 371898 479062 372134
rect 479146 371898 479382 372134
rect 478826 336218 479062 336454
rect 479146 336218 479382 336454
rect 478826 335898 479062 336134
rect 479146 335898 479382 336134
rect 478826 300218 479062 300454
rect 479146 300218 479382 300454
rect 478826 299898 479062 300134
rect 479146 299898 479382 300134
rect 478826 264218 479062 264454
rect 479146 264218 479382 264454
rect 478826 263898 479062 264134
rect 479146 263898 479382 264134
rect 478826 228218 479062 228454
rect 479146 228218 479382 228454
rect 478826 227898 479062 228134
rect 479146 227898 479382 228134
rect 478826 192218 479062 192454
rect 479146 192218 479382 192454
rect 478826 191898 479062 192134
rect 479146 191898 479382 192134
rect 478826 156218 479062 156454
rect 479146 156218 479382 156454
rect 478826 155898 479062 156134
rect 479146 155898 479382 156134
rect 478826 120218 479062 120454
rect 479146 120218 479382 120454
rect 478826 119898 479062 120134
rect 479146 119898 479382 120134
rect 478826 84218 479062 84454
rect 479146 84218 479382 84454
rect 478826 83898 479062 84134
rect 479146 83898 479382 84134
rect 478826 48218 479062 48454
rect 479146 48218 479382 48454
rect 478826 47898 479062 48134
rect 479146 47898 479382 48134
rect 478826 12218 479062 12454
rect 479146 12218 479382 12454
rect 478826 11898 479062 12134
rect 479146 11898 479382 12134
rect 478826 -2502 479062 -2266
rect 479146 -2502 479382 -2266
rect 478826 -2822 479062 -2586
rect 479146 -2822 479382 -2586
rect 483326 707482 483562 707718
rect 483646 707482 483882 707718
rect 483326 707162 483562 707398
rect 483646 707162 483882 707398
rect 483326 700718 483562 700954
rect 483646 700718 483882 700954
rect 483326 700398 483562 700634
rect 483646 700398 483882 700634
rect 483326 664718 483562 664954
rect 483646 664718 483882 664954
rect 483326 664398 483562 664634
rect 483646 664398 483882 664634
rect 483326 628718 483562 628954
rect 483646 628718 483882 628954
rect 483326 628398 483562 628634
rect 483646 628398 483882 628634
rect 483326 592718 483562 592954
rect 483646 592718 483882 592954
rect 483326 592398 483562 592634
rect 483646 592398 483882 592634
rect 483326 556718 483562 556954
rect 483646 556718 483882 556954
rect 483326 556398 483562 556634
rect 483646 556398 483882 556634
rect 483326 520718 483562 520954
rect 483646 520718 483882 520954
rect 483326 520398 483562 520634
rect 483646 520398 483882 520634
rect 483326 484718 483562 484954
rect 483646 484718 483882 484954
rect 483326 484398 483562 484634
rect 483646 484398 483882 484634
rect 483326 448718 483562 448954
rect 483646 448718 483882 448954
rect 483326 448398 483562 448634
rect 483646 448398 483882 448634
rect 483326 412718 483562 412954
rect 483646 412718 483882 412954
rect 483326 412398 483562 412634
rect 483646 412398 483882 412634
rect 483326 376718 483562 376954
rect 483646 376718 483882 376954
rect 483326 376398 483562 376634
rect 483646 376398 483882 376634
rect 483326 340718 483562 340954
rect 483646 340718 483882 340954
rect 483326 340398 483562 340634
rect 483646 340398 483882 340634
rect 483326 304718 483562 304954
rect 483646 304718 483882 304954
rect 483326 304398 483562 304634
rect 483646 304398 483882 304634
rect 483326 268718 483562 268954
rect 483646 268718 483882 268954
rect 483326 268398 483562 268634
rect 483646 268398 483882 268634
rect 483326 232718 483562 232954
rect 483646 232718 483882 232954
rect 483326 232398 483562 232634
rect 483646 232398 483882 232634
rect 483326 196718 483562 196954
rect 483646 196718 483882 196954
rect 483326 196398 483562 196634
rect 483646 196398 483882 196634
rect 483326 160718 483562 160954
rect 483646 160718 483882 160954
rect 483326 160398 483562 160634
rect 483646 160398 483882 160634
rect 483326 124718 483562 124954
rect 483646 124718 483882 124954
rect 483326 124398 483562 124634
rect 483646 124398 483882 124634
rect 483326 88718 483562 88954
rect 483646 88718 483882 88954
rect 483326 88398 483562 88634
rect 483646 88398 483882 88634
rect 483326 52718 483562 52954
rect 483646 52718 483882 52954
rect 483326 52398 483562 52634
rect 483646 52398 483882 52634
rect 483326 16718 483562 16954
rect 483646 16718 483882 16954
rect 483326 16398 483562 16634
rect 483646 16398 483882 16634
rect 483326 -3462 483562 -3226
rect 483646 -3462 483882 -3226
rect 483326 -3782 483562 -3546
rect 483646 -3782 483882 -3546
rect 487826 708442 488062 708678
rect 488146 708442 488382 708678
rect 487826 708122 488062 708358
rect 488146 708122 488382 708358
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -4422 488062 -4186
rect 488146 -4422 488382 -4186
rect 487826 -4742 488062 -4506
rect 488146 -4742 488382 -4506
rect 492326 709402 492562 709638
rect 492646 709402 492882 709638
rect 492326 709082 492562 709318
rect 492646 709082 492882 709318
rect 492326 673718 492562 673954
rect 492646 673718 492882 673954
rect 492326 673398 492562 673634
rect 492646 673398 492882 673634
rect 492326 637718 492562 637954
rect 492646 637718 492882 637954
rect 492326 637398 492562 637634
rect 492646 637398 492882 637634
rect 492326 601718 492562 601954
rect 492646 601718 492882 601954
rect 492326 601398 492562 601634
rect 492646 601398 492882 601634
rect 492326 565718 492562 565954
rect 492646 565718 492882 565954
rect 492326 565398 492562 565634
rect 492646 565398 492882 565634
rect 492326 529718 492562 529954
rect 492646 529718 492882 529954
rect 492326 529398 492562 529634
rect 492646 529398 492882 529634
rect 492326 493718 492562 493954
rect 492646 493718 492882 493954
rect 492326 493398 492562 493634
rect 492646 493398 492882 493634
rect 492326 457718 492562 457954
rect 492646 457718 492882 457954
rect 492326 457398 492562 457634
rect 492646 457398 492882 457634
rect 492326 421718 492562 421954
rect 492646 421718 492882 421954
rect 492326 421398 492562 421634
rect 492646 421398 492882 421634
rect 492326 385718 492562 385954
rect 492646 385718 492882 385954
rect 492326 385398 492562 385634
rect 492646 385398 492882 385634
rect 492326 349718 492562 349954
rect 492646 349718 492882 349954
rect 492326 349398 492562 349634
rect 492646 349398 492882 349634
rect 492326 313718 492562 313954
rect 492646 313718 492882 313954
rect 492326 313398 492562 313634
rect 492646 313398 492882 313634
rect 492326 277718 492562 277954
rect 492646 277718 492882 277954
rect 492326 277398 492562 277634
rect 492646 277398 492882 277634
rect 492326 241718 492562 241954
rect 492646 241718 492882 241954
rect 492326 241398 492562 241634
rect 492646 241398 492882 241634
rect 492326 205718 492562 205954
rect 492646 205718 492882 205954
rect 492326 205398 492562 205634
rect 492646 205398 492882 205634
rect 492326 169718 492562 169954
rect 492646 169718 492882 169954
rect 492326 169398 492562 169634
rect 492646 169398 492882 169634
rect 492326 133718 492562 133954
rect 492646 133718 492882 133954
rect 492326 133398 492562 133634
rect 492646 133398 492882 133634
rect 492326 97718 492562 97954
rect 492646 97718 492882 97954
rect 492326 97398 492562 97634
rect 492646 97398 492882 97634
rect 492326 61718 492562 61954
rect 492646 61718 492882 61954
rect 492326 61398 492562 61634
rect 492646 61398 492882 61634
rect 492326 25718 492562 25954
rect 492646 25718 492882 25954
rect 492326 25398 492562 25634
rect 492646 25398 492882 25634
rect 492326 -5382 492562 -5146
rect 492646 -5382 492882 -5146
rect 492326 -5702 492562 -5466
rect 492646 -5702 492882 -5466
rect 496826 710362 497062 710598
rect 497146 710362 497382 710598
rect 496826 710042 497062 710278
rect 497146 710042 497382 710278
rect 496826 678218 497062 678454
rect 497146 678218 497382 678454
rect 496826 677898 497062 678134
rect 497146 677898 497382 678134
rect 496826 642218 497062 642454
rect 497146 642218 497382 642454
rect 496826 641898 497062 642134
rect 497146 641898 497382 642134
rect 496826 606218 497062 606454
rect 497146 606218 497382 606454
rect 496826 605898 497062 606134
rect 497146 605898 497382 606134
rect 496826 570218 497062 570454
rect 497146 570218 497382 570454
rect 496826 569898 497062 570134
rect 497146 569898 497382 570134
rect 496826 534218 497062 534454
rect 497146 534218 497382 534454
rect 496826 533898 497062 534134
rect 497146 533898 497382 534134
rect 496826 498218 497062 498454
rect 497146 498218 497382 498454
rect 496826 497898 497062 498134
rect 497146 497898 497382 498134
rect 496826 462218 497062 462454
rect 497146 462218 497382 462454
rect 496826 461898 497062 462134
rect 497146 461898 497382 462134
rect 496826 426218 497062 426454
rect 497146 426218 497382 426454
rect 496826 425898 497062 426134
rect 497146 425898 497382 426134
rect 496826 390218 497062 390454
rect 497146 390218 497382 390454
rect 496826 389898 497062 390134
rect 497146 389898 497382 390134
rect 496826 354218 497062 354454
rect 497146 354218 497382 354454
rect 496826 353898 497062 354134
rect 497146 353898 497382 354134
rect 496826 318218 497062 318454
rect 497146 318218 497382 318454
rect 496826 317898 497062 318134
rect 497146 317898 497382 318134
rect 496826 282218 497062 282454
rect 497146 282218 497382 282454
rect 496826 281898 497062 282134
rect 497146 281898 497382 282134
rect 496826 246218 497062 246454
rect 497146 246218 497382 246454
rect 496826 245898 497062 246134
rect 497146 245898 497382 246134
rect 496826 210218 497062 210454
rect 497146 210218 497382 210454
rect 496826 209898 497062 210134
rect 497146 209898 497382 210134
rect 496826 174218 497062 174454
rect 497146 174218 497382 174454
rect 496826 173898 497062 174134
rect 497146 173898 497382 174134
rect 496826 138218 497062 138454
rect 497146 138218 497382 138454
rect 496826 137898 497062 138134
rect 497146 137898 497382 138134
rect 496826 102218 497062 102454
rect 497146 102218 497382 102454
rect 496826 101898 497062 102134
rect 497146 101898 497382 102134
rect 496826 66218 497062 66454
rect 497146 66218 497382 66454
rect 496826 65898 497062 66134
rect 497146 65898 497382 66134
rect 496826 30218 497062 30454
rect 497146 30218 497382 30454
rect 496826 29898 497062 30134
rect 497146 29898 497382 30134
rect 496826 -6342 497062 -6106
rect 497146 -6342 497382 -6106
rect 496826 -6662 497062 -6426
rect 497146 -6662 497382 -6426
rect 501326 711322 501562 711558
rect 501646 711322 501882 711558
rect 501326 711002 501562 711238
rect 501646 711002 501882 711238
rect 501326 682718 501562 682954
rect 501646 682718 501882 682954
rect 501326 682398 501562 682634
rect 501646 682398 501882 682634
rect 501326 646718 501562 646954
rect 501646 646718 501882 646954
rect 501326 646398 501562 646634
rect 501646 646398 501882 646634
rect 501326 610718 501562 610954
rect 501646 610718 501882 610954
rect 501326 610398 501562 610634
rect 501646 610398 501882 610634
rect 501326 574718 501562 574954
rect 501646 574718 501882 574954
rect 501326 574398 501562 574634
rect 501646 574398 501882 574634
rect 501326 538718 501562 538954
rect 501646 538718 501882 538954
rect 501326 538398 501562 538634
rect 501646 538398 501882 538634
rect 501326 502718 501562 502954
rect 501646 502718 501882 502954
rect 501326 502398 501562 502634
rect 501646 502398 501882 502634
rect 501326 466718 501562 466954
rect 501646 466718 501882 466954
rect 501326 466398 501562 466634
rect 501646 466398 501882 466634
rect 501326 430718 501562 430954
rect 501646 430718 501882 430954
rect 501326 430398 501562 430634
rect 501646 430398 501882 430634
rect 501326 394718 501562 394954
rect 501646 394718 501882 394954
rect 501326 394398 501562 394634
rect 501646 394398 501882 394634
rect 501326 358718 501562 358954
rect 501646 358718 501882 358954
rect 501326 358398 501562 358634
rect 501646 358398 501882 358634
rect 501326 322718 501562 322954
rect 501646 322718 501882 322954
rect 501326 322398 501562 322634
rect 501646 322398 501882 322634
rect 501326 286718 501562 286954
rect 501646 286718 501882 286954
rect 501326 286398 501562 286634
rect 501646 286398 501882 286634
rect 501326 250718 501562 250954
rect 501646 250718 501882 250954
rect 501326 250398 501562 250634
rect 501646 250398 501882 250634
rect 501326 214718 501562 214954
rect 501646 214718 501882 214954
rect 501326 214398 501562 214634
rect 501646 214398 501882 214634
rect 501326 178718 501562 178954
rect 501646 178718 501882 178954
rect 501326 178398 501562 178634
rect 501646 178398 501882 178634
rect 501326 142718 501562 142954
rect 501646 142718 501882 142954
rect 501326 142398 501562 142634
rect 501646 142398 501882 142634
rect 501326 106718 501562 106954
rect 501646 106718 501882 106954
rect 501326 106398 501562 106634
rect 501646 106398 501882 106634
rect 501326 70718 501562 70954
rect 501646 70718 501882 70954
rect 501326 70398 501562 70634
rect 501646 70398 501882 70634
rect 501326 34718 501562 34954
rect 501646 34718 501882 34954
rect 501326 34398 501562 34634
rect 501646 34398 501882 34634
rect 501326 -7302 501562 -7066
rect 501646 -7302 501882 -7066
rect 501326 -7622 501562 -7386
rect 501646 -7622 501882 -7386
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 510326 705562 510562 705798
rect 510646 705562 510882 705798
rect 510326 705242 510562 705478
rect 510646 705242 510882 705478
rect 510326 691718 510562 691954
rect 510646 691718 510882 691954
rect 510326 691398 510562 691634
rect 510646 691398 510882 691634
rect 510326 655718 510562 655954
rect 510646 655718 510882 655954
rect 510326 655398 510562 655634
rect 510646 655398 510882 655634
rect 510326 619718 510562 619954
rect 510646 619718 510882 619954
rect 510326 619398 510562 619634
rect 510646 619398 510882 619634
rect 510326 583718 510562 583954
rect 510646 583718 510882 583954
rect 510326 583398 510562 583634
rect 510646 583398 510882 583634
rect 510326 547718 510562 547954
rect 510646 547718 510882 547954
rect 510326 547398 510562 547634
rect 510646 547398 510882 547634
rect 510326 511718 510562 511954
rect 510646 511718 510882 511954
rect 510326 511398 510562 511634
rect 510646 511398 510882 511634
rect 510326 475718 510562 475954
rect 510646 475718 510882 475954
rect 510326 475398 510562 475634
rect 510646 475398 510882 475634
rect 510326 439718 510562 439954
rect 510646 439718 510882 439954
rect 510326 439398 510562 439634
rect 510646 439398 510882 439634
rect 510326 403718 510562 403954
rect 510646 403718 510882 403954
rect 510326 403398 510562 403634
rect 510646 403398 510882 403634
rect 510326 367718 510562 367954
rect 510646 367718 510882 367954
rect 510326 367398 510562 367634
rect 510646 367398 510882 367634
rect 510326 331718 510562 331954
rect 510646 331718 510882 331954
rect 510326 331398 510562 331634
rect 510646 331398 510882 331634
rect 510326 295718 510562 295954
rect 510646 295718 510882 295954
rect 510326 295398 510562 295634
rect 510646 295398 510882 295634
rect 510326 259718 510562 259954
rect 510646 259718 510882 259954
rect 510326 259398 510562 259634
rect 510646 259398 510882 259634
rect 510326 223718 510562 223954
rect 510646 223718 510882 223954
rect 510326 223398 510562 223634
rect 510646 223398 510882 223634
rect 510326 187718 510562 187954
rect 510646 187718 510882 187954
rect 510326 187398 510562 187634
rect 510646 187398 510882 187634
rect 510326 151718 510562 151954
rect 510646 151718 510882 151954
rect 510326 151398 510562 151634
rect 510646 151398 510882 151634
rect 510326 115718 510562 115954
rect 510646 115718 510882 115954
rect 510326 115398 510562 115634
rect 510646 115398 510882 115634
rect 510326 79718 510562 79954
rect 510646 79718 510882 79954
rect 510326 79398 510562 79634
rect 510646 79398 510882 79634
rect 510326 43718 510562 43954
rect 510646 43718 510882 43954
rect 510326 43398 510562 43634
rect 510646 43398 510882 43634
rect 510326 7718 510562 7954
rect 510646 7718 510882 7954
rect 510326 7398 510562 7634
rect 510646 7398 510882 7634
rect 510326 -1542 510562 -1306
rect 510646 -1542 510882 -1306
rect 510326 -1862 510562 -1626
rect 510646 -1862 510882 -1626
rect 514826 706522 515062 706758
rect 515146 706522 515382 706758
rect 514826 706202 515062 706438
rect 515146 706202 515382 706438
rect 514826 696218 515062 696454
rect 515146 696218 515382 696454
rect 514826 695898 515062 696134
rect 515146 695898 515382 696134
rect 514826 660218 515062 660454
rect 515146 660218 515382 660454
rect 514826 659898 515062 660134
rect 515146 659898 515382 660134
rect 514826 624218 515062 624454
rect 515146 624218 515382 624454
rect 514826 623898 515062 624134
rect 515146 623898 515382 624134
rect 514826 588218 515062 588454
rect 515146 588218 515382 588454
rect 514826 587898 515062 588134
rect 515146 587898 515382 588134
rect 514826 552218 515062 552454
rect 515146 552218 515382 552454
rect 514826 551898 515062 552134
rect 515146 551898 515382 552134
rect 514826 516218 515062 516454
rect 515146 516218 515382 516454
rect 514826 515898 515062 516134
rect 515146 515898 515382 516134
rect 514826 480218 515062 480454
rect 515146 480218 515382 480454
rect 514826 479898 515062 480134
rect 515146 479898 515382 480134
rect 514826 444218 515062 444454
rect 515146 444218 515382 444454
rect 514826 443898 515062 444134
rect 515146 443898 515382 444134
rect 514826 408218 515062 408454
rect 515146 408218 515382 408454
rect 514826 407898 515062 408134
rect 515146 407898 515382 408134
rect 514826 372218 515062 372454
rect 515146 372218 515382 372454
rect 514826 371898 515062 372134
rect 515146 371898 515382 372134
rect 514826 336218 515062 336454
rect 515146 336218 515382 336454
rect 514826 335898 515062 336134
rect 515146 335898 515382 336134
rect 514826 300218 515062 300454
rect 515146 300218 515382 300454
rect 514826 299898 515062 300134
rect 515146 299898 515382 300134
rect 514826 264218 515062 264454
rect 515146 264218 515382 264454
rect 514826 263898 515062 264134
rect 515146 263898 515382 264134
rect 514826 228218 515062 228454
rect 515146 228218 515382 228454
rect 514826 227898 515062 228134
rect 515146 227898 515382 228134
rect 514826 192218 515062 192454
rect 515146 192218 515382 192454
rect 514826 191898 515062 192134
rect 515146 191898 515382 192134
rect 514826 156218 515062 156454
rect 515146 156218 515382 156454
rect 514826 155898 515062 156134
rect 515146 155898 515382 156134
rect 514826 120218 515062 120454
rect 515146 120218 515382 120454
rect 514826 119898 515062 120134
rect 515146 119898 515382 120134
rect 514826 84218 515062 84454
rect 515146 84218 515382 84454
rect 514826 83898 515062 84134
rect 515146 83898 515382 84134
rect 514826 48218 515062 48454
rect 515146 48218 515382 48454
rect 514826 47898 515062 48134
rect 515146 47898 515382 48134
rect 514826 12218 515062 12454
rect 515146 12218 515382 12454
rect 514826 11898 515062 12134
rect 515146 11898 515382 12134
rect 514826 -2502 515062 -2266
rect 515146 -2502 515382 -2266
rect 514826 -2822 515062 -2586
rect 515146 -2822 515382 -2586
rect 519326 707482 519562 707718
rect 519646 707482 519882 707718
rect 519326 707162 519562 707398
rect 519646 707162 519882 707398
rect 519326 700718 519562 700954
rect 519646 700718 519882 700954
rect 519326 700398 519562 700634
rect 519646 700398 519882 700634
rect 519326 664718 519562 664954
rect 519646 664718 519882 664954
rect 519326 664398 519562 664634
rect 519646 664398 519882 664634
rect 519326 628718 519562 628954
rect 519646 628718 519882 628954
rect 519326 628398 519562 628634
rect 519646 628398 519882 628634
rect 519326 592718 519562 592954
rect 519646 592718 519882 592954
rect 519326 592398 519562 592634
rect 519646 592398 519882 592634
rect 519326 556718 519562 556954
rect 519646 556718 519882 556954
rect 519326 556398 519562 556634
rect 519646 556398 519882 556634
rect 519326 520718 519562 520954
rect 519646 520718 519882 520954
rect 519326 520398 519562 520634
rect 519646 520398 519882 520634
rect 519326 484718 519562 484954
rect 519646 484718 519882 484954
rect 519326 484398 519562 484634
rect 519646 484398 519882 484634
rect 519326 448718 519562 448954
rect 519646 448718 519882 448954
rect 519326 448398 519562 448634
rect 519646 448398 519882 448634
rect 519326 412718 519562 412954
rect 519646 412718 519882 412954
rect 519326 412398 519562 412634
rect 519646 412398 519882 412634
rect 519326 376718 519562 376954
rect 519646 376718 519882 376954
rect 519326 376398 519562 376634
rect 519646 376398 519882 376634
rect 519326 340718 519562 340954
rect 519646 340718 519882 340954
rect 519326 340398 519562 340634
rect 519646 340398 519882 340634
rect 519326 304718 519562 304954
rect 519646 304718 519882 304954
rect 519326 304398 519562 304634
rect 519646 304398 519882 304634
rect 519326 268718 519562 268954
rect 519646 268718 519882 268954
rect 519326 268398 519562 268634
rect 519646 268398 519882 268634
rect 519326 232718 519562 232954
rect 519646 232718 519882 232954
rect 519326 232398 519562 232634
rect 519646 232398 519882 232634
rect 519326 196718 519562 196954
rect 519646 196718 519882 196954
rect 519326 196398 519562 196634
rect 519646 196398 519882 196634
rect 519326 160718 519562 160954
rect 519646 160718 519882 160954
rect 519326 160398 519562 160634
rect 519646 160398 519882 160634
rect 519326 124718 519562 124954
rect 519646 124718 519882 124954
rect 519326 124398 519562 124634
rect 519646 124398 519882 124634
rect 519326 88718 519562 88954
rect 519646 88718 519882 88954
rect 519326 88398 519562 88634
rect 519646 88398 519882 88634
rect 519326 52718 519562 52954
rect 519646 52718 519882 52954
rect 519326 52398 519562 52634
rect 519646 52398 519882 52634
rect 519326 16718 519562 16954
rect 519646 16718 519882 16954
rect 519326 16398 519562 16634
rect 519646 16398 519882 16634
rect 519326 -3462 519562 -3226
rect 519646 -3462 519882 -3226
rect 519326 -3782 519562 -3546
rect 519646 -3782 519882 -3546
rect 523826 708442 524062 708678
rect 524146 708442 524382 708678
rect 523826 708122 524062 708358
rect 524146 708122 524382 708358
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -4422 524062 -4186
rect 524146 -4422 524382 -4186
rect 523826 -4742 524062 -4506
rect 524146 -4742 524382 -4506
rect 528326 709402 528562 709638
rect 528646 709402 528882 709638
rect 528326 709082 528562 709318
rect 528646 709082 528882 709318
rect 528326 673718 528562 673954
rect 528646 673718 528882 673954
rect 528326 673398 528562 673634
rect 528646 673398 528882 673634
rect 528326 637718 528562 637954
rect 528646 637718 528882 637954
rect 528326 637398 528562 637634
rect 528646 637398 528882 637634
rect 528326 601718 528562 601954
rect 528646 601718 528882 601954
rect 528326 601398 528562 601634
rect 528646 601398 528882 601634
rect 528326 565718 528562 565954
rect 528646 565718 528882 565954
rect 528326 565398 528562 565634
rect 528646 565398 528882 565634
rect 528326 529718 528562 529954
rect 528646 529718 528882 529954
rect 528326 529398 528562 529634
rect 528646 529398 528882 529634
rect 528326 493718 528562 493954
rect 528646 493718 528882 493954
rect 528326 493398 528562 493634
rect 528646 493398 528882 493634
rect 528326 457718 528562 457954
rect 528646 457718 528882 457954
rect 528326 457398 528562 457634
rect 528646 457398 528882 457634
rect 528326 421718 528562 421954
rect 528646 421718 528882 421954
rect 528326 421398 528562 421634
rect 528646 421398 528882 421634
rect 528326 385718 528562 385954
rect 528646 385718 528882 385954
rect 528326 385398 528562 385634
rect 528646 385398 528882 385634
rect 528326 349718 528562 349954
rect 528646 349718 528882 349954
rect 528326 349398 528562 349634
rect 528646 349398 528882 349634
rect 528326 313718 528562 313954
rect 528646 313718 528882 313954
rect 528326 313398 528562 313634
rect 528646 313398 528882 313634
rect 528326 277718 528562 277954
rect 528646 277718 528882 277954
rect 528326 277398 528562 277634
rect 528646 277398 528882 277634
rect 528326 241718 528562 241954
rect 528646 241718 528882 241954
rect 528326 241398 528562 241634
rect 528646 241398 528882 241634
rect 528326 205718 528562 205954
rect 528646 205718 528882 205954
rect 528326 205398 528562 205634
rect 528646 205398 528882 205634
rect 528326 169718 528562 169954
rect 528646 169718 528882 169954
rect 528326 169398 528562 169634
rect 528646 169398 528882 169634
rect 528326 133718 528562 133954
rect 528646 133718 528882 133954
rect 528326 133398 528562 133634
rect 528646 133398 528882 133634
rect 528326 97718 528562 97954
rect 528646 97718 528882 97954
rect 528326 97398 528562 97634
rect 528646 97398 528882 97634
rect 528326 61718 528562 61954
rect 528646 61718 528882 61954
rect 528326 61398 528562 61634
rect 528646 61398 528882 61634
rect 528326 25718 528562 25954
rect 528646 25718 528882 25954
rect 528326 25398 528562 25634
rect 528646 25398 528882 25634
rect 528326 -5382 528562 -5146
rect 528646 -5382 528882 -5146
rect 528326 -5702 528562 -5466
rect 528646 -5702 528882 -5466
rect 532826 710362 533062 710598
rect 533146 710362 533382 710598
rect 532826 710042 533062 710278
rect 533146 710042 533382 710278
rect 532826 678218 533062 678454
rect 533146 678218 533382 678454
rect 532826 677898 533062 678134
rect 533146 677898 533382 678134
rect 532826 642218 533062 642454
rect 533146 642218 533382 642454
rect 532826 641898 533062 642134
rect 533146 641898 533382 642134
rect 532826 606218 533062 606454
rect 533146 606218 533382 606454
rect 532826 605898 533062 606134
rect 533146 605898 533382 606134
rect 532826 570218 533062 570454
rect 533146 570218 533382 570454
rect 532826 569898 533062 570134
rect 533146 569898 533382 570134
rect 532826 534218 533062 534454
rect 533146 534218 533382 534454
rect 532826 533898 533062 534134
rect 533146 533898 533382 534134
rect 532826 498218 533062 498454
rect 533146 498218 533382 498454
rect 532826 497898 533062 498134
rect 533146 497898 533382 498134
rect 532826 462218 533062 462454
rect 533146 462218 533382 462454
rect 532826 461898 533062 462134
rect 533146 461898 533382 462134
rect 532826 426218 533062 426454
rect 533146 426218 533382 426454
rect 532826 425898 533062 426134
rect 533146 425898 533382 426134
rect 532826 390218 533062 390454
rect 533146 390218 533382 390454
rect 532826 389898 533062 390134
rect 533146 389898 533382 390134
rect 532826 354218 533062 354454
rect 533146 354218 533382 354454
rect 532826 353898 533062 354134
rect 533146 353898 533382 354134
rect 532826 318218 533062 318454
rect 533146 318218 533382 318454
rect 532826 317898 533062 318134
rect 533146 317898 533382 318134
rect 532826 282218 533062 282454
rect 533146 282218 533382 282454
rect 532826 281898 533062 282134
rect 533146 281898 533382 282134
rect 532826 246218 533062 246454
rect 533146 246218 533382 246454
rect 532826 245898 533062 246134
rect 533146 245898 533382 246134
rect 532826 210218 533062 210454
rect 533146 210218 533382 210454
rect 532826 209898 533062 210134
rect 533146 209898 533382 210134
rect 532826 174218 533062 174454
rect 533146 174218 533382 174454
rect 532826 173898 533062 174134
rect 533146 173898 533382 174134
rect 532826 138218 533062 138454
rect 533146 138218 533382 138454
rect 532826 137898 533062 138134
rect 533146 137898 533382 138134
rect 532826 102218 533062 102454
rect 533146 102218 533382 102454
rect 532826 101898 533062 102134
rect 533146 101898 533382 102134
rect 532826 66218 533062 66454
rect 533146 66218 533382 66454
rect 532826 65898 533062 66134
rect 533146 65898 533382 66134
rect 532826 30218 533062 30454
rect 533146 30218 533382 30454
rect 532826 29898 533062 30134
rect 533146 29898 533382 30134
rect 532826 -6342 533062 -6106
rect 533146 -6342 533382 -6106
rect 532826 -6662 533062 -6426
rect 533146 -6662 533382 -6426
rect 537326 711322 537562 711558
rect 537646 711322 537882 711558
rect 537326 711002 537562 711238
rect 537646 711002 537882 711238
rect 537326 682718 537562 682954
rect 537646 682718 537882 682954
rect 537326 682398 537562 682634
rect 537646 682398 537882 682634
rect 537326 646718 537562 646954
rect 537646 646718 537882 646954
rect 537326 646398 537562 646634
rect 537646 646398 537882 646634
rect 537326 610718 537562 610954
rect 537646 610718 537882 610954
rect 537326 610398 537562 610634
rect 537646 610398 537882 610634
rect 537326 574718 537562 574954
rect 537646 574718 537882 574954
rect 537326 574398 537562 574634
rect 537646 574398 537882 574634
rect 537326 538718 537562 538954
rect 537646 538718 537882 538954
rect 537326 538398 537562 538634
rect 537646 538398 537882 538634
rect 537326 502718 537562 502954
rect 537646 502718 537882 502954
rect 537326 502398 537562 502634
rect 537646 502398 537882 502634
rect 537326 466718 537562 466954
rect 537646 466718 537882 466954
rect 537326 466398 537562 466634
rect 537646 466398 537882 466634
rect 537326 430718 537562 430954
rect 537646 430718 537882 430954
rect 537326 430398 537562 430634
rect 537646 430398 537882 430634
rect 537326 394718 537562 394954
rect 537646 394718 537882 394954
rect 537326 394398 537562 394634
rect 537646 394398 537882 394634
rect 537326 358718 537562 358954
rect 537646 358718 537882 358954
rect 537326 358398 537562 358634
rect 537646 358398 537882 358634
rect 537326 322718 537562 322954
rect 537646 322718 537882 322954
rect 537326 322398 537562 322634
rect 537646 322398 537882 322634
rect 537326 286718 537562 286954
rect 537646 286718 537882 286954
rect 537326 286398 537562 286634
rect 537646 286398 537882 286634
rect 537326 250718 537562 250954
rect 537646 250718 537882 250954
rect 537326 250398 537562 250634
rect 537646 250398 537882 250634
rect 537326 214718 537562 214954
rect 537646 214718 537882 214954
rect 537326 214398 537562 214634
rect 537646 214398 537882 214634
rect 537326 178718 537562 178954
rect 537646 178718 537882 178954
rect 537326 178398 537562 178634
rect 537646 178398 537882 178634
rect 537326 142718 537562 142954
rect 537646 142718 537882 142954
rect 537326 142398 537562 142634
rect 537646 142398 537882 142634
rect 537326 106718 537562 106954
rect 537646 106718 537882 106954
rect 537326 106398 537562 106634
rect 537646 106398 537882 106634
rect 537326 70718 537562 70954
rect 537646 70718 537882 70954
rect 537326 70398 537562 70634
rect 537646 70398 537882 70634
rect 537326 34718 537562 34954
rect 537646 34718 537882 34954
rect 537326 34398 537562 34634
rect 537646 34398 537882 34634
rect 537326 -7302 537562 -7066
rect 537646 -7302 537882 -7066
rect 537326 -7622 537562 -7386
rect 537646 -7622 537882 -7386
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 546326 705562 546562 705798
rect 546646 705562 546882 705798
rect 546326 705242 546562 705478
rect 546646 705242 546882 705478
rect 546326 691718 546562 691954
rect 546646 691718 546882 691954
rect 546326 691398 546562 691634
rect 546646 691398 546882 691634
rect 546326 655718 546562 655954
rect 546646 655718 546882 655954
rect 546326 655398 546562 655634
rect 546646 655398 546882 655634
rect 546326 619718 546562 619954
rect 546646 619718 546882 619954
rect 546326 619398 546562 619634
rect 546646 619398 546882 619634
rect 546326 583718 546562 583954
rect 546646 583718 546882 583954
rect 546326 583398 546562 583634
rect 546646 583398 546882 583634
rect 546326 547718 546562 547954
rect 546646 547718 546882 547954
rect 546326 547398 546562 547634
rect 546646 547398 546882 547634
rect 546326 511718 546562 511954
rect 546646 511718 546882 511954
rect 546326 511398 546562 511634
rect 546646 511398 546882 511634
rect 546326 475718 546562 475954
rect 546646 475718 546882 475954
rect 546326 475398 546562 475634
rect 546646 475398 546882 475634
rect 546326 439718 546562 439954
rect 546646 439718 546882 439954
rect 546326 439398 546562 439634
rect 546646 439398 546882 439634
rect 546326 403718 546562 403954
rect 546646 403718 546882 403954
rect 546326 403398 546562 403634
rect 546646 403398 546882 403634
rect 546326 367718 546562 367954
rect 546646 367718 546882 367954
rect 546326 367398 546562 367634
rect 546646 367398 546882 367634
rect 546326 331718 546562 331954
rect 546646 331718 546882 331954
rect 546326 331398 546562 331634
rect 546646 331398 546882 331634
rect 546326 295718 546562 295954
rect 546646 295718 546882 295954
rect 546326 295398 546562 295634
rect 546646 295398 546882 295634
rect 546326 259718 546562 259954
rect 546646 259718 546882 259954
rect 546326 259398 546562 259634
rect 546646 259398 546882 259634
rect 546326 223718 546562 223954
rect 546646 223718 546882 223954
rect 546326 223398 546562 223634
rect 546646 223398 546882 223634
rect 546326 187718 546562 187954
rect 546646 187718 546882 187954
rect 546326 187398 546562 187634
rect 546646 187398 546882 187634
rect 546326 151718 546562 151954
rect 546646 151718 546882 151954
rect 546326 151398 546562 151634
rect 546646 151398 546882 151634
rect 546326 115718 546562 115954
rect 546646 115718 546882 115954
rect 546326 115398 546562 115634
rect 546646 115398 546882 115634
rect 546326 79718 546562 79954
rect 546646 79718 546882 79954
rect 546326 79398 546562 79634
rect 546646 79398 546882 79634
rect 546326 43718 546562 43954
rect 546646 43718 546882 43954
rect 546326 43398 546562 43634
rect 546646 43398 546882 43634
rect 546326 7718 546562 7954
rect 546646 7718 546882 7954
rect 546326 7398 546562 7634
rect 546646 7398 546882 7634
rect 546326 -1542 546562 -1306
rect 546646 -1542 546882 -1306
rect 546326 -1862 546562 -1626
rect 546646 -1862 546882 -1626
rect 550826 706522 551062 706758
rect 551146 706522 551382 706758
rect 550826 706202 551062 706438
rect 551146 706202 551382 706438
rect 550826 696218 551062 696454
rect 551146 696218 551382 696454
rect 550826 695898 551062 696134
rect 551146 695898 551382 696134
rect 550826 660218 551062 660454
rect 551146 660218 551382 660454
rect 550826 659898 551062 660134
rect 551146 659898 551382 660134
rect 550826 624218 551062 624454
rect 551146 624218 551382 624454
rect 550826 623898 551062 624134
rect 551146 623898 551382 624134
rect 550826 588218 551062 588454
rect 551146 588218 551382 588454
rect 550826 587898 551062 588134
rect 551146 587898 551382 588134
rect 550826 552218 551062 552454
rect 551146 552218 551382 552454
rect 550826 551898 551062 552134
rect 551146 551898 551382 552134
rect 550826 516218 551062 516454
rect 551146 516218 551382 516454
rect 550826 515898 551062 516134
rect 551146 515898 551382 516134
rect 550826 480218 551062 480454
rect 551146 480218 551382 480454
rect 550826 479898 551062 480134
rect 551146 479898 551382 480134
rect 550826 444218 551062 444454
rect 551146 444218 551382 444454
rect 550826 443898 551062 444134
rect 551146 443898 551382 444134
rect 550826 408218 551062 408454
rect 551146 408218 551382 408454
rect 550826 407898 551062 408134
rect 551146 407898 551382 408134
rect 550826 372218 551062 372454
rect 551146 372218 551382 372454
rect 550826 371898 551062 372134
rect 551146 371898 551382 372134
rect 550826 336218 551062 336454
rect 551146 336218 551382 336454
rect 550826 335898 551062 336134
rect 551146 335898 551382 336134
rect 550826 300218 551062 300454
rect 551146 300218 551382 300454
rect 550826 299898 551062 300134
rect 551146 299898 551382 300134
rect 550826 264218 551062 264454
rect 551146 264218 551382 264454
rect 550826 263898 551062 264134
rect 551146 263898 551382 264134
rect 550826 228218 551062 228454
rect 551146 228218 551382 228454
rect 550826 227898 551062 228134
rect 551146 227898 551382 228134
rect 550826 192218 551062 192454
rect 551146 192218 551382 192454
rect 550826 191898 551062 192134
rect 551146 191898 551382 192134
rect 550826 156218 551062 156454
rect 551146 156218 551382 156454
rect 550826 155898 551062 156134
rect 551146 155898 551382 156134
rect 550826 120218 551062 120454
rect 551146 120218 551382 120454
rect 550826 119898 551062 120134
rect 551146 119898 551382 120134
rect 550826 84218 551062 84454
rect 551146 84218 551382 84454
rect 550826 83898 551062 84134
rect 551146 83898 551382 84134
rect 550826 48218 551062 48454
rect 551146 48218 551382 48454
rect 550826 47898 551062 48134
rect 551146 47898 551382 48134
rect 550826 12218 551062 12454
rect 551146 12218 551382 12454
rect 550826 11898 551062 12134
rect 551146 11898 551382 12134
rect 550826 -2502 551062 -2266
rect 551146 -2502 551382 -2266
rect 550826 -2822 551062 -2586
rect 551146 -2822 551382 -2586
rect 555326 707482 555562 707718
rect 555646 707482 555882 707718
rect 555326 707162 555562 707398
rect 555646 707162 555882 707398
rect 555326 700718 555562 700954
rect 555646 700718 555882 700954
rect 555326 700398 555562 700634
rect 555646 700398 555882 700634
rect 555326 664718 555562 664954
rect 555646 664718 555882 664954
rect 555326 664398 555562 664634
rect 555646 664398 555882 664634
rect 555326 628718 555562 628954
rect 555646 628718 555882 628954
rect 555326 628398 555562 628634
rect 555646 628398 555882 628634
rect 555326 592718 555562 592954
rect 555646 592718 555882 592954
rect 555326 592398 555562 592634
rect 555646 592398 555882 592634
rect 555326 556718 555562 556954
rect 555646 556718 555882 556954
rect 555326 556398 555562 556634
rect 555646 556398 555882 556634
rect 555326 520718 555562 520954
rect 555646 520718 555882 520954
rect 555326 520398 555562 520634
rect 555646 520398 555882 520634
rect 555326 484718 555562 484954
rect 555646 484718 555882 484954
rect 555326 484398 555562 484634
rect 555646 484398 555882 484634
rect 555326 448718 555562 448954
rect 555646 448718 555882 448954
rect 555326 448398 555562 448634
rect 555646 448398 555882 448634
rect 555326 412718 555562 412954
rect 555646 412718 555882 412954
rect 555326 412398 555562 412634
rect 555646 412398 555882 412634
rect 555326 376718 555562 376954
rect 555646 376718 555882 376954
rect 555326 376398 555562 376634
rect 555646 376398 555882 376634
rect 555326 340718 555562 340954
rect 555646 340718 555882 340954
rect 555326 340398 555562 340634
rect 555646 340398 555882 340634
rect 555326 304718 555562 304954
rect 555646 304718 555882 304954
rect 555326 304398 555562 304634
rect 555646 304398 555882 304634
rect 555326 268718 555562 268954
rect 555646 268718 555882 268954
rect 555326 268398 555562 268634
rect 555646 268398 555882 268634
rect 555326 232718 555562 232954
rect 555646 232718 555882 232954
rect 555326 232398 555562 232634
rect 555646 232398 555882 232634
rect 555326 196718 555562 196954
rect 555646 196718 555882 196954
rect 555326 196398 555562 196634
rect 555646 196398 555882 196634
rect 555326 160718 555562 160954
rect 555646 160718 555882 160954
rect 555326 160398 555562 160634
rect 555646 160398 555882 160634
rect 555326 124718 555562 124954
rect 555646 124718 555882 124954
rect 555326 124398 555562 124634
rect 555646 124398 555882 124634
rect 555326 88718 555562 88954
rect 555646 88718 555882 88954
rect 555326 88398 555562 88634
rect 555646 88398 555882 88634
rect 555326 52718 555562 52954
rect 555646 52718 555882 52954
rect 555326 52398 555562 52634
rect 555646 52398 555882 52634
rect 555326 16718 555562 16954
rect 555646 16718 555882 16954
rect 555326 16398 555562 16634
rect 555646 16398 555882 16634
rect 555326 -3462 555562 -3226
rect 555646 -3462 555882 -3226
rect 555326 -3782 555562 -3546
rect 555646 -3782 555882 -3546
rect 559826 708442 560062 708678
rect 560146 708442 560382 708678
rect 559826 708122 560062 708358
rect 560146 708122 560382 708358
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -4422 560062 -4186
rect 560146 -4422 560382 -4186
rect 559826 -4742 560062 -4506
rect 560146 -4742 560382 -4506
rect 564326 709402 564562 709638
rect 564646 709402 564882 709638
rect 564326 709082 564562 709318
rect 564646 709082 564882 709318
rect 564326 673718 564562 673954
rect 564646 673718 564882 673954
rect 564326 673398 564562 673634
rect 564646 673398 564882 673634
rect 564326 637718 564562 637954
rect 564646 637718 564882 637954
rect 564326 637398 564562 637634
rect 564646 637398 564882 637634
rect 564326 601718 564562 601954
rect 564646 601718 564882 601954
rect 564326 601398 564562 601634
rect 564646 601398 564882 601634
rect 564326 565718 564562 565954
rect 564646 565718 564882 565954
rect 564326 565398 564562 565634
rect 564646 565398 564882 565634
rect 564326 529718 564562 529954
rect 564646 529718 564882 529954
rect 564326 529398 564562 529634
rect 564646 529398 564882 529634
rect 564326 493718 564562 493954
rect 564646 493718 564882 493954
rect 564326 493398 564562 493634
rect 564646 493398 564882 493634
rect 564326 457718 564562 457954
rect 564646 457718 564882 457954
rect 564326 457398 564562 457634
rect 564646 457398 564882 457634
rect 564326 421718 564562 421954
rect 564646 421718 564882 421954
rect 564326 421398 564562 421634
rect 564646 421398 564882 421634
rect 564326 385718 564562 385954
rect 564646 385718 564882 385954
rect 564326 385398 564562 385634
rect 564646 385398 564882 385634
rect 564326 349718 564562 349954
rect 564646 349718 564882 349954
rect 564326 349398 564562 349634
rect 564646 349398 564882 349634
rect 564326 313718 564562 313954
rect 564646 313718 564882 313954
rect 564326 313398 564562 313634
rect 564646 313398 564882 313634
rect 564326 277718 564562 277954
rect 564646 277718 564882 277954
rect 564326 277398 564562 277634
rect 564646 277398 564882 277634
rect 564326 241718 564562 241954
rect 564646 241718 564882 241954
rect 564326 241398 564562 241634
rect 564646 241398 564882 241634
rect 564326 205718 564562 205954
rect 564646 205718 564882 205954
rect 564326 205398 564562 205634
rect 564646 205398 564882 205634
rect 564326 169718 564562 169954
rect 564646 169718 564882 169954
rect 564326 169398 564562 169634
rect 564646 169398 564882 169634
rect 564326 133718 564562 133954
rect 564646 133718 564882 133954
rect 564326 133398 564562 133634
rect 564646 133398 564882 133634
rect 564326 97718 564562 97954
rect 564646 97718 564882 97954
rect 564326 97398 564562 97634
rect 564646 97398 564882 97634
rect 564326 61718 564562 61954
rect 564646 61718 564882 61954
rect 564326 61398 564562 61634
rect 564646 61398 564882 61634
rect 564326 25718 564562 25954
rect 564646 25718 564882 25954
rect 564326 25398 564562 25634
rect 564646 25398 564882 25634
rect 564326 -5382 564562 -5146
rect 564646 -5382 564882 -5146
rect 564326 -5702 564562 -5466
rect 564646 -5702 564882 -5466
rect 568826 710362 569062 710598
rect 569146 710362 569382 710598
rect 568826 710042 569062 710278
rect 569146 710042 569382 710278
rect 568826 678218 569062 678454
rect 569146 678218 569382 678454
rect 568826 677898 569062 678134
rect 569146 677898 569382 678134
rect 568826 642218 569062 642454
rect 569146 642218 569382 642454
rect 568826 641898 569062 642134
rect 569146 641898 569382 642134
rect 568826 606218 569062 606454
rect 569146 606218 569382 606454
rect 568826 605898 569062 606134
rect 569146 605898 569382 606134
rect 568826 570218 569062 570454
rect 569146 570218 569382 570454
rect 568826 569898 569062 570134
rect 569146 569898 569382 570134
rect 568826 534218 569062 534454
rect 569146 534218 569382 534454
rect 568826 533898 569062 534134
rect 569146 533898 569382 534134
rect 568826 498218 569062 498454
rect 569146 498218 569382 498454
rect 568826 497898 569062 498134
rect 569146 497898 569382 498134
rect 568826 462218 569062 462454
rect 569146 462218 569382 462454
rect 568826 461898 569062 462134
rect 569146 461898 569382 462134
rect 568826 426218 569062 426454
rect 569146 426218 569382 426454
rect 568826 425898 569062 426134
rect 569146 425898 569382 426134
rect 568826 390218 569062 390454
rect 569146 390218 569382 390454
rect 568826 389898 569062 390134
rect 569146 389898 569382 390134
rect 568826 354218 569062 354454
rect 569146 354218 569382 354454
rect 568826 353898 569062 354134
rect 569146 353898 569382 354134
rect 568826 318218 569062 318454
rect 569146 318218 569382 318454
rect 568826 317898 569062 318134
rect 569146 317898 569382 318134
rect 568826 282218 569062 282454
rect 569146 282218 569382 282454
rect 568826 281898 569062 282134
rect 569146 281898 569382 282134
rect 568826 246218 569062 246454
rect 569146 246218 569382 246454
rect 568826 245898 569062 246134
rect 569146 245898 569382 246134
rect 568826 210218 569062 210454
rect 569146 210218 569382 210454
rect 568826 209898 569062 210134
rect 569146 209898 569382 210134
rect 568826 174218 569062 174454
rect 569146 174218 569382 174454
rect 568826 173898 569062 174134
rect 569146 173898 569382 174134
rect 568826 138218 569062 138454
rect 569146 138218 569382 138454
rect 568826 137898 569062 138134
rect 569146 137898 569382 138134
rect 568826 102218 569062 102454
rect 569146 102218 569382 102454
rect 568826 101898 569062 102134
rect 569146 101898 569382 102134
rect 568826 66218 569062 66454
rect 569146 66218 569382 66454
rect 568826 65898 569062 66134
rect 569146 65898 569382 66134
rect 568826 30218 569062 30454
rect 569146 30218 569382 30454
rect 568826 29898 569062 30134
rect 569146 29898 569382 30134
rect 568826 -6342 569062 -6106
rect 569146 -6342 569382 -6106
rect 568826 -6662 569062 -6426
rect 569146 -6662 569382 -6426
rect 573326 711322 573562 711558
rect 573646 711322 573882 711558
rect 573326 711002 573562 711238
rect 573646 711002 573882 711238
rect 573326 682718 573562 682954
rect 573646 682718 573882 682954
rect 573326 682398 573562 682634
rect 573646 682398 573882 682634
rect 573326 646718 573562 646954
rect 573646 646718 573882 646954
rect 573326 646398 573562 646634
rect 573646 646398 573882 646634
rect 573326 610718 573562 610954
rect 573646 610718 573882 610954
rect 573326 610398 573562 610634
rect 573646 610398 573882 610634
rect 573326 574718 573562 574954
rect 573646 574718 573882 574954
rect 573326 574398 573562 574634
rect 573646 574398 573882 574634
rect 573326 538718 573562 538954
rect 573646 538718 573882 538954
rect 573326 538398 573562 538634
rect 573646 538398 573882 538634
rect 573326 502718 573562 502954
rect 573646 502718 573882 502954
rect 573326 502398 573562 502634
rect 573646 502398 573882 502634
rect 573326 466718 573562 466954
rect 573646 466718 573882 466954
rect 573326 466398 573562 466634
rect 573646 466398 573882 466634
rect 573326 430718 573562 430954
rect 573646 430718 573882 430954
rect 573326 430398 573562 430634
rect 573646 430398 573882 430634
rect 573326 394718 573562 394954
rect 573646 394718 573882 394954
rect 573326 394398 573562 394634
rect 573646 394398 573882 394634
rect 573326 358718 573562 358954
rect 573646 358718 573882 358954
rect 573326 358398 573562 358634
rect 573646 358398 573882 358634
rect 573326 322718 573562 322954
rect 573646 322718 573882 322954
rect 573326 322398 573562 322634
rect 573646 322398 573882 322634
rect 573326 286718 573562 286954
rect 573646 286718 573882 286954
rect 573326 286398 573562 286634
rect 573646 286398 573882 286634
rect 573326 250718 573562 250954
rect 573646 250718 573882 250954
rect 573326 250398 573562 250634
rect 573646 250398 573882 250634
rect 573326 214718 573562 214954
rect 573646 214718 573882 214954
rect 573326 214398 573562 214634
rect 573646 214398 573882 214634
rect 573326 178718 573562 178954
rect 573646 178718 573882 178954
rect 573326 178398 573562 178634
rect 573646 178398 573882 178634
rect 573326 142718 573562 142954
rect 573646 142718 573882 142954
rect 573326 142398 573562 142634
rect 573646 142398 573882 142634
rect 573326 106718 573562 106954
rect 573646 106718 573882 106954
rect 573326 106398 573562 106634
rect 573646 106398 573882 106634
rect 573326 70718 573562 70954
rect 573646 70718 573882 70954
rect 573326 70398 573562 70634
rect 573646 70398 573882 70634
rect 573326 34718 573562 34954
rect 573646 34718 573882 34954
rect 573326 34398 573562 34634
rect 573646 34398 573882 34634
rect 573326 -7302 573562 -7066
rect 573646 -7302 573882 -7066
rect 573326 -7622 573562 -7386
rect 573646 -7622 573882 -7386
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 582326 705562 582562 705798
rect 582646 705562 582882 705798
rect 582326 705242 582562 705478
rect 582646 705242 582882 705478
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 582326 691718 582562 691954
rect 582646 691718 582882 691954
rect 582326 691398 582562 691634
rect 582646 691398 582882 691634
rect 582326 655718 582562 655954
rect 582646 655718 582882 655954
rect 582326 655398 582562 655634
rect 582646 655398 582882 655634
rect 582326 619718 582562 619954
rect 582646 619718 582882 619954
rect 582326 619398 582562 619634
rect 582646 619398 582882 619634
rect 582326 583718 582562 583954
rect 582646 583718 582882 583954
rect 582326 583398 582562 583634
rect 582646 583398 582882 583634
rect 582326 547718 582562 547954
rect 582646 547718 582882 547954
rect 582326 547398 582562 547634
rect 582646 547398 582882 547634
rect 582326 511718 582562 511954
rect 582646 511718 582882 511954
rect 582326 511398 582562 511634
rect 582646 511398 582882 511634
rect 582326 475718 582562 475954
rect 582646 475718 582882 475954
rect 582326 475398 582562 475634
rect 582646 475398 582882 475634
rect 582326 439718 582562 439954
rect 582646 439718 582882 439954
rect 582326 439398 582562 439634
rect 582646 439398 582882 439634
rect 582326 403718 582562 403954
rect 582646 403718 582882 403954
rect 582326 403398 582562 403634
rect 582646 403398 582882 403634
rect 582326 367718 582562 367954
rect 582646 367718 582882 367954
rect 582326 367398 582562 367634
rect 582646 367398 582882 367634
rect 582326 331718 582562 331954
rect 582646 331718 582882 331954
rect 582326 331398 582562 331634
rect 582646 331398 582882 331634
rect 582326 295718 582562 295954
rect 582646 295718 582882 295954
rect 582326 295398 582562 295634
rect 582646 295398 582882 295634
rect 582326 259718 582562 259954
rect 582646 259718 582882 259954
rect 582326 259398 582562 259634
rect 582646 259398 582882 259634
rect 582326 223718 582562 223954
rect 582646 223718 582882 223954
rect 582326 223398 582562 223634
rect 582646 223398 582882 223634
rect 582326 187718 582562 187954
rect 582646 187718 582882 187954
rect 582326 187398 582562 187634
rect 582646 187398 582882 187634
rect 582326 151718 582562 151954
rect 582646 151718 582882 151954
rect 582326 151398 582562 151634
rect 582646 151398 582882 151634
rect 582326 115718 582562 115954
rect 582646 115718 582882 115954
rect 582326 115398 582562 115634
rect 582646 115398 582882 115634
rect 582326 79718 582562 79954
rect 582646 79718 582882 79954
rect 582326 79398 582562 79634
rect 582646 79398 582882 79634
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 582326 43718 582562 43954
rect 582646 43718 582882 43954
rect 582326 43398 582562 43634
rect 582646 43398 582882 43634
rect 582326 7718 582562 7954
rect 582646 7718 582882 7954
rect 582326 7398 582562 7634
rect 582646 7398 582882 7634
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 691718 586538 691954
rect 586622 691718 586858 691954
rect 586302 691398 586538 691634
rect 586622 691398 586858 691634
rect 586302 655718 586538 655954
rect 586622 655718 586858 655954
rect 586302 655398 586538 655634
rect 586622 655398 586858 655634
rect 586302 619718 586538 619954
rect 586622 619718 586858 619954
rect 586302 619398 586538 619634
rect 586622 619398 586858 619634
rect 586302 583718 586538 583954
rect 586622 583718 586858 583954
rect 586302 583398 586538 583634
rect 586622 583398 586858 583634
rect 586302 547718 586538 547954
rect 586622 547718 586858 547954
rect 586302 547398 586538 547634
rect 586622 547398 586858 547634
rect 586302 511718 586538 511954
rect 586622 511718 586858 511954
rect 586302 511398 586538 511634
rect 586622 511398 586858 511634
rect 586302 475718 586538 475954
rect 586622 475718 586858 475954
rect 586302 475398 586538 475634
rect 586622 475398 586858 475634
rect 586302 439718 586538 439954
rect 586622 439718 586858 439954
rect 586302 439398 586538 439634
rect 586622 439398 586858 439634
rect 586302 403718 586538 403954
rect 586622 403718 586858 403954
rect 586302 403398 586538 403634
rect 586622 403398 586858 403634
rect 586302 367718 586538 367954
rect 586622 367718 586858 367954
rect 586302 367398 586538 367634
rect 586622 367398 586858 367634
rect 586302 331718 586538 331954
rect 586622 331718 586858 331954
rect 586302 331398 586538 331634
rect 586622 331398 586858 331634
rect 586302 295718 586538 295954
rect 586622 295718 586858 295954
rect 586302 295398 586538 295634
rect 586622 295398 586858 295634
rect 586302 259718 586538 259954
rect 586622 259718 586858 259954
rect 586302 259398 586538 259634
rect 586622 259398 586858 259634
rect 586302 223718 586538 223954
rect 586622 223718 586858 223954
rect 586302 223398 586538 223634
rect 586622 223398 586858 223634
rect 586302 187718 586538 187954
rect 586622 187718 586858 187954
rect 586302 187398 586538 187634
rect 586622 187398 586858 187634
rect 586302 151718 586538 151954
rect 586622 151718 586858 151954
rect 586302 151398 586538 151634
rect 586622 151398 586858 151634
rect 586302 115718 586538 115954
rect 586622 115718 586858 115954
rect 586302 115398 586538 115634
rect 586622 115398 586858 115634
rect 586302 79718 586538 79954
rect 586622 79718 586858 79954
rect 586302 79398 586538 79634
rect 586622 79398 586858 79634
rect 586302 43718 586538 43954
rect 586622 43718 586858 43954
rect 586302 43398 586538 43634
rect 586622 43398 586858 43634
rect 586302 7718 586538 7954
rect 586622 7718 586858 7954
rect 586302 7398 586538 7634
rect 586622 7398 586858 7634
rect 582326 -1542 582562 -1306
rect 582646 -1542 582882 -1306
rect 582326 -1862 582562 -1626
rect 582646 -1862 582882 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 696218 587498 696454
rect 587582 696218 587818 696454
rect 587262 695898 587498 696134
rect 587582 695898 587818 696134
rect 587262 660218 587498 660454
rect 587582 660218 587818 660454
rect 587262 659898 587498 660134
rect 587582 659898 587818 660134
rect 587262 624218 587498 624454
rect 587582 624218 587818 624454
rect 587262 623898 587498 624134
rect 587582 623898 587818 624134
rect 587262 588218 587498 588454
rect 587582 588218 587818 588454
rect 587262 587898 587498 588134
rect 587582 587898 587818 588134
rect 587262 552218 587498 552454
rect 587582 552218 587818 552454
rect 587262 551898 587498 552134
rect 587582 551898 587818 552134
rect 587262 516218 587498 516454
rect 587582 516218 587818 516454
rect 587262 515898 587498 516134
rect 587582 515898 587818 516134
rect 587262 480218 587498 480454
rect 587582 480218 587818 480454
rect 587262 479898 587498 480134
rect 587582 479898 587818 480134
rect 587262 444218 587498 444454
rect 587582 444218 587818 444454
rect 587262 443898 587498 444134
rect 587582 443898 587818 444134
rect 587262 408218 587498 408454
rect 587582 408218 587818 408454
rect 587262 407898 587498 408134
rect 587582 407898 587818 408134
rect 587262 372218 587498 372454
rect 587582 372218 587818 372454
rect 587262 371898 587498 372134
rect 587582 371898 587818 372134
rect 587262 336218 587498 336454
rect 587582 336218 587818 336454
rect 587262 335898 587498 336134
rect 587582 335898 587818 336134
rect 587262 300218 587498 300454
rect 587582 300218 587818 300454
rect 587262 299898 587498 300134
rect 587582 299898 587818 300134
rect 587262 264218 587498 264454
rect 587582 264218 587818 264454
rect 587262 263898 587498 264134
rect 587582 263898 587818 264134
rect 587262 228218 587498 228454
rect 587582 228218 587818 228454
rect 587262 227898 587498 228134
rect 587582 227898 587818 228134
rect 587262 192218 587498 192454
rect 587582 192218 587818 192454
rect 587262 191898 587498 192134
rect 587582 191898 587818 192134
rect 587262 156218 587498 156454
rect 587582 156218 587818 156454
rect 587262 155898 587498 156134
rect 587582 155898 587818 156134
rect 587262 120218 587498 120454
rect 587582 120218 587818 120454
rect 587262 119898 587498 120134
rect 587582 119898 587818 120134
rect 587262 84218 587498 84454
rect 587582 84218 587818 84454
rect 587262 83898 587498 84134
rect 587582 83898 587818 84134
rect 587262 48218 587498 48454
rect 587582 48218 587818 48454
rect 587262 47898 587498 48134
rect 587582 47898 587818 48134
rect 587262 12218 587498 12454
rect 587582 12218 587818 12454
rect 587262 11898 587498 12134
rect 587582 11898 587818 12134
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 700718 588458 700954
rect 588542 700718 588778 700954
rect 588222 700398 588458 700634
rect 588542 700398 588778 700634
rect 588222 664718 588458 664954
rect 588542 664718 588778 664954
rect 588222 664398 588458 664634
rect 588542 664398 588778 664634
rect 588222 628718 588458 628954
rect 588542 628718 588778 628954
rect 588222 628398 588458 628634
rect 588542 628398 588778 628634
rect 588222 592718 588458 592954
rect 588542 592718 588778 592954
rect 588222 592398 588458 592634
rect 588542 592398 588778 592634
rect 588222 556718 588458 556954
rect 588542 556718 588778 556954
rect 588222 556398 588458 556634
rect 588542 556398 588778 556634
rect 588222 520718 588458 520954
rect 588542 520718 588778 520954
rect 588222 520398 588458 520634
rect 588542 520398 588778 520634
rect 588222 484718 588458 484954
rect 588542 484718 588778 484954
rect 588222 484398 588458 484634
rect 588542 484398 588778 484634
rect 588222 448718 588458 448954
rect 588542 448718 588778 448954
rect 588222 448398 588458 448634
rect 588542 448398 588778 448634
rect 588222 412718 588458 412954
rect 588542 412718 588778 412954
rect 588222 412398 588458 412634
rect 588542 412398 588778 412634
rect 588222 376718 588458 376954
rect 588542 376718 588778 376954
rect 588222 376398 588458 376634
rect 588542 376398 588778 376634
rect 588222 340718 588458 340954
rect 588542 340718 588778 340954
rect 588222 340398 588458 340634
rect 588542 340398 588778 340634
rect 588222 304718 588458 304954
rect 588542 304718 588778 304954
rect 588222 304398 588458 304634
rect 588542 304398 588778 304634
rect 588222 268718 588458 268954
rect 588542 268718 588778 268954
rect 588222 268398 588458 268634
rect 588542 268398 588778 268634
rect 588222 232718 588458 232954
rect 588542 232718 588778 232954
rect 588222 232398 588458 232634
rect 588542 232398 588778 232634
rect 588222 196718 588458 196954
rect 588542 196718 588778 196954
rect 588222 196398 588458 196634
rect 588542 196398 588778 196634
rect 588222 160718 588458 160954
rect 588542 160718 588778 160954
rect 588222 160398 588458 160634
rect 588542 160398 588778 160634
rect 588222 124718 588458 124954
rect 588542 124718 588778 124954
rect 588222 124398 588458 124634
rect 588542 124398 588778 124634
rect 588222 88718 588458 88954
rect 588542 88718 588778 88954
rect 588222 88398 588458 88634
rect 588542 88398 588778 88634
rect 588222 52718 588458 52954
rect 588542 52718 588778 52954
rect 588222 52398 588458 52634
rect 588542 52398 588778 52634
rect 588222 16718 588458 16954
rect 588542 16718 588778 16954
rect 588222 16398 588458 16634
rect 588542 16398 588778 16634
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 669218 589418 669454
rect 589502 669218 589738 669454
rect 589182 668898 589418 669134
rect 589502 668898 589738 669134
rect 589182 633218 589418 633454
rect 589502 633218 589738 633454
rect 589182 632898 589418 633134
rect 589502 632898 589738 633134
rect 589182 597218 589418 597454
rect 589502 597218 589738 597454
rect 589182 596898 589418 597134
rect 589502 596898 589738 597134
rect 589182 561218 589418 561454
rect 589502 561218 589738 561454
rect 589182 560898 589418 561134
rect 589502 560898 589738 561134
rect 589182 525218 589418 525454
rect 589502 525218 589738 525454
rect 589182 524898 589418 525134
rect 589502 524898 589738 525134
rect 589182 489218 589418 489454
rect 589502 489218 589738 489454
rect 589182 488898 589418 489134
rect 589502 488898 589738 489134
rect 589182 453218 589418 453454
rect 589502 453218 589738 453454
rect 589182 452898 589418 453134
rect 589502 452898 589738 453134
rect 589182 417218 589418 417454
rect 589502 417218 589738 417454
rect 589182 416898 589418 417134
rect 589502 416898 589738 417134
rect 589182 381218 589418 381454
rect 589502 381218 589738 381454
rect 589182 380898 589418 381134
rect 589502 380898 589738 381134
rect 589182 345218 589418 345454
rect 589502 345218 589738 345454
rect 589182 344898 589418 345134
rect 589502 344898 589738 345134
rect 589182 309218 589418 309454
rect 589502 309218 589738 309454
rect 589182 308898 589418 309134
rect 589502 308898 589738 309134
rect 589182 273218 589418 273454
rect 589502 273218 589738 273454
rect 589182 272898 589418 273134
rect 589502 272898 589738 273134
rect 589182 237218 589418 237454
rect 589502 237218 589738 237454
rect 589182 236898 589418 237134
rect 589502 236898 589738 237134
rect 589182 201218 589418 201454
rect 589502 201218 589738 201454
rect 589182 200898 589418 201134
rect 589502 200898 589738 201134
rect 589182 165218 589418 165454
rect 589502 165218 589738 165454
rect 589182 164898 589418 165134
rect 589502 164898 589738 165134
rect 589182 129218 589418 129454
rect 589502 129218 589738 129454
rect 589182 128898 589418 129134
rect 589502 128898 589738 129134
rect 589182 93218 589418 93454
rect 589502 93218 589738 93454
rect 589182 92898 589418 93134
rect 589502 92898 589738 93134
rect 589182 57218 589418 57454
rect 589502 57218 589738 57454
rect 589182 56898 589418 57134
rect 589502 56898 589738 57134
rect 589182 21218 589418 21454
rect 589502 21218 589738 21454
rect 589182 20898 589418 21134
rect 589502 20898 589738 21134
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 673718 590378 673954
rect 590462 673718 590698 673954
rect 590142 673398 590378 673634
rect 590462 673398 590698 673634
rect 590142 637718 590378 637954
rect 590462 637718 590698 637954
rect 590142 637398 590378 637634
rect 590462 637398 590698 637634
rect 590142 601718 590378 601954
rect 590462 601718 590698 601954
rect 590142 601398 590378 601634
rect 590462 601398 590698 601634
rect 590142 565718 590378 565954
rect 590462 565718 590698 565954
rect 590142 565398 590378 565634
rect 590462 565398 590698 565634
rect 590142 529718 590378 529954
rect 590462 529718 590698 529954
rect 590142 529398 590378 529634
rect 590462 529398 590698 529634
rect 590142 493718 590378 493954
rect 590462 493718 590698 493954
rect 590142 493398 590378 493634
rect 590462 493398 590698 493634
rect 590142 457718 590378 457954
rect 590462 457718 590698 457954
rect 590142 457398 590378 457634
rect 590462 457398 590698 457634
rect 590142 421718 590378 421954
rect 590462 421718 590698 421954
rect 590142 421398 590378 421634
rect 590462 421398 590698 421634
rect 590142 385718 590378 385954
rect 590462 385718 590698 385954
rect 590142 385398 590378 385634
rect 590462 385398 590698 385634
rect 590142 349718 590378 349954
rect 590462 349718 590698 349954
rect 590142 349398 590378 349634
rect 590462 349398 590698 349634
rect 590142 313718 590378 313954
rect 590462 313718 590698 313954
rect 590142 313398 590378 313634
rect 590462 313398 590698 313634
rect 590142 277718 590378 277954
rect 590462 277718 590698 277954
rect 590142 277398 590378 277634
rect 590462 277398 590698 277634
rect 590142 241718 590378 241954
rect 590462 241718 590698 241954
rect 590142 241398 590378 241634
rect 590462 241398 590698 241634
rect 590142 205718 590378 205954
rect 590462 205718 590698 205954
rect 590142 205398 590378 205634
rect 590462 205398 590698 205634
rect 590142 169718 590378 169954
rect 590462 169718 590698 169954
rect 590142 169398 590378 169634
rect 590462 169398 590698 169634
rect 590142 133718 590378 133954
rect 590462 133718 590698 133954
rect 590142 133398 590378 133634
rect 590462 133398 590698 133634
rect 590142 97718 590378 97954
rect 590462 97718 590698 97954
rect 590142 97398 590378 97634
rect 590462 97398 590698 97634
rect 590142 61718 590378 61954
rect 590462 61718 590698 61954
rect 590142 61398 590378 61634
rect 590462 61398 590698 61634
rect 590142 25718 590378 25954
rect 590462 25718 590698 25954
rect 590142 25398 590378 25634
rect 590462 25398 590698 25634
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 678218 591338 678454
rect 591422 678218 591658 678454
rect 591102 677898 591338 678134
rect 591422 677898 591658 678134
rect 591102 642218 591338 642454
rect 591422 642218 591658 642454
rect 591102 641898 591338 642134
rect 591422 641898 591658 642134
rect 591102 606218 591338 606454
rect 591422 606218 591658 606454
rect 591102 605898 591338 606134
rect 591422 605898 591658 606134
rect 591102 570218 591338 570454
rect 591422 570218 591658 570454
rect 591102 569898 591338 570134
rect 591422 569898 591658 570134
rect 591102 534218 591338 534454
rect 591422 534218 591658 534454
rect 591102 533898 591338 534134
rect 591422 533898 591658 534134
rect 591102 498218 591338 498454
rect 591422 498218 591658 498454
rect 591102 497898 591338 498134
rect 591422 497898 591658 498134
rect 591102 462218 591338 462454
rect 591422 462218 591658 462454
rect 591102 461898 591338 462134
rect 591422 461898 591658 462134
rect 591102 426218 591338 426454
rect 591422 426218 591658 426454
rect 591102 425898 591338 426134
rect 591422 425898 591658 426134
rect 591102 390218 591338 390454
rect 591422 390218 591658 390454
rect 591102 389898 591338 390134
rect 591422 389898 591658 390134
rect 591102 354218 591338 354454
rect 591422 354218 591658 354454
rect 591102 353898 591338 354134
rect 591422 353898 591658 354134
rect 591102 318218 591338 318454
rect 591422 318218 591658 318454
rect 591102 317898 591338 318134
rect 591422 317898 591658 318134
rect 591102 282218 591338 282454
rect 591422 282218 591658 282454
rect 591102 281898 591338 282134
rect 591422 281898 591658 282134
rect 591102 246218 591338 246454
rect 591422 246218 591658 246454
rect 591102 245898 591338 246134
rect 591422 245898 591658 246134
rect 591102 210218 591338 210454
rect 591422 210218 591658 210454
rect 591102 209898 591338 210134
rect 591422 209898 591658 210134
rect 591102 174218 591338 174454
rect 591422 174218 591658 174454
rect 591102 173898 591338 174134
rect 591422 173898 591658 174134
rect 591102 138218 591338 138454
rect 591422 138218 591658 138454
rect 591102 137898 591338 138134
rect 591422 137898 591658 138134
rect 591102 102218 591338 102454
rect 591422 102218 591658 102454
rect 591102 101898 591338 102134
rect 591422 101898 591658 102134
rect 591102 66218 591338 66454
rect 591422 66218 591658 66454
rect 591102 65898 591338 66134
rect 591422 65898 591658 66134
rect 591102 30218 591338 30454
rect 591422 30218 591658 30454
rect 591102 29898 591338 30134
rect 591422 29898 591658 30134
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 682718 592298 682954
rect 592382 682718 592618 682954
rect 592062 682398 592298 682634
rect 592382 682398 592618 682634
rect 592062 646718 592298 646954
rect 592382 646718 592618 646954
rect 592062 646398 592298 646634
rect 592382 646398 592618 646634
rect 592062 610718 592298 610954
rect 592382 610718 592618 610954
rect 592062 610398 592298 610634
rect 592382 610398 592618 610634
rect 592062 574718 592298 574954
rect 592382 574718 592618 574954
rect 592062 574398 592298 574634
rect 592382 574398 592618 574634
rect 592062 538718 592298 538954
rect 592382 538718 592618 538954
rect 592062 538398 592298 538634
rect 592382 538398 592618 538634
rect 592062 502718 592298 502954
rect 592382 502718 592618 502954
rect 592062 502398 592298 502634
rect 592382 502398 592618 502634
rect 592062 466718 592298 466954
rect 592382 466718 592618 466954
rect 592062 466398 592298 466634
rect 592382 466398 592618 466634
rect 592062 430718 592298 430954
rect 592382 430718 592618 430954
rect 592062 430398 592298 430634
rect 592382 430398 592618 430634
rect 592062 394718 592298 394954
rect 592382 394718 592618 394954
rect 592062 394398 592298 394634
rect 592382 394398 592618 394634
rect 592062 358718 592298 358954
rect 592382 358718 592618 358954
rect 592062 358398 592298 358634
rect 592382 358398 592618 358634
rect 592062 322718 592298 322954
rect 592382 322718 592618 322954
rect 592062 322398 592298 322634
rect 592382 322398 592618 322634
rect 592062 286718 592298 286954
rect 592382 286718 592618 286954
rect 592062 286398 592298 286634
rect 592382 286398 592618 286634
rect 592062 250718 592298 250954
rect 592382 250718 592618 250954
rect 592062 250398 592298 250634
rect 592382 250398 592618 250634
rect 592062 214718 592298 214954
rect 592382 214718 592618 214954
rect 592062 214398 592298 214634
rect 592382 214398 592618 214634
rect 592062 178718 592298 178954
rect 592382 178718 592618 178954
rect 592062 178398 592298 178634
rect 592382 178398 592618 178634
rect 592062 142718 592298 142954
rect 592382 142718 592618 142954
rect 592062 142398 592298 142634
rect 592382 142398 592618 142634
rect 592062 106718 592298 106954
rect 592382 106718 592618 106954
rect 592062 106398 592298 106634
rect 592382 106398 592618 106634
rect 592062 70718 592298 70954
rect 592382 70718 592618 70954
rect 592062 70398 592298 70634
rect 592382 70398 592618 70634
rect 592062 34718 592298 34954
rect 592382 34718 592618 34954
rect 592062 34398 592298 34634
rect 592382 34398 592618 34634
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 700954 592650 700986
rect -8726 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 592650 700954
rect -8726 700634 592650 700718
rect -8726 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 592650 700634
rect -8726 700366 592650 700398
rect -8726 696454 592650 696486
rect -8726 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 592650 696454
rect -8726 696134 592650 696218
rect -8726 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 592650 696134
rect -8726 695866 592650 695898
rect -8726 691954 592650 691986
rect -8726 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 592650 691954
rect -8726 691634 592650 691718
rect -8726 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 592650 691634
rect -8726 691366 592650 691398
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 682954 592650 682986
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect -8726 682634 592650 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect -8726 682366 592650 682398
rect -8726 678454 592650 678486
rect -8726 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 592650 678454
rect -8726 678134 592650 678218
rect -8726 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 592650 678134
rect -8726 677866 592650 677898
rect -8726 673954 592650 673986
rect -8726 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 592650 673954
rect -8726 673634 592650 673718
rect -8726 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 592650 673634
rect -8726 673366 592650 673398
rect -8726 669454 592650 669486
rect -8726 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 592650 669454
rect -8726 669134 592650 669218
rect -8726 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 592650 669134
rect -8726 668866 592650 668898
rect -8726 664954 592650 664986
rect -8726 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 592650 664954
rect -8726 664634 592650 664718
rect -8726 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 592650 664634
rect -8726 664366 592650 664398
rect -8726 660454 592650 660486
rect -8726 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 592650 660454
rect -8726 660134 592650 660218
rect -8726 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 592650 660134
rect -8726 659866 592650 659898
rect -8726 655954 592650 655986
rect -8726 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 592650 655954
rect -8726 655634 592650 655718
rect -8726 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 592650 655634
rect -8726 655366 592650 655398
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 646954 592650 646986
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect -8726 646634 592650 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect -8726 646366 592650 646398
rect -8726 642454 592650 642486
rect -8726 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 592650 642454
rect -8726 642134 592650 642218
rect -8726 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 592650 642134
rect -8726 641866 592650 641898
rect -8726 637954 592650 637986
rect -8726 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 592650 637954
rect -8726 637634 592650 637718
rect -8726 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 592650 637634
rect -8726 637366 592650 637398
rect -8726 633454 592650 633486
rect -8726 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 592650 633454
rect -8726 633134 592650 633218
rect -8726 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 592650 633134
rect -8726 632866 592650 632898
rect -8726 628954 592650 628986
rect -8726 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 592650 628954
rect -8726 628634 592650 628718
rect -8726 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 592650 628634
rect -8726 628366 592650 628398
rect -8726 624454 592650 624486
rect -8726 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 592650 624454
rect -8726 624134 592650 624218
rect -8726 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 592650 624134
rect -8726 623866 592650 623898
rect -8726 619954 592650 619986
rect -8726 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 592650 619954
rect -8726 619634 592650 619718
rect -8726 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 592650 619634
rect -8726 619366 592650 619398
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 610954 592650 610986
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect -8726 610634 592650 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect -8726 610366 592650 610398
rect -8726 606454 592650 606486
rect -8726 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 592650 606454
rect -8726 606134 592650 606218
rect -8726 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 592650 606134
rect -8726 605866 592650 605898
rect -8726 601954 592650 601986
rect -8726 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 592650 601954
rect -8726 601634 592650 601718
rect -8726 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 592650 601634
rect -8726 601366 592650 601398
rect -8726 597454 592650 597486
rect -8726 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 592650 597454
rect -8726 597134 592650 597218
rect -8726 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 592650 597134
rect -8726 596866 592650 596898
rect -8726 592954 592650 592986
rect -8726 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 592650 592954
rect -8726 592634 592650 592718
rect -8726 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 592650 592634
rect -8726 592366 592650 592398
rect -8726 588454 592650 588486
rect -8726 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 592650 588454
rect -8726 588134 592650 588218
rect -8726 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 592650 588134
rect -8726 587866 592650 587898
rect -8726 583954 592650 583986
rect -8726 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 592650 583954
rect -8726 583634 592650 583718
rect -8726 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 592650 583634
rect -8726 583366 592650 583398
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 574954 592650 574986
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect -8726 574634 592650 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect -8726 574366 592650 574398
rect -8726 570454 592650 570486
rect -8726 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 592650 570454
rect -8726 570134 592650 570218
rect -8726 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 592650 570134
rect -8726 569866 592650 569898
rect -8726 565954 592650 565986
rect -8726 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 592650 565954
rect -8726 565634 592650 565718
rect -8726 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 592650 565634
rect -8726 565366 592650 565398
rect -8726 561454 592650 561486
rect -8726 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 592650 561454
rect -8726 561134 592650 561218
rect -8726 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 592650 561134
rect -8726 560866 592650 560898
rect -8726 556954 592650 556986
rect -8726 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 592650 556954
rect -8726 556634 592650 556718
rect -8726 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 592650 556634
rect -8726 556366 592650 556398
rect -8726 552454 592650 552486
rect -8726 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 592650 552454
rect -8726 552134 592650 552218
rect -8726 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 592650 552134
rect -8726 551866 592650 551898
rect -8726 547954 592650 547986
rect -8726 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 592650 547954
rect -8726 547634 592650 547718
rect -8726 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 592650 547634
rect -8726 547366 592650 547398
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 538954 592650 538986
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect -8726 538634 592650 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect -8726 538366 592650 538398
rect -8726 534454 592650 534486
rect -8726 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 592650 534454
rect -8726 534134 592650 534218
rect -8726 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 592650 534134
rect -8726 533866 592650 533898
rect -8726 529954 592650 529986
rect -8726 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 592650 529954
rect -8726 529634 592650 529718
rect -8726 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 592650 529634
rect -8726 529366 592650 529398
rect -8726 525454 592650 525486
rect -8726 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 592650 525454
rect -8726 525134 592650 525218
rect -8726 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 592650 525134
rect -8726 524866 592650 524898
rect -8726 520954 592650 520986
rect -8726 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 592650 520954
rect -8726 520634 592650 520718
rect -8726 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 592650 520634
rect -8726 520366 592650 520398
rect -8726 516454 592650 516486
rect -8726 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 592650 516454
rect -8726 516134 592650 516218
rect -8726 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 592650 516134
rect -8726 515866 592650 515898
rect -8726 511954 592650 511986
rect -8726 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 592650 511954
rect -8726 511634 592650 511718
rect -8726 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 592650 511634
rect -8726 511366 592650 511398
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 502954 592650 502986
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect -8726 502634 592650 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect -8726 502366 592650 502398
rect -8726 498454 592650 498486
rect -8726 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 592650 498454
rect -8726 498134 592650 498218
rect -8726 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 592650 498134
rect -8726 497866 592650 497898
rect -8726 493954 592650 493986
rect -8726 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 592650 493954
rect -8726 493634 592650 493718
rect -8726 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 592650 493634
rect -8726 493366 592650 493398
rect -8726 489454 592650 489486
rect -8726 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 592650 489454
rect -8726 489134 592650 489218
rect -8726 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 592650 489134
rect -8726 488866 592650 488898
rect -8726 484954 592650 484986
rect -8726 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 592650 484954
rect -8726 484634 592650 484718
rect -8726 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 592650 484634
rect -8726 484366 592650 484398
rect -8726 480454 592650 480486
rect -8726 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 592650 480454
rect -8726 480134 592650 480218
rect -8726 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 592650 480134
rect -8726 479866 592650 479898
rect -8726 475954 592650 475986
rect -8726 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 592650 475954
rect -8726 475634 592650 475718
rect -8726 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 592650 475634
rect -8726 475366 592650 475398
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 466954 592650 466986
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect -8726 466634 592650 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect -8726 466366 592650 466398
rect -8726 462454 592650 462486
rect -8726 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 592650 462454
rect -8726 462134 592650 462218
rect -8726 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 592650 462134
rect -8726 461866 592650 461898
rect -8726 457954 592650 457986
rect -8726 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 592650 457954
rect -8726 457634 592650 457718
rect -8726 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 592650 457634
rect -8726 457366 592650 457398
rect -8726 453454 592650 453486
rect -8726 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 592650 453454
rect -8726 453134 592650 453218
rect -8726 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 592650 453134
rect -8726 452866 592650 452898
rect -8726 448954 592650 448986
rect -8726 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 592650 448954
rect -8726 448634 592650 448718
rect -8726 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 592650 448634
rect -8726 448366 592650 448398
rect -8726 444454 592650 444486
rect -8726 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 592650 444454
rect -8726 444134 592650 444218
rect -8726 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 592650 444134
rect -8726 443866 592650 443898
rect -8726 439954 592650 439986
rect -8726 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 592650 439954
rect -8726 439634 592650 439718
rect -8726 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 592650 439634
rect -8726 439366 592650 439398
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 430954 592650 430986
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect -8726 430634 592650 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect -8726 430366 592650 430398
rect -8726 426454 592650 426486
rect -8726 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 592650 426454
rect -8726 426134 592650 426218
rect -8726 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 592650 426134
rect -8726 425866 592650 425898
rect -8726 421954 592650 421986
rect -8726 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 592650 421954
rect -8726 421634 592650 421718
rect -8726 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 592650 421634
rect -8726 421366 592650 421398
rect -8726 417454 592650 417486
rect -8726 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 592650 417454
rect -8726 417134 592650 417218
rect -8726 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 592650 417134
rect -8726 416866 592650 416898
rect -8726 412954 592650 412986
rect -8726 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 592650 412954
rect -8726 412634 592650 412718
rect -8726 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 592650 412634
rect -8726 412366 592650 412398
rect -8726 408454 592650 408486
rect -8726 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 592650 408454
rect -8726 408134 592650 408218
rect -8726 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 592650 408134
rect -8726 407866 592650 407898
rect -8726 403954 592650 403986
rect -8726 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 592650 403954
rect -8726 403634 592650 403718
rect -8726 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 592650 403634
rect -8726 403366 592650 403398
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 394954 592650 394986
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect -8726 394634 592650 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect -8726 394366 592650 394398
rect -8726 390454 592650 390486
rect -8726 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 592650 390454
rect -8726 390134 592650 390218
rect -8726 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 592650 390134
rect -8726 389866 592650 389898
rect -8726 385954 592650 385986
rect -8726 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 592650 385954
rect -8726 385634 592650 385718
rect -8726 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 592650 385634
rect -8726 385366 592650 385398
rect -8726 381454 592650 381486
rect -8726 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 592650 381454
rect -8726 381134 592650 381218
rect -8726 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 592650 381134
rect -8726 380866 592650 380898
rect -8726 376954 592650 376986
rect -8726 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 592650 376954
rect -8726 376634 592650 376718
rect -8726 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 592650 376634
rect -8726 376366 592650 376398
rect -8726 372454 592650 372486
rect -8726 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 592650 372454
rect -8726 372134 592650 372218
rect -8726 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 592650 372134
rect -8726 371866 592650 371898
rect -8726 367954 592650 367986
rect -8726 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 592650 367954
rect -8726 367634 592650 367718
rect -8726 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 592650 367634
rect -8726 367366 592650 367398
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 358954 592650 358986
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect -8726 358634 592650 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect -8726 358366 592650 358398
rect -8726 354454 592650 354486
rect -8726 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 244826 354454
rect 245062 354218 245146 354454
rect 245382 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 592650 354454
rect -8726 354134 592650 354218
rect -8726 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 244826 354134
rect 245062 353898 245146 354134
rect 245382 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 592650 354134
rect -8726 353866 592650 353898
rect -8726 349954 592650 349986
rect -8726 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 240326 349954
rect 240562 349718 240646 349954
rect 240882 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 592650 349954
rect -8726 349634 592650 349718
rect -8726 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 240326 349634
rect 240562 349398 240646 349634
rect 240882 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 592650 349634
rect -8726 349366 592650 349398
rect -8726 345454 592650 345486
rect -8726 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 592650 345454
rect -8726 345134 592650 345218
rect -8726 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 592650 345134
rect -8726 344866 592650 344898
rect -8726 340954 592650 340986
rect -8726 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 592650 340954
rect -8726 340634 592650 340718
rect -8726 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 592650 340634
rect -8726 340366 592650 340398
rect -8726 336454 592650 336486
rect -8726 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 592650 336454
rect -8726 336134 592650 336218
rect -8726 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 592650 336134
rect -8726 335866 592650 335898
rect -8726 331954 592650 331986
rect -8726 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 592650 331954
rect -8726 331634 592650 331718
rect -8726 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 592650 331634
rect -8726 331366 592650 331398
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 322954 592650 322986
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect -8726 322634 592650 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect -8726 322366 592650 322398
rect -8726 318454 592650 318486
rect -8726 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 592650 318454
rect -8726 318134 592650 318218
rect -8726 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 592650 318134
rect -8726 317866 592650 317898
rect -8726 313954 592650 313986
rect -8726 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 592650 313954
rect -8726 313634 592650 313718
rect -8726 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 592650 313634
rect -8726 313366 592650 313398
rect -8726 309454 592650 309486
rect -8726 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 592650 309454
rect -8726 309134 592650 309218
rect -8726 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 592650 309134
rect -8726 308866 592650 308898
rect -8726 304954 592650 304986
rect -8726 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 592650 304954
rect -8726 304634 592650 304718
rect -8726 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 592650 304634
rect -8726 304366 592650 304398
rect -8726 300454 592650 300486
rect -8726 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 592650 300454
rect -8726 300134 592650 300218
rect -8726 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 592650 300134
rect -8726 299866 592650 299898
rect -8726 295954 592650 295986
rect -8726 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 592650 295954
rect -8726 295634 592650 295718
rect -8726 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 592650 295634
rect -8726 295366 592650 295398
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 286954 592650 286986
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect -8726 286634 592650 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect -8726 286366 592650 286398
rect -8726 282454 592650 282486
rect -8726 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 592650 282454
rect -8726 282134 592650 282218
rect -8726 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 592650 282134
rect -8726 281866 592650 281898
rect -8726 277954 592650 277986
rect -8726 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 592650 277954
rect -8726 277634 592650 277718
rect -8726 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 592650 277634
rect -8726 277366 592650 277398
rect -8726 273454 592650 273486
rect -8726 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 592650 273454
rect -8726 273134 592650 273218
rect -8726 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 592650 273134
rect -8726 272866 592650 272898
rect -8726 268954 592650 268986
rect -8726 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 592650 268954
rect -8726 268634 592650 268718
rect -8726 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 592650 268634
rect -8726 268366 592650 268398
rect -8726 264454 592650 264486
rect -8726 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 592650 264454
rect -8726 264134 592650 264218
rect -8726 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 592650 264134
rect -8726 263866 592650 263898
rect -8726 259954 592650 259986
rect -8726 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 592650 259954
rect -8726 259634 592650 259718
rect -8726 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 592650 259634
rect -8726 259366 592650 259398
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 250954 592650 250986
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect -8726 250634 592650 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect -8726 250366 592650 250398
rect -8726 246454 592650 246486
rect -8726 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246303 424826 246454
rect 29382 246218 65342 246303
rect -8726 246134 65342 246218
rect -8726 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 246067 65342 246134
rect 65578 246067 65662 246303
rect 65898 246067 65982 246303
rect 66218 246067 66302 246303
rect 66538 246067 66622 246303
rect 66858 246067 66942 246303
rect 67178 246067 67262 246303
rect 67498 246067 67582 246303
rect 67818 246067 67902 246303
rect 68138 246067 68222 246303
rect 68458 246067 68542 246303
rect 68778 246067 68862 246303
rect 69098 246067 69182 246303
rect 69418 246067 69502 246303
rect 69738 246067 69822 246303
rect 70058 246218 424826 246303
rect 425062 246218 425146 246454
rect 425382 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 592650 246454
rect 70058 246134 592650 246218
rect 70058 246067 424826 246134
rect 29382 245898 424826 246067
rect 425062 245898 425146 246134
rect 425382 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 592650 246134
rect -8726 245866 592650 245898
rect -8726 241954 592650 241986
rect -8726 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241953 420326 241954
rect 24882 241718 65462 241953
rect -8726 241717 65462 241718
rect 65698 241717 65782 241953
rect 66018 241717 66102 241953
rect 66338 241717 66422 241953
rect 66658 241717 66742 241953
rect 66978 241717 67062 241953
rect 67298 241717 67382 241953
rect 67618 241717 67702 241953
rect 67938 241717 68022 241953
rect 68258 241717 68342 241953
rect 68578 241717 68662 241953
rect 68898 241717 68982 241953
rect 69218 241717 69302 241953
rect 69538 241717 69622 241953
rect 69858 241717 69942 241953
rect 70178 241717 70262 241953
rect 70498 241717 70582 241953
rect 70818 241717 70902 241953
rect 71138 241718 420326 241953
rect 420562 241718 420646 241954
rect 420882 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 592650 241954
rect 71138 241717 592650 241718
rect -8726 241634 592650 241717
rect -8726 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241633 420326 241634
rect 24882 241398 65462 241633
rect -8726 241397 65462 241398
rect 65698 241397 65782 241633
rect 66018 241397 66102 241633
rect 66338 241397 66422 241633
rect 66658 241397 66742 241633
rect 66978 241397 67062 241633
rect 67298 241397 67382 241633
rect 67618 241397 67702 241633
rect 67938 241397 68022 241633
rect 68258 241397 68342 241633
rect 68578 241397 68662 241633
rect 68898 241397 68982 241633
rect 69218 241397 69302 241633
rect 69538 241397 69622 241633
rect 69858 241397 69942 241633
rect 70178 241397 70262 241633
rect 70498 241397 70582 241633
rect 70818 241397 70902 241633
rect 71138 241398 420326 241633
rect 420562 241398 420646 241634
rect 420882 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 592650 241634
rect 71138 241397 592650 241398
rect -8726 241366 592650 241397
rect -8726 237454 592650 237486
rect -8726 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 592650 237454
rect -8726 237134 592650 237218
rect -8726 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 592650 237134
rect -8726 236866 592650 236898
rect -8726 232954 592650 232986
rect -8726 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 592650 232954
rect -8726 232634 592650 232718
rect -8726 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 592650 232634
rect -8726 232366 592650 232398
rect -8726 228454 592650 228486
rect -8726 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228453 406826 228454
rect 11382 228218 46826 228453
rect -8726 228217 46826 228218
rect 47062 228217 47146 228453
rect 47382 228217 82826 228453
rect 83062 228217 83146 228453
rect 83382 228217 118826 228453
rect 119062 228217 119146 228453
rect 119382 228217 190826 228453
rect 191062 228217 191146 228453
rect 191382 228217 226826 228453
rect 227062 228217 227146 228453
rect 227382 228217 262826 228453
rect 263062 228217 263146 228453
rect 263382 228217 298826 228453
rect 299062 228217 299146 228453
rect 299382 228217 334826 228453
rect 335062 228217 335146 228453
rect 335382 228217 370826 228453
rect 371062 228217 371146 228453
rect 371382 228218 406826 228453
rect 407062 228218 407146 228454
rect 407382 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 592650 228454
rect 371382 228217 592650 228218
rect -8726 228134 592650 228217
rect -8726 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 228133 406826 228134
rect 11382 227898 46826 228133
rect -8726 227897 46826 227898
rect 47062 227897 47146 228133
rect 47382 227897 82826 228133
rect 83062 227897 83146 228133
rect 83382 227897 118826 228133
rect 119062 227897 119146 228133
rect 119382 227897 190826 228133
rect 191062 227897 191146 228133
rect 191382 227897 226826 228133
rect 227062 227897 227146 228133
rect 227382 227897 262826 228133
rect 263062 227897 263146 228133
rect 263382 227897 298826 228133
rect 299062 227897 299146 228133
rect 299382 227897 334826 228133
rect 335062 227897 335146 228133
rect 335382 227897 370826 228133
rect 371062 227897 371146 228133
rect 371382 227898 406826 228133
rect 407062 227898 407146 228134
rect 407382 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 592650 228134
rect 371382 227897 592650 227898
rect -8726 227866 592650 227897
rect -8726 223954 592650 223986
rect -8726 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 592650 223954
rect -8726 223634 592650 223718
rect -8726 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 592650 223634
rect -8726 223366 592650 223398
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 214954 592650 214986
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect -8726 214634 592650 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect -8726 214366 592650 214398
rect -8726 210454 592650 210486
rect -8726 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 592650 210454
rect -8726 210134 592650 210218
rect -8726 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 592650 210134
rect -8726 209866 592650 209898
rect -8726 205954 592650 205986
rect -8726 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205861 204326 205954
rect 132882 205718 136036 205861
rect -8726 205634 136036 205718
rect -8726 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205625 136036 205634
rect 136272 205625 136356 205861
rect 136592 205625 136676 205861
rect 136912 205625 136996 205861
rect 137232 205625 137316 205861
rect 137552 205625 137636 205861
rect 137872 205625 137956 205861
rect 138192 205625 138276 205861
rect 138512 205625 138596 205861
rect 138832 205625 138916 205861
rect 139152 205625 139236 205861
rect 139472 205625 139556 205861
rect 139792 205625 139876 205861
rect 140112 205625 140196 205861
rect 140432 205625 140516 205861
rect 140752 205625 140836 205861
rect 141072 205625 141156 205861
rect 141392 205625 141476 205861
rect 141712 205625 141796 205861
rect 142032 205625 142116 205861
rect 142352 205625 142436 205861
rect 142672 205625 142756 205861
rect 142992 205625 143076 205861
rect 143312 205625 143396 205861
rect 143632 205625 143716 205861
rect 143952 205625 144036 205861
rect 144272 205625 144356 205861
rect 144592 205625 144676 205861
rect 144912 205625 144996 205861
rect 145232 205625 145316 205861
rect 145552 205625 145636 205861
rect 145872 205625 145956 205861
rect 146192 205625 146276 205861
rect 146512 205625 146596 205861
rect 146832 205625 146916 205861
rect 147152 205625 147236 205861
rect 147472 205625 147556 205861
rect 147792 205625 147876 205861
rect 148112 205625 148196 205861
rect 148432 205625 148516 205861
rect 148752 205625 148836 205861
rect 149072 205625 149156 205861
rect 149392 205625 149476 205861
rect 149712 205625 149796 205861
rect 150032 205625 150116 205861
rect 150352 205625 150436 205861
rect 150672 205625 150756 205861
rect 150992 205625 151076 205861
rect 151312 205625 151396 205861
rect 151632 205625 151716 205861
rect 151952 205625 152036 205861
rect 152272 205625 152356 205861
rect 152592 205625 152676 205861
rect 152912 205625 152996 205861
rect 153232 205625 153316 205861
rect 153552 205625 153636 205861
rect 153872 205625 153956 205861
rect 154192 205625 154276 205861
rect 154512 205625 154596 205861
rect 154832 205625 154916 205861
rect 155152 205625 155236 205861
rect 155472 205625 155556 205861
rect 155792 205625 155876 205861
rect 156112 205625 156196 205861
rect 156432 205625 156516 205861
rect 156752 205625 156836 205861
rect 157072 205625 157156 205861
rect 157392 205625 157476 205861
rect 157712 205625 157796 205861
rect 158032 205625 158116 205861
rect 158352 205625 158436 205861
rect 158672 205625 158756 205861
rect 158992 205625 159076 205861
rect 159312 205625 159396 205861
rect 159632 205625 159716 205861
rect 159952 205625 160036 205861
rect 160272 205625 160356 205861
rect 160592 205625 160676 205861
rect 160912 205625 160996 205861
rect 161232 205625 161316 205861
rect 161552 205625 161636 205861
rect 161872 205625 161956 205861
rect 162192 205625 162276 205861
rect 162512 205625 162596 205861
rect 162832 205625 162916 205861
rect 163152 205625 163236 205861
rect 163472 205625 163556 205861
rect 163792 205625 163876 205861
rect 164112 205625 164196 205861
rect 164432 205625 164516 205861
rect 164752 205625 164836 205861
rect 165072 205625 165156 205861
rect 165392 205718 204326 205861
rect 204562 205718 204646 205954
rect 204882 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 592650 205954
rect 165392 205634 592650 205718
rect 165392 205625 204326 205634
rect 132882 205398 204326 205625
rect 204562 205398 204646 205634
rect 204882 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 592650 205634
rect -8726 205366 592650 205398
rect -8726 201454 592650 201486
rect -8726 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201411 199826 201454
rect 128382 201218 137376 201411
rect -8726 201175 137376 201218
rect 137612 201175 137696 201411
rect 137932 201175 138016 201411
rect 138252 201175 138336 201411
rect 138572 201175 138656 201411
rect 138892 201175 138976 201411
rect 139212 201175 139296 201411
rect 139532 201175 139616 201411
rect 139852 201175 139936 201411
rect 140172 201175 140256 201411
rect 140492 201175 140576 201411
rect 140812 201175 140896 201411
rect 141132 201175 141216 201411
rect 141452 201175 141536 201411
rect 141772 201175 141856 201411
rect 142092 201175 142176 201411
rect 142412 201175 142496 201411
rect 142732 201175 142816 201411
rect 143052 201175 143136 201411
rect 143372 201175 143456 201411
rect 143692 201175 143776 201411
rect 144012 201175 144096 201411
rect 144332 201175 144416 201411
rect 144652 201175 144736 201411
rect 144972 201175 145056 201411
rect 145292 201175 145376 201411
rect 145612 201175 145696 201411
rect 145932 201175 146016 201411
rect 146252 201175 146336 201411
rect 146572 201175 146656 201411
rect 146892 201175 146976 201411
rect 147212 201175 147296 201411
rect 147532 201175 147616 201411
rect 147852 201175 147936 201411
rect 148172 201175 148256 201411
rect 148492 201175 148576 201411
rect 148812 201175 148896 201411
rect 149132 201175 149216 201411
rect 149452 201175 149536 201411
rect 149772 201175 149856 201411
rect 150092 201175 150176 201411
rect 150412 201175 150496 201411
rect 150732 201175 150816 201411
rect 151052 201175 151136 201411
rect 151372 201175 151456 201411
rect 151692 201175 151776 201411
rect 152012 201175 152096 201411
rect 152332 201175 152416 201411
rect 152652 201175 152736 201411
rect 152972 201175 153056 201411
rect 153292 201175 153376 201411
rect 153612 201175 153696 201411
rect 153932 201175 154016 201411
rect 154252 201175 154336 201411
rect 154572 201175 154656 201411
rect 154892 201175 154976 201411
rect 155212 201175 155296 201411
rect 155532 201175 155616 201411
rect 155852 201175 155936 201411
rect 156172 201175 156256 201411
rect 156492 201175 156576 201411
rect 156812 201175 156896 201411
rect 157132 201175 157216 201411
rect 157452 201175 157536 201411
rect 157772 201175 157856 201411
rect 158092 201175 158176 201411
rect 158412 201175 158496 201411
rect 158732 201175 158816 201411
rect 159052 201175 159136 201411
rect 159372 201175 159456 201411
rect 159692 201175 159776 201411
rect 160012 201175 160096 201411
rect 160332 201175 160416 201411
rect 160652 201175 160736 201411
rect 160972 201175 161056 201411
rect 161292 201175 161376 201411
rect 161612 201175 161696 201411
rect 161932 201175 162016 201411
rect 162252 201175 162336 201411
rect 162572 201175 162656 201411
rect 162892 201175 162976 201411
rect 163212 201175 163296 201411
rect 163532 201175 163616 201411
rect 163852 201175 163936 201411
rect 164172 201175 164256 201411
rect 164492 201175 164576 201411
rect 164812 201175 164896 201411
rect 165132 201175 165216 201411
rect 165452 201218 199826 201411
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 592650 201454
rect 165452 201175 592650 201218
rect -8726 201134 592650 201175
rect -8726 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 592650 201134
rect -8726 200866 592650 200898
rect -8726 196954 592650 196986
rect -8726 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 592650 196954
rect -8726 196634 592650 196718
rect -8726 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 592650 196634
rect -8726 196366 592650 196398
rect -8726 192454 592650 192486
rect -8726 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 592650 192454
rect -8726 192134 592650 192218
rect -8726 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 592650 192134
rect -8726 191866 592650 191898
rect -8726 187954 592650 187986
rect -8726 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 592650 187954
rect -8726 187634 592650 187718
rect -8726 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 592650 187634
rect -8726 187366 592650 187398
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 178954 592650 178986
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect -8726 178634 592650 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect -8726 178366 592650 178398
rect -8726 174454 592650 174486
rect -8726 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 137066 174454
rect 137302 174218 137386 174454
rect 137622 174218 137706 174454
rect 137942 174218 138026 174454
rect 138262 174218 138346 174454
rect 138582 174218 138666 174454
rect 138902 174218 138986 174454
rect 139222 174218 139306 174454
rect 139542 174218 139626 174454
rect 139862 174218 139946 174454
rect 140182 174218 140266 174454
rect 140502 174218 140586 174454
rect 140822 174218 140906 174454
rect 141142 174218 141226 174454
rect 141462 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 316826 174454
rect 317062 174218 317146 174454
rect 317382 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 592650 174454
rect -8726 174134 592650 174218
rect -8726 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 137066 174134
rect 137302 173898 137386 174134
rect 137622 173898 137706 174134
rect 137942 173898 138026 174134
rect 138262 173898 138346 174134
rect 138582 173898 138666 174134
rect 138902 173898 138986 174134
rect 139222 173898 139306 174134
rect 139542 173898 139626 174134
rect 139862 173898 139946 174134
rect 140182 173898 140266 174134
rect 140502 173898 140586 174134
rect 140822 173898 140906 174134
rect 141142 173898 141226 174134
rect 141462 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 316826 174134
rect 317062 173898 317146 174134
rect 317382 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 592650 174134
rect -8726 173866 592650 173898
rect -8726 169954 592650 169986
rect -8726 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 132326 169954
rect 132562 169718 132646 169954
rect 132882 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 312326 169954
rect 312562 169718 312646 169954
rect 312882 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 592650 169954
rect -8726 169634 592650 169718
rect -8726 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 132326 169634
rect 132562 169398 132646 169634
rect 132882 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 312326 169634
rect 312562 169398 312646 169634
rect 312882 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 592650 169634
rect -8726 169366 592650 169398
rect -8726 165454 592650 165486
rect -8726 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 592650 165454
rect -8726 165134 592650 165218
rect -8726 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 592650 165134
rect -8726 164866 592650 164898
rect -8726 160954 592650 160986
rect -8726 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 592650 160954
rect -8726 160634 592650 160718
rect -8726 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 592650 160634
rect -8726 160366 592650 160398
rect -8726 156454 592650 156486
rect -8726 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 592650 156454
rect -8726 156134 592650 156218
rect -8726 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 592650 156134
rect -8726 155866 592650 155898
rect -8726 151954 592650 151986
rect -8726 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 592650 151954
rect -8726 151634 592650 151718
rect -8726 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 592650 151634
rect -8726 151366 592650 151398
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 142954 592650 142986
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect -8726 142634 592650 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect -8726 142366 592650 142398
rect -8726 138454 592650 138486
rect -8726 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 172826 138454
rect 173062 138218 173146 138454
rect 173382 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 592650 138454
rect -8726 138134 592650 138218
rect -8726 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 172826 138134
rect 173062 137898 173146 138134
rect 173382 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 592650 138134
rect -8726 137866 592650 137898
rect -8726 133954 592650 133986
rect -8726 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 592650 133954
rect -8726 133634 592650 133718
rect -8726 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 592650 133634
rect -8726 133366 592650 133398
rect -8726 129454 592650 129486
rect -8726 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 592650 129454
rect -8726 129134 592650 129218
rect -8726 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 592650 129134
rect -8726 128866 592650 128898
rect -8726 124954 592650 124986
rect -8726 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 592650 124954
rect -8726 124634 592650 124718
rect -8726 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 592650 124634
rect -8726 124366 592650 124398
rect -8726 120454 592650 120486
rect -8726 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 592650 120454
rect -8726 120134 592650 120218
rect -8726 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 592650 120134
rect -8726 119866 592650 119898
rect -8726 115954 592650 115986
rect -8726 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 135610 115954
rect 135846 115718 166330 115954
rect 166566 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 592650 115954
rect -8726 115634 592650 115718
rect -8726 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 135610 115634
rect 135846 115398 166330 115634
rect 166566 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 592650 115634
rect -8726 115366 592650 115398
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 120250 111454
rect 120486 111218 150970 111454
rect 151206 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 120250 111134
rect 120486 110898 150970 111134
rect 151206 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 106954 592650 106986
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect -8726 106634 592650 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect -8726 106366 592650 106398
rect -8726 102454 592650 102486
rect -8726 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 592650 102454
rect -8726 102134 592650 102218
rect -8726 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 592650 102134
rect -8726 101866 592650 101898
rect -8726 97954 592650 97986
rect -8726 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 592650 97954
rect -8726 97634 592650 97718
rect -8726 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 592650 97634
rect -8726 97366 592650 97398
rect -8726 93454 592650 93486
rect -8726 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 592650 93454
rect -8726 93134 592650 93218
rect -8726 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 592650 93134
rect -8726 92866 592650 92898
rect -8726 88954 592650 88986
rect -8726 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 592650 88954
rect -8726 88634 592650 88718
rect -8726 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 592650 88634
rect -8726 88366 592650 88398
rect -8726 84454 592650 84486
rect -8726 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 592650 84454
rect -8726 84134 592650 84218
rect -8726 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 592650 84134
rect -8726 83866 592650 83898
rect -8726 79954 592650 79986
rect -8726 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 135610 79954
rect 135846 79718 166330 79954
rect 166566 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 592650 79954
rect -8726 79634 592650 79718
rect -8726 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 135610 79634
rect 135846 79398 166330 79634
rect 166566 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 592650 79634
rect -8726 79366 592650 79398
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 70954 592650 70986
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect -8726 70634 592650 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect -8726 70366 592650 70398
rect -8726 66454 592650 66486
rect -8726 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 592650 66454
rect -8726 66134 592650 66218
rect -8726 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 592650 66134
rect -8726 65866 592650 65898
rect -8726 61954 592650 61986
rect -8726 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 592650 61954
rect -8726 61634 592650 61718
rect -8726 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 592650 61634
rect -8726 61366 592650 61398
rect -8726 57454 592650 57486
rect -8726 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 592650 57454
rect -8726 57134 592650 57218
rect -8726 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 592650 57134
rect -8726 56866 592650 56898
rect -8726 52954 592650 52986
rect -8726 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 592650 52954
rect -8726 52634 592650 52718
rect -8726 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 592650 52634
rect -8726 52366 592650 52398
rect -8726 48454 592650 48486
rect -8726 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 592650 48454
rect -8726 48134 592650 48218
rect -8726 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 592650 48134
rect -8726 47866 592650 47898
rect -8726 43954 592650 43986
rect -8726 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 592650 43954
rect -8726 43634 592650 43718
rect -8726 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 592650 43634
rect -8726 43366 592650 43398
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 34954 592650 34986
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect -8726 34634 592650 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect -8726 34366 592650 34398
rect -8726 30454 592650 30486
rect -8726 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 592650 30454
rect -8726 30134 592650 30218
rect -8726 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 592650 30134
rect -8726 29866 592650 29898
rect -8726 25954 592650 25986
rect -8726 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 592650 25954
rect -8726 25634 592650 25718
rect -8726 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 592650 25634
rect -8726 25366 592650 25398
rect -8726 21454 592650 21486
rect -8726 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 592650 21454
rect -8726 21134 592650 21218
rect -8726 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 592650 21134
rect -8726 20866 592650 20898
rect -8726 16954 592650 16986
rect -8726 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 592650 16954
rect -8726 16634 592650 16718
rect -8726 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 592650 16634
rect -8726 16366 592650 16398
rect -8726 12454 592650 12486
rect -8726 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 592650 12454
rect -8726 12134 592650 12218
rect -8726 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 592650 12134
rect -8726 11866 592650 11898
rect -8726 7954 592650 7986
rect -8726 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 592650 7954
rect -8726 7634 592650 7718
rect -8726 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 592650 7634
rect -8726 7366 592650 7398
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use PD_M1_M2  PD_M1_M2_macro0
timestamp 0
transform 1 0 16000 0 1 232484
box 30000 -2000 380500 14200
use rlbp_macro  rlbp_macro0
timestamp 0
transform 1 0 116000 0 1 75000
box 0 0 60000 60000
use SystemLevel  sl_macro0
timestamp 0
transform 1 0 148914 0 1 188300
box -13000 -15200 17500 18000
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 248684 74414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 248684 110414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 73000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 248684 146414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 248684 182414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 248684 218414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 248684 254414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 248684 290414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 248684 326414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 248684 362414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 248684 398414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 10794 -7654 11414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 46794 -7654 47414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 46794 248684 47414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 -7654 83414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 248684 83414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 -7654 119414 73000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 137000 119414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 248684 119414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 -7654 155414 73000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 248684 155414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 -7654 191414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 248684 191414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 -7654 227414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 248684 227414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 -7654 263414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 248684 263414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 -7654 299414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 248684 299414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 -7654 335414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 248684 335414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 -7654 371414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 248684 371414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 406794 -7654 407414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 442794 -7654 443414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 478794 -7654 479414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 514794 -7654 515414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 550794 -7654 551414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 11866 592650 12486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 47866 592650 48486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 83866 592650 84486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 119866 592650 120486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 155866 592650 156486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 191866 592650 192486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 227866 592650 228486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 263866 592650 264486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 299866 592650 300486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 335866 592650 336486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 371866 592650 372486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 407866 592650 408486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 443866 592650 444486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 479866 592650 480486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 515866 592650 516486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 551866 592650 552486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 587866 592650 588486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 623866 592650 624486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 659866 592650 660486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 695866 592650 696486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 19794 -7654 20414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 55794 -7654 56414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 55794 248684 56414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 -7654 92414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 248684 92414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 -7654 128414 73000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 137000 128414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 248684 128414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 -7654 164414 73000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 248684 164414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 -7654 200414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 248684 200414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 -7654 236414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 248684 236414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 271794 -7654 272414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 271794 248684 272414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 -7654 308414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 248684 308414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 343794 -7654 344414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 343794 248684 344414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 -7654 380414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 248684 380414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 415794 -7654 416414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 451794 -7654 452414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 487794 -7654 488414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 523794 -7654 524414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 559794 -7654 560414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 20866 592650 21486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 56866 592650 57486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 92866 592650 93486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 128866 592650 129486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 164866 592650 165486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 200866 592650 201486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 236866 592650 237486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 272866 592650 273486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 308866 592650 309486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 344866 592650 345486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 380866 592650 381486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 416866 592650 417486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 452866 592650 453486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 488866 592650 489486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 524866 592650 525486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 560866 592650 561486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 596866 592650 597486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 632866 592650 633486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 668866 592650 669486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 28794 -7654 29414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 64794 -7654 65414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 64794 248684 65414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 100794 -7654 101414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 100794 248684 101414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 -7654 137414 73000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 248684 137414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 -7654 173414 73000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 137000 173414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 248684 173414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 208794 -7654 209414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 208794 248684 209414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 244794 -7654 245414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 244794 248684 245414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 280794 -7654 281414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 280794 248684 281414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 316794 -7654 317414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 316794 248684 317414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 352794 -7654 353414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 352794 248684 353414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 388794 -7654 389414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 388794 248684 389414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 424794 -7654 425414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 460794 -7654 461414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 496794 -7654 497414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 532794 -7654 533414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 568794 -7654 569414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 29866 592650 30486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 65866 592650 66486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 101866 592650 102486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 137866 592650 138486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 173866 592650 174486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 209866 592650 210486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 245866 592650 246486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 281866 592650 282486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 317866 592650 318486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 353866 592650 354486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 389866 592650 390486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 425866 592650 426486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 461866 592650 462486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 497866 592650 498486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 533866 592650 534486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 569866 592650 570486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 605866 592650 606486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 641866 592650 642486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 677866 592650 678486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 24294 -7654 24914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 60294 -7654 60914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 60294 248684 60914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 96294 -7654 96914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 96294 248684 96914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 -7654 132914 73000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 137000 132914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 248684 132914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 -7654 168914 73000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 248684 168914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 204294 -7654 204914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 204294 248684 204914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 240294 -7654 240914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 240294 248684 240914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 276294 -7654 276914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 276294 248684 276914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 -7654 312914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 248684 312914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 348294 -7654 348914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 348294 248684 348914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 384294 -7654 384914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 384294 248684 384914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 420294 -7654 420914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 456294 -7654 456914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 492294 -7654 492914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 528294 -7654 528914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 564294 -7654 564914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 25366 592650 25986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 61366 592650 61986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 97366 592650 97986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 133366 592650 133986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 169366 592650 169986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 205366 592650 205986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 241366 592650 241986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 277366 592650 277986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 313366 592650 313986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 349366 592650 349986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 385366 592650 385986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 421366 592650 421986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 457366 592650 457986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 493366 592650 493986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 529366 592650 529986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 565366 592650 565986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 601366 592650 601986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 637366 592650 637986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 673366 592650 673986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 33294 -7654 33914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 69294 -7654 69914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 69294 248684 69914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 -7654 105914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 248684 105914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 -7654 141914 73000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 248684 141914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 -7654 177914 73000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 137000 177914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 248684 177914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 213294 -7654 213914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 213294 248684 213914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 -7654 249914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 248684 249914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 285294 -7654 285914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 285294 248684 285914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 321294 -7654 321914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 321294 248684 321914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 357294 -7654 357914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 357294 248684 357914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 393294 -7654 393914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 393294 248684 393914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 429294 -7654 429914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 465294 -7654 465914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 501294 -7654 501914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 537294 -7654 537914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 573294 -7654 573914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 34366 592650 34986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 70366 592650 70986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 106366 592650 106986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 142366 592650 142986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 178366 592650 178986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 214366 592650 214986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 250366 592650 250986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 286366 592650 286986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 322366 592650 322986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 358366 592650 358986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 394366 592650 394986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 430366 592650 430986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 466366 592650 466986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 502366 592650 502986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 538366 592650 538986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 574366 592650 574986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 610366 592650 610986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 646366 592650 646986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 682366 592650 682986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 6294 -7654 6914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 42294 -7654 42914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 -7654 78914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 248684 78914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 -7654 114914 73000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 137000 114914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 248684 114914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 -7654 150914 73000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 248684 150914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 -7654 186914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 248684 186914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 -7654 222914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 248684 222914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 -7654 258914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 248684 258914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 -7654 294914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 248684 294914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 -7654 330914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 248684 330914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 -7654 366914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 248684 366914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 402294 -7654 402914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 438294 -7654 438914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 474294 -7654 474914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 510294 -7654 510914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 546294 -7654 546914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 582294 -7654 582914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 7366 592650 7986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 43366 592650 43986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 79366 592650 79986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 115366 592650 115986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 151366 592650 151986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 187366 592650 187986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 223366 592650 223986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 259366 592650 259986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 295366 592650 295986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 331366 592650 331986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 367366 592650 367986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 403366 592650 403986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 439366 592650 439986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 475366 592650 475986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 511366 592650 511986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 547366 592650 547986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 583366 592650 583986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 619366 592650 619986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 655366 592650 655986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 691366 592650 691986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 15294 -7654 15914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 51294 -7654 51914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 51294 248684 51914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 -7654 87914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 248684 87914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 -7654 123914 73000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 137000 123914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 248684 123914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 -7654 159914 73000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 248684 159914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 -7654 195914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 248684 195914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 -7654 231914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 248684 231914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 -7654 267914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 248684 267914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 -7654 303914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 248684 303914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 -7654 339914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 248684 339914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 -7654 375914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 248684 375914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 411294 -7654 411914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 447294 -7654 447914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 483294 -7654 483914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 519294 -7654 519914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 555294 -7654 555914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 16366 592650 16986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 52366 592650 52986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 88366 592650 88986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 124366 592650 124986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 160366 592650 160986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 196366 592650 196986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 232366 592650 232986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 268366 592650 268986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 304366 592650 304986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 340366 592650 340986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 376366 592650 376986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 412366 592650 412986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 448366 592650 448986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 484366 592650 484986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 520366 592650 520986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 556366 592650 556986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 592366 592650 592986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 628366 592650 628986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 664366 592650 664986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 700366 592650 700986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
