VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1426.380 2924.800 1427.580 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3486.100 2.400 3487.300 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3224.980 2.400 3226.180 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2964.540 2.400 2965.740 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1692.260 2924.800 1693.460 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2703.420 2.400 2704.620 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2442.980 2.400 2444.180 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2182.540 2.400 2183.740 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1921.420 2.400 1922.620 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1660.980 2.400 1662.180 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1399.860 2.400 1401.060 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1139.420 2.400 1140.620 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 878.980 2.400 880.180 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 617.860 2.400 619.060 ;
    END
  END analog_io[28]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1958.140 2924.800 1959.340 ;
    END
  END analog_io[2]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2223.340 2924.800 2224.540 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2489.220 2924.800 2490.420 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2755.100 2924.800 2756.300 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3020.300 2924.800 3021.500 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3286.180 2924.800 3287.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 32.380 2924.800 33.580 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2289.980 2924.800 2291.180 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2555.860 2924.800 2557.060 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2821.060 2924.800 2822.260 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3086.940 2924.800 3088.140 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3352.820 2924.800 3354.020 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 230.940 2924.800 232.140 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3420.820 2.400 3422.020 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3159.700 2.400 3160.900 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2899.260 2.400 2900.460 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2638.820 2.400 2640.020 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2377.700 2.400 2378.900 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2117.260 2.400 2118.460 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 430.180 2924.800 431.380 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1856.140 2.400 1857.340 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1595.700 2.400 1596.900 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1335.260 2.400 1336.460 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1074.140 2.400 1075.340 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 813.700 2.400 814.900 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 552.580 2.400 553.780 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 357.420 2.400 358.620 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 161.580 2.400 162.780 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 629.420 2924.800 630.620 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 828.660 2924.800 829.860 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1027.900 2924.800 1029.100 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1227.140 2924.800 1228.340 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1493.020 2924.800 1494.220 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1758.900 2924.800 1760.100 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2024.100 2924.800 2025.300 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 164.980 2924.800 166.180 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2422.580 2924.800 2423.780 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2688.460 2924.800 2689.660 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2954.340 2924.800 2955.540 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3219.540 2924.800 3220.740 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3485.420 2924.800 3486.620 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 364.220 2924.800 365.420 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3290.260 2.400 3291.460 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3029.820 2.400 3031.020 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2768.700 2.400 2769.900 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2508.260 2.400 2509.460 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2247.140 2.400 2248.340 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1986.700 2.400 1987.900 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 563.460 2924.800 564.660 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1726.260 2.400 1727.460 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1465.140 2.400 1466.340 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1204.700 2.400 1205.900 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 943.580 2.400 944.780 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 683.140 2.400 684.340 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 422.700 2.400 423.900 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 226.860 2.400 228.060 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 31.700 2.400 32.900 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 762.700 2924.800 763.900 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 961.940 2924.800 963.140 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1161.180 2924.800 1162.380 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1360.420 2924.800 1361.620 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1625.620 2924.800 1626.820 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1891.500 2924.800 1892.700 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2157.380 2924.800 2158.580 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 98.340 2924.800 99.540 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2356.620 2924.800 2357.820 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2621.820 2924.800 2623.020 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2887.700 2924.800 2888.900 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3153.580 2924.800 3154.780 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3418.780 2924.800 3419.980 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 297.580 2924.800 298.780 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3355.540 2.400 3356.740 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3095.100 2.400 3096.300 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2833.980 2.400 2835.180 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2573.540 2.400 2574.740 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2312.420 2.400 2313.620 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2051.980 2.400 2053.180 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 496.820 2924.800 498.020 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1791.540 2.400 1792.740 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1530.420 2.400 1531.620 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1269.980 2.400 1271.180 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1008.860 2.400 1010.060 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 748.420 2.400 749.620 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 487.300 2.400 488.500 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 292.140 2.400 293.340 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 96.300 2.400 97.500 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 696.060 2924.800 697.260 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 895.300 2924.800 896.500 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1094.540 2924.800 1095.740 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1293.780 2924.800 1294.980 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1559.660 2924.800 1560.860 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1824.860 2924.800 1826.060 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2090.740 2924.800 2091.940 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.230 -4.800 629.790 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2402.530 -4.800 2403.090 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2420.010 -4.800 2420.570 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2437.950 -4.800 2438.510 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2455.430 -4.800 2455.990 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2473.370 -4.800 2473.930 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2490.850 -4.800 2491.410 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2508.790 -4.800 2509.350 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2526.730 -4.800 2527.290 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2544.210 -4.800 2544.770 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2562.150 -4.800 2562.710 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.330 -4.800 806.890 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2579.630 -4.800 2580.190 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2597.570 -4.800 2598.130 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2615.050 -4.800 2615.610 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2632.990 -4.800 2633.550 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2650.470 -4.800 2651.030 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2668.410 -4.800 2668.970 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2685.890 -4.800 2686.450 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2703.830 -4.800 2704.390 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2721.770 -4.800 2722.330 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2739.250 -4.800 2739.810 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.270 -4.800 824.830 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2757.190 -4.800 2757.750 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2774.670 -4.800 2775.230 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2792.610 -4.800 2793.170 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2810.090 -4.800 2810.650 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2828.030 -4.800 2828.590 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2845.510 -4.800 2846.070 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2863.450 -4.800 2864.010 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2881.390 -4.800 2881.950 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 841.750 -4.800 842.310 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.690 -4.800 860.250 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 877.170 -4.800 877.730 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.110 -4.800 895.670 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 912.590 -4.800 913.150 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 930.530 -4.800 931.090 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 948.470 -4.800 949.030 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.710 -4.800 647.270 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 983.890 -4.800 984.450 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.370 -4.800 1001.930 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1036.790 -4.800 1037.350 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1054.730 -4.800 1055.290 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1072.210 -4.800 1072.770 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1090.150 -4.800 1090.710 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1107.630 -4.800 1108.190 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1125.570 -4.800 1126.130 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1143.510 -4.800 1144.070 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.650 -4.800 665.210 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1160.990 -4.800 1161.550 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1178.930 -4.800 1179.490 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1196.410 -4.800 1196.970 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1214.350 -4.800 1214.910 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1231.830 -4.800 1232.390 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1249.770 -4.800 1250.330 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1267.250 -4.800 1267.810 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1285.190 -4.800 1285.750 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1303.130 -4.800 1303.690 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1320.610 -4.800 1321.170 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.130 -4.800 682.690 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1338.550 -4.800 1339.110 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1356.030 -4.800 1356.590 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1373.970 -4.800 1374.530 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1391.450 -4.800 1392.010 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1409.390 -4.800 1409.950 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1426.870 -4.800 1427.430 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1444.810 -4.800 1445.370 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1462.750 -4.800 1463.310 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1480.230 -4.800 1480.790 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1498.170 -4.800 1498.730 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.070 -4.800 700.630 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1515.650 -4.800 1516.210 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1533.590 -4.800 1534.150 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1551.070 -4.800 1551.630 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1569.010 -4.800 1569.570 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1586.490 -4.800 1587.050 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1604.430 -4.800 1604.990 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1621.910 -4.800 1622.470 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1639.850 -4.800 1640.410 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1657.790 -4.800 1658.350 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1675.270 -4.800 1675.830 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.550 -4.800 718.110 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1693.210 -4.800 1693.770 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1710.690 -4.800 1711.250 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1728.630 -4.800 1729.190 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1746.110 -4.800 1746.670 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1764.050 -4.800 1764.610 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1781.530 -4.800 1782.090 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1799.470 -4.800 1800.030 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1817.410 -4.800 1817.970 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1834.890 -4.800 1835.450 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1852.830 -4.800 1853.390 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.490 -4.800 736.050 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1870.310 -4.800 1870.870 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1888.250 -4.800 1888.810 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1923.670 -4.800 1924.230 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1976.570 -4.800 1977.130 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1994.510 -4.800 1995.070 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2029.930 -4.800 2030.490 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.970 -4.800 753.530 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2047.870 -4.800 2048.430 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2065.350 -4.800 2065.910 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2083.290 -4.800 2083.850 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2100.770 -4.800 2101.330 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2118.710 -4.800 2119.270 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2136.190 -4.800 2136.750 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2154.130 -4.800 2154.690 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2172.070 -4.800 2172.630 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2189.550 -4.800 2190.110 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2207.490 -4.800 2208.050 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.910 -4.800 771.470 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2224.970 -4.800 2225.530 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2242.910 -4.800 2243.470 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2260.390 -4.800 2260.950 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2278.330 -4.800 2278.890 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2295.810 -4.800 2296.370 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2313.750 -4.800 2314.310 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2331.230 -4.800 2331.790 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2349.170 -4.800 2349.730 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2367.110 -4.800 2367.670 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2384.590 -4.800 2385.150 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.850 -4.800 789.410 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.750 -4.800 635.310 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2408.510 -4.800 2409.070 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2425.990 -4.800 2426.550 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2443.930 -4.800 2444.490 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2461.410 -4.800 2461.970 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2479.350 -4.800 2479.910 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2496.830 -4.800 2497.390 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2514.770 -4.800 2515.330 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2532.250 -4.800 2532.810 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2550.190 -4.800 2550.750 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2567.670 -4.800 2568.230 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 812.310 -4.800 812.870 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2585.610 -4.800 2586.170 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2603.550 -4.800 2604.110 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2621.030 -4.800 2621.590 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2638.970 -4.800 2639.530 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2656.450 -4.800 2657.010 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2674.390 -4.800 2674.950 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2691.870 -4.800 2692.430 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2709.810 -4.800 2710.370 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2727.290 -4.800 2727.850 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2745.230 -4.800 2745.790 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.250 -4.800 830.810 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2763.170 -4.800 2763.730 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2780.650 -4.800 2781.210 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2798.590 -4.800 2799.150 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2816.070 -4.800 2816.630 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2834.010 -4.800 2834.570 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2851.490 -4.800 2852.050 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2869.430 -4.800 2869.990 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 847.730 -4.800 848.290 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 865.670 -4.800 866.230 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 883.150 -4.800 883.710 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 901.090 -4.800 901.650 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 918.570 -4.800 919.130 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 936.510 -4.800 937.070 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 953.990 -4.800 954.550 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 971.930 -4.800 972.490 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.690 -4.800 653.250 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 989.410 -4.800 989.970 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1042.770 -4.800 1043.330 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1060.710 -4.800 1061.270 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1078.190 -4.800 1078.750 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1096.130 -4.800 1096.690 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1113.610 -4.800 1114.170 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1131.550 -4.800 1132.110 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1149.030 -4.800 1149.590 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.630 -4.800 671.190 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1166.970 -4.800 1167.530 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1184.910 -4.800 1185.470 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1202.390 -4.800 1202.950 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1220.330 -4.800 1220.890 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1237.810 -4.800 1238.370 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1255.750 -4.800 1256.310 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1273.230 -4.800 1273.790 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1291.170 -4.800 1291.730 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1308.650 -4.800 1309.210 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1326.590 -4.800 1327.150 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.110 -4.800 688.670 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1344.070 -4.800 1344.630 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1362.010 -4.800 1362.570 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1379.950 -4.800 1380.510 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1397.430 -4.800 1397.990 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1415.370 -4.800 1415.930 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1432.850 -4.800 1433.410 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1450.790 -4.800 1451.350 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1468.270 -4.800 1468.830 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1486.210 -4.800 1486.770 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1503.690 -4.800 1504.250 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.050 -4.800 706.610 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1521.630 -4.800 1522.190 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1539.570 -4.800 1540.130 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1557.050 -4.800 1557.610 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1574.990 -4.800 1575.550 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1592.470 -4.800 1593.030 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1610.410 -4.800 1610.970 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1627.890 -4.800 1628.450 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1645.830 -4.800 1646.390 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1663.310 -4.800 1663.870 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1681.250 -4.800 1681.810 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 723.530 -4.800 724.090 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1699.190 -4.800 1699.750 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1716.670 -4.800 1717.230 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1734.610 -4.800 1735.170 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1752.090 -4.800 1752.650 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1770.030 -4.800 1770.590 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1787.510 -4.800 1788.070 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1805.450 -4.800 1806.010 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1822.930 -4.800 1823.490 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1840.870 -4.800 1841.430 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1858.350 -4.800 1858.910 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.470 -4.800 742.030 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1876.290 -4.800 1876.850 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1894.230 -4.800 1894.790 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1929.650 -4.800 1930.210 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1982.550 -4.800 1983.110 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2000.490 -4.800 2001.050 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2017.970 -4.800 2018.530 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2035.910 -4.800 2036.470 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 758.950 -4.800 759.510 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2053.850 -4.800 2054.410 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2071.330 -4.800 2071.890 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2089.270 -4.800 2089.830 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2106.750 -4.800 2107.310 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2124.690 -4.800 2125.250 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2142.170 -4.800 2142.730 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2160.110 -4.800 2160.670 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2177.590 -4.800 2178.150 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2195.530 -4.800 2196.090 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2213.010 -4.800 2213.570 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.890 -4.800 777.450 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2230.950 -4.800 2231.510 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2248.890 -4.800 2249.450 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2266.370 -4.800 2266.930 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2284.310 -4.800 2284.870 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2301.790 -4.800 2302.350 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2319.730 -4.800 2320.290 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2337.210 -4.800 2337.770 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2355.150 -4.800 2355.710 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2372.630 -4.800 2373.190 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2390.570 -4.800 2391.130 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.370 -4.800 794.930 2.400 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.730 -4.800 641.290 2.400 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2414.030 -4.800 2414.590 2.400 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2431.970 -4.800 2432.530 2.400 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2449.450 -4.800 2450.010 2.400 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2467.390 -4.800 2467.950 2.400 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2485.330 -4.800 2485.890 2.400 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2502.810 -4.800 2503.370 2.400 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2520.750 -4.800 2521.310 2.400 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2538.230 -4.800 2538.790 2.400 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2556.170 -4.800 2556.730 2.400 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2573.650 -4.800 2574.210 2.400 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 818.290 -4.800 818.850 2.400 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2591.590 -4.800 2592.150 2.400 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2609.070 -4.800 2609.630 2.400 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2627.010 -4.800 2627.570 2.400 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2644.950 -4.800 2645.510 2.400 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2662.430 -4.800 2662.990 2.400 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2680.370 -4.800 2680.930 2.400 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2697.850 -4.800 2698.410 2.400 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2715.790 -4.800 2716.350 2.400 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2733.270 -4.800 2733.830 2.400 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2751.210 -4.800 2751.770 2.400 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 835.770 -4.800 836.330 2.400 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2768.690 -4.800 2769.250 2.400 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2786.630 -4.800 2787.190 2.400 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2804.110 -4.800 2804.670 2.400 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2822.050 -4.800 2822.610 2.400 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2839.990 -4.800 2840.550 2.400 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2857.470 -4.800 2858.030 2.400 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2875.410 -4.800 2875.970 2.400 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.710 -4.800 854.270 2.400 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 871.190 -4.800 871.750 2.400 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 889.130 -4.800 889.690 2.400 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 907.070 -4.800 907.630 2.400 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.550 -4.800 925.110 2.400 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.490 -4.800 943.050 2.400 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.970 -4.800 960.530 2.400 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 977.910 -4.800 978.470 2.400 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.670 -4.800 659.230 2.400 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.390 -4.800 995.950 2.400 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1030.810 -4.800 1031.370 2.400 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1048.750 -4.800 1049.310 2.400 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1066.690 -4.800 1067.250 2.400 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1084.170 -4.800 1084.730 2.400 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1102.110 -4.800 1102.670 2.400 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1119.590 -4.800 1120.150 2.400 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1137.530 -4.800 1138.090 2.400 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1155.010 -4.800 1155.570 2.400 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.150 -4.800 676.710 2.400 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1172.950 -4.800 1173.510 2.400 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1190.430 -4.800 1190.990 2.400 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1208.370 -4.800 1208.930 2.400 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1225.850 -4.800 1226.410 2.400 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1243.790 -4.800 1244.350 2.400 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1261.730 -4.800 1262.290 2.400 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1279.210 -4.800 1279.770 2.400 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1297.150 -4.800 1297.710 2.400 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1314.630 -4.800 1315.190 2.400 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1332.570 -4.800 1333.130 2.400 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.090 -4.800 694.650 2.400 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1350.050 -4.800 1350.610 2.400 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1367.990 -4.800 1368.550 2.400 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1385.470 -4.800 1386.030 2.400 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1403.410 -4.800 1403.970 2.400 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1421.350 -4.800 1421.910 2.400 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1438.830 -4.800 1439.390 2.400 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1456.770 -4.800 1457.330 2.400 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1474.250 -4.800 1474.810 2.400 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1492.190 -4.800 1492.750 2.400 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1509.670 -4.800 1510.230 2.400 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.030 -4.800 712.590 2.400 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1527.610 -4.800 1528.170 2.400 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1545.090 -4.800 1545.650 2.400 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1563.030 -4.800 1563.590 2.400 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1580.970 -4.800 1581.530 2.400 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1598.450 -4.800 1599.010 2.400 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1616.390 -4.800 1616.950 2.400 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1633.870 -4.800 1634.430 2.400 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1651.810 -4.800 1652.370 2.400 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1669.290 -4.800 1669.850 2.400 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1687.230 -4.800 1687.790 2.400 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.510 -4.800 730.070 2.400 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1704.710 -4.800 1705.270 2.400 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1722.650 -4.800 1723.210 2.400 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1740.130 -4.800 1740.690 2.400 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1758.070 -4.800 1758.630 2.400 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1776.010 -4.800 1776.570 2.400 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1793.490 -4.800 1794.050 2.400 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1811.430 -4.800 1811.990 2.400 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1828.910 -4.800 1829.470 2.400 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1846.850 -4.800 1847.410 2.400 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1864.330 -4.800 1864.890 2.400 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.450 -4.800 748.010 2.400 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1882.270 -4.800 1882.830 2.400 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1935.630 -4.800 1936.190 2.400 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1988.530 -4.800 1989.090 2.400 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2023.950 -4.800 2024.510 2.400 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2041.890 -4.800 2042.450 2.400 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 764.930 -4.800 765.490 2.400 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2059.370 -4.800 2059.930 2.400 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2077.310 -4.800 2077.870 2.400 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2094.790 -4.800 2095.350 2.400 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2112.730 -4.800 2113.290 2.400 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2130.670 -4.800 2131.230 2.400 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2148.150 -4.800 2148.710 2.400 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2166.090 -4.800 2166.650 2.400 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2183.570 -4.800 2184.130 2.400 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2201.510 -4.800 2202.070 2.400 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2218.990 -4.800 2219.550 2.400 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.870 -4.800 783.430 2.400 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2236.930 -4.800 2237.490 2.400 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2254.410 -4.800 2254.970 2.400 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2272.350 -4.800 2272.910 2.400 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2290.290 -4.800 2290.850 2.400 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2307.770 -4.800 2308.330 2.400 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2325.710 -4.800 2326.270 2.400 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2343.190 -4.800 2343.750 2.400 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2361.130 -4.800 2361.690 2.400 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2378.610 -4.800 2379.170 2.400 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2396.550 -4.800 2397.110 2.400 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.350 -4.800 800.910 2.400 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
    END
  END user_clock2
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
    END
  END user_irq[2]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -10.030 -4.670 -6.930 3524.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -10.030 -4.670 2929.650 -1.570 ;
    END
    PORT
      LAYER met5 ;
        RECT -10.030 3521.250 2929.650 3524.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2926.550 -4.670 2929.650 3524.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 8.970 -38.270 12.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.970 -38.270 192.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.970 -38.270 372.070 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.970 1243.420 372.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 548.970 -38.270 552.070 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 548.970 1243.420 552.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 728.970 -38.270 732.070 365.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 728.970 1243.420 732.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 908.970 -38.270 912.070 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 908.970 1243.420 912.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.970 -38.270 1092.070 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.970 1243.420 1092.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1268.970 -38.270 1272.070 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 1268.970 1243.420 1272.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1448.970 -38.270 1452.070 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 1448.970 1243.420 1452.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1628.970 -38.270 1632.070 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 1628.970 1243.420 1632.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1808.970 -38.270 1812.070 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 1808.970 1243.420 1812.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1988.970 -38.270 1992.070 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 1988.970 1243.420 1992.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2168.970 -38.270 2172.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2348.970 -38.270 2352.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2528.970 -38.270 2532.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2708.970 -38.270 2712.070 1500.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2708.970 1604.000 2712.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2888.970 -38.270 2892.070 3557.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 14.330 2963.250 17.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 194.330 2963.250 197.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 374.330 2963.250 377.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 554.330 2963.250 557.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 734.330 2963.250 737.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 914.330 2963.250 917.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1094.330 2963.250 1097.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1274.330 2963.250 1277.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1454.330 2963.250 1457.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1634.330 2963.250 1637.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1814.330 2963.250 1817.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1994.330 2963.250 1997.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2174.330 2963.250 2177.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2354.330 2963.250 2357.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2534.330 2963.250 2537.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2714.330 2963.250 2717.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2894.330 2963.250 2897.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3074.330 2963.250 3077.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3254.330 2963.250 3257.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3434.330 2963.250 3437.430 ;
    END
  END vccd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -19.630 -14.270 -16.530 3533.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -19.630 -14.270 2939.250 -11.170 ;
    END
    PORT
      LAYER met5 ;
        RECT -19.630 3530.850 2939.250 3533.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2936.150 -14.270 2939.250 3533.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 53.970 -38.270 57.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 233.970 -38.270 237.070 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 233.970 1243.420 237.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 413.970 -38.270 417.070 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 413.970 1243.420 417.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 593.970 -38.270 597.070 365.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 593.970 685.000 597.070 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 593.970 1243.420 597.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 773.970 -38.270 777.070 365.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 773.970 1243.420 777.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 953.970 -38.270 957.070 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 953.970 1243.420 957.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1133.970 -38.270 1137.070 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 1133.970 1243.420 1137.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1313.970 -38.270 1317.070 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 1313.970 1243.420 1317.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1493.970 -38.270 1497.070 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 1493.970 1243.420 1497.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1673.970 -38.270 1677.070 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 1673.970 1243.420 1677.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1853.970 -38.270 1857.070 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 1853.970 1243.420 1857.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2033.970 -38.270 2037.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2213.970 -38.270 2217.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2393.970 -38.270 2397.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2573.970 -38.270 2577.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2753.970 -38.270 2757.070 1500.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2753.970 1604.000 2757.070 3557.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 59.330 2963.250 62.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 239.330 2963.250 242.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 419.330 2963.250 422.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 599.330 2963.250 602.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 779.330 2963.250 782.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 959.330 2963.250 962.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1139.330 2963.250 1142.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1319.330 2963.250 1322.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1499.330 2963.250 1502.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1679.330 2963.250 1682.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1859.330 2963.250 1862.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2039.330 2963.250 2042.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2219.330 2963.250 2222.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2399.330 2963.250 2402.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2579.330 2963.250 2582.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2759.330 2963.250 2762.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2939.330 2963.250 2942.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3119.330 2963.250 3122.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3299.330 2963.250 3302.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3479.330 2963.250 3482.430 ;
    END
  END vccd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -29.230 -23.870 -26.130 3543.550 ;
    END
    PORT
      LAYER met5 ;
        RECT -29.230 -23.870 2948.850 -20.770 ;
    END
    PORT
      LAYER met5 ;
        RECT -29.230 3540.450 2948.850 3543.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 2945.750 -23.870 2948.850 3543.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 98.970 -38.270 102.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 278.970 -38.270 282.070 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 278.970 1243.420 282.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.970 -38.270 462.070 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.970 1243.420 462.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.970 -38.270 642.070 365.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.970 685.000 642.070 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.970 1243.420 642.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 818.970 -38.270 822.070 365.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 818.970 1243.420 822.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 998.970 -38.270 1002.070 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 998.970 1243.420 1002.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1178.970 -38.270 1182.070 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 1178.970 1243.420 1182.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1358.970 -38.270 1362.070 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 1358.970 1243.420 1362.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1538.970 -38.270 1542.070 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 1538.970 1243.420 1542.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1718.970 -38.270 1722.070 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 1718.970 1243.420 1722.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1898.970 -38.270 1902.070 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 1898.970 1243.420 1902.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2078.970 -38.270 2082.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2258.970 -38.270 2262.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2438.970 -38.270 2442.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2618.970 -38.270 2622.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2798.970 -38.270 2802.070 1500.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2798.970 1604.000 2802.070 3557.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 104.330 2963.250 107.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 284.330 2963.250 287.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 464.330 2963.250 467.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 644.330 2963.250 647.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 824.330 2963.250 827.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1004.330 2963.250 1007.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1184.330 2963.250 1187.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1364.330 2963.250 1367.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1544.330 2963.250 1547.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1724.330 2963.250 1727.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1904.330 2963.250 1907.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2084.330 2963.250 2087.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2264.330 2963.250 2267.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2444.330 2963.250 2447.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2624.330 2963.250 2627.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2804.330 2963.250 2807.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2984.330 2963.250 2987.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3164.330 2963.250 3167.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3344.330 2963.250 3347.430 ;
    END
  END vdda1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -38.830 -33.470 -35.730 3553.150 ;
    END
    PORT
      LAYER met5 ;
        RECT -38.830 -33.470 2958.450 -30.370 ;
    END
    PORT
      LAYER met5 ;
        RECT -38.830 3550.050 2958.450 3553.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2955.350 -33.470 2958.450 3553.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 143.970 -38.270 147.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 323.970 -38.270 327.070 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 323.970 1243.420 327.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 503.970 -38.270 507.070 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 503.970 1243.420 507.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 683.970 -38.270 687.070 365.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 683.970 1243.420 687.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 863.970 -38.270 867.070 365.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 863.970 685.000 867.070 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 863.970 1243.420 867.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1043.970 -38.270 1047.070 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 1043.970 1243.420 1047.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1223.970 -38.270 1227.070 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 1223.970 1243.420 1227.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.970 -38.270 1407.070 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.970 1243.420 1407.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1583.970 -38.270 1587.070 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 1583.970 1243.420 1587.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1763.970 -38.270 1767.070 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 1763.970 1243.420 1767.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1943.970 -38.270 1947.070 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 1943.970 1243.420 1947.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2123.970 -38.270 2127.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2303.970 -38.270 2307.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2483.970 -38.270 2487.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2663.970 -38.270 2667.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2843.970 -38.270 2847.070 1500.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2843.970 1604.000 2847.070 3557.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 149.330 2963.250 152.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 329.330 2963.250 332.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 509.330 2963.250 512.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 689.330 2963.250 692.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 869.330 2963.250 872.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1049.330 2963.250 1052.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1229.330 2963.250 1232.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1409.330 2963.250 1412.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1589.330 2963.250 1592.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1769.330 2963.250 1772.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1949.330 2963.250 1952.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2129.330 2963.250 2132.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2309.330 2963.250 2312.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2489.330 2963.250 2492.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2669.330 2963.250 2672.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2849.330 2963.250 2852.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3029.330 2963.250 3032.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3209.330 2963.250 3212.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3389.330 2963.250 3392.430 ;
    END
  END vdda2
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -34.030 -28.670 -30.930 3548.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 -28.670 2953.650 -25.570 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3545.250 2953.650 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2950.550 -28.670 2953.650 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 121.470 -38.270 124.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 301.470 -38.270 304.570 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 301.470 1243.420 304.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.470 -38.270 484.570 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.470 1243.420 484.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 661.470 -38.270 664.570 365.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 661.470 685.000 664.570 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 661.470 1243.420 664.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 841.470 -38.270 844.570 365.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 841.470 1243.420 844.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1021.470 -38.270 1024.570 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 1021.470 1243.420 1024.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1201.470 -38.270 1204.570 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 1201.470 1243.420 1204.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1381.470 -38.270 1384.570 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 1381.470 1243.420 1384.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1561.470 -38.270 1564.570 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 1561.470 1243.420 1564.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1741.470 -38.270 1744.570 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 1741.470 1243.420 1744.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1921.470 -38.270 1924.570 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 1921.470 1243.420 1924.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2101.470 -38.270 2104.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2281.470 -38.270 2284.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2461.470 -38.270 2464.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2641.470 -38.270 2644.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2821.470 -38.270 2824.570 1500.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2821.470 1604.000 2824.570 3557.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 126.830 2963.250 129.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 306.830 2963.250 309.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 486.830 2963.250 489.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 666.830 2963.250 669.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 846.830 2963.250 849.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1026.830 2963.250 1029.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1206.830 2963.250 1209.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1386.830 2963.250 1389.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1566.830 2963.250 1569.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1746.830 2963.250 1749.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1926.830 2963.250 1929.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2106.830 2963.250 2109.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2286.830 2963.250 2289.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2466.830 2963.250 2469.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2646.830 2963.250 2649.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2826.830 2963.250 2829.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3006.830 2963.250 3009.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3186.830 2963.250 3189.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3366.830 2963.250 3369.930 ;
    END
  END vssa1
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -43.630 -38.270 -40.530 3557.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 -38.270 2963.250 -35.170 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3554.850 2963.250 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2960.150 -38.270 2963.250 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 166.470 -38.270 169.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 346.470 -38.270 349.570 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 346.470 1243.420 349.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 526.470 -38.270 529.570 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 526.470 1243.420 529.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 706.470 -38.270 709.570 365.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 706.470 1243.420 709.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 886.470 -38.270 889.570 365.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 886.470 685.000 889.570 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 886.470 1243.420 889.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1066.470 -38.270 1069.570 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 1066.470 1243.420 1069.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1246.470 -38.270 1249.570 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 1246.470 1243.420 1249.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1426.470 -38.270 1429.570 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 1426.470 1243.420 1429.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1606.470 -38.270 1609.570 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 1606.470 1243.420 1609.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1786.470 -38.270 1789.570 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 1786.470 1243.420 1789.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1966.470 -38.270 1969.570 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 1966.470 1243.420 1969.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2146.470 -38.270 2149.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2326.470 -38.270 2329.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2506.470 -38.270 2509.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2686.470 -38.270 2689.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2866.470 -38.270 2869.570 3557.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 171.830 2963.250 174.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 351.830 2963.250 354.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 531.830 2963.250 534.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 711.830 2963.250 714.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 891.830 2963.250 894.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1071.830 2963.250 1074.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1251.830 2963.250 1254.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1431.830 2963.250 1434.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1611.830 2963.250 1614.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1791.830 2963.250 1794.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1971.830 2963.250 1974.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2151.830 2963.250 2154.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2331.830 2963.250 2334.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2511.830 2963.250 2514.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2691.830 2963.250 2694.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2871.830 2963.250 2874.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3051.830 2963.250 3054.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3231.830 2963.250 3234.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3411.830 2963.250 3414.930 ;
    END
  END vssa2
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -14.830 -9.470 -11.730 3529.150 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 -9.470 2934.450 -6.370 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 3526.050 2934.450 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2931.350 -9.470 2934.450 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 31.470 -38.270 34.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 211.470 -38.270 214.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 391.470 -38.270 394.570 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 391.470 1243.420 394.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 571.470 -38.270 574.570 365.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 571.470 685.000 574.570 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 571.470 1243.420 574.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 751.470 -38.270 754.570 365.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 751.470 1243.420 754.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 931.470 -38.270 934.570 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 931.470 1243.420 934.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1111.470 -38.270 1114.570 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 1111.470 1243.420 1114.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1291.470 -38.270 1294.570 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 1291.470 1243.420 1294.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1471.470 -38.270 1474.570 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 1471.470 1243.420 1474.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1651.470 -38.270 1654.570 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 1651.470 1243.420 1654.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1831.470 -38.270 1834.570 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 1831.470 1243.420 1834.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2011.470 -38.270 2014.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2191.470 -38.270 2194.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2371.470 -38.270 2374.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2551.470 -38.270 2554.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2731.470 -38.270 2734.570 1500.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2731.470 1604.000 2734.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2911.470 -38.270 2914.570 3557.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 36.830 2963.250 39.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 216.830 2963.250 219.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 396.830 2963.250 399.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 576.830 2963.250 579.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 756.830 2963.250 759.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 936.830 2963.250 939.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1116.830 2963.250 1119.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1296.830 2963.250 1299.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1476.830 2963.250 1479.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1656.830 2963.250 1659.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1836.830 2963.250 1839.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2016.830 2963.250 2019.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2196.830 2963.250 2199.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2376.830 2963.250 2379.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2556.830 2963.250 2559.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2736.830 2963.250 2739.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2916.830 2963.250 2919.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3096.830 2963.250 3099.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3276.830 2963.250 3279.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3456.830 2963.250 3459.930 ;
    END
  END vssd1
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -24.430 -19.070 -21.330 3538.750 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 -19.070 2944.050 -15.970 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3535.650 2944.050 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2940.950 -19.070 2944.050 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 76.470 -38.270 79.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 256.470 -38.270 259.570 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 256.470 1243.420 259.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 436.470 -38.270 439.570 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 436.470 1243.420 439.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 616.470 -38.270 619.570 365.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 616.470 685.000 619.570 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 616.470 1243.420 619.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 796.470 -38.270 799.570 365.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 796.470 1243.420 799.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 976.470 -38.270 979.570 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 976.470 1243.420 979.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1156.470 -38.270 1159.570 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 1156.470 1243.420 1159.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1336.470 -38.270 1339.570 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 1336.470 1243.420 1339.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1516.470 -38.270 1519.570 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 1516.470 1243.420 1519.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1696.470 -38.270 1699.570 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 1696.470 1243.420 1699.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1876.470 -38.270 1879.570 1142.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 1876.470 1243.420 1879.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2056.470 -38.270 2059.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2236.470 -38.270 2239.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2416.470 -38.270 2419.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2596.470 -38.270 2599.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2776.470 -38.270 2779.570 1500.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2776.470 1604.000 2779.570 3557.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 81.830 2963.250 84.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 261.830 2963.250 264.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 441.830 2963.250 444.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 621.830 2963.250 624.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 801.830 2963.250 804.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 981.830 2963.250 984.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1161.830 2963.250 1164.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1341.830 2963.250 1344.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1521.830 2963.250 1524.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1701.830 2963.250 1704.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1881.830 2963.250 1884.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2061.830 2963.250 2064.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2241.830 2963.250 2244.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2421.830 2963.250 2424.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2601.830 2963.250 2604.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2781.830 2963.250 2784.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2961.830 2963.250 2964.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3141.830 2963.250 3144.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3321.830 2963.250 3324.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3501.830 2963.250 3504.930 ;
    END
  END vssd2
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.710 -4.800 3.270 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.230 -4.800 8.790 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.210 -4.800 14.770 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.130 -4.800 38.690 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.150 -4.800 239.710 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.630 -4.800 257.190 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.570 -4.800 275.130 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.050 -4.800 292.610 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.990 -4.800 310.550 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.470 -4.800 328.030 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.410 -4.800 345.970 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.890 -4.800 363.450 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.830 -4.800 381.390 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.310 -4.800 398.870 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.590 -4.800 62.150 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.250 -4.800 416.810 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.190 -4.800 434.750 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.670 -4.800 452.230 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.610 -4.800 470.170 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.090 -4.800 487.650 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.030 -4.800 505.590 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.510 -4.800 523.070 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.450 -4.800 541.010 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.930 -4.800 558.490 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.870 -4.800 576.430 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.050 -4.800 85.610 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.810 -4.800 594.370 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.290 -4.800 611.850 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.970 -4.800 109.530 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.430 -4.800 132.990 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.370 -4.800 150.930 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.850 -4.800 168.410 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.790 -4.800 186.350 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.270 -4.800 203.830 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.210 -4.800 221.770 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.190 -4.800 20.750 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.650 -4.800 44.210 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.670 -4.800 245.230 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.610 -4.800 263.170 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.090 -4.800 280.650 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.030 -4.800 298.590 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.970 -4.800 316.530 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.450 -4.800 334.010 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.390 -4.800 351.950 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.870 -4.800 369.430 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.810 -4.800 387.370 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.290 -4.800 404.850 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.570 -4.800 68.130 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.230 -4.800 422.790 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.710 -4.800 440.270 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.650 -4.800 458.210 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.590 -4.800 476.150 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.070 -4.800 493.630 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.010 -4.800 511.570 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.490 -4.800 529.050 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.430 -4.800 546.990 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.910 -4.800 564.470 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.850 -4.800 582.410 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.030 -4.800 91.590 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.330 -4.800 599.890 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.270 -4.800 617.830 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.950 -4.800 115.510 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.410 -4.800 138.970 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.350 -4.800 156.910 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.830 -4.800 174.390 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.770 -4.800 192.330 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.250 -4.800 209.810 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.190 -4.800 227.750 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.630 -4.800 50.190 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.650 -4.800 251.210 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.590 -4.800 269.150 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.070 -4.800 286.630 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.010 -4.800 304.570 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.490 -4.800 322.050 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.430 -4.800 339.990 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.370 -4.800 357.930 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.850 -4.800 375.410 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.790 -4.800 393.350 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.270 -4.800 410.830 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.550 -4.800 74.110 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.210 -4.800 428.770 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.690 -4.800 446.250 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.630 -4.800 464.190 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.110 -4.800 481.670 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.050 -4.800 499.610 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.530 -4.800 517.090 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.470 -4.800 535.030 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.410 -4.800 552.970 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.890 -4.800 570.450 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.830 -4.800 588.390 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.010 -4.800 97.570 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.310 -4.800 605.870 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.250 -4.800 623.810 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.930 -4.800 121.490 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.390 -4.800 144.950 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.870 -4.800 162.430 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.810 -4.800 180.370 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.750 -4.800 198.310 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.230 -4.800 215.790 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.170 -4.800 233.730 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.610 -4.800 56.170 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.530 -4.800 80.090 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.990 -4.800 103.550 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.450 -4.800 127.010 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.170 -4.800 26.730 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.150 -4.800 32.710 2.400 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 230.500 385.795 2826.000 1570.500 ;
      LAYER met1 ;
        RECT 13.870 6.160 2905.290 3515.220 ;
      LAYER met2 ;
        RECT 2.850 3517.320 40.150 3518.050 ;
        RECT 41.270 3517.320 121.110 3518.050 ;
        RECT 122.230 3517.320 202.070 3518.050 ;
        RECT 203.190 3517.320 283.490 3518.050 ;
        RECT 284.610 3517.320 364.450 3518.050 ;
        RECT 365.570 3517.320 445.410 3518.050 ;
        RECT 446.530 3517.320 526.830 3518.050 ;
        RECT 527.950 3517.320 607.790 3518.050 ;
        RECT 608.910 3517.320 688.750 3518.050 ;
        RECT 689.870 3517.320 770.170 3518.050 ;
        RECT 771.290 3517.320 851.130 3518.050 ;
        RECT 852.250 3517.320 932.090 3518.050 ;
        RECT 933.210 3517.320 1013.510 3518.050 ;
        RECT 1014.630 3517.320 1094.470 3518.050 ;
        RECT 1095.590 3517.320 1175.430 3518.050 ;
        RECT 1176.550 3517.320 1256.850 3518.050 ;
        RECT 1257.970 3517.320 1337.810 3518.050 ;
        RECT 1338.930 3517.320 1418.770 3518.050 ;
        RECT 1419.890 3517.320 1500.190 3518.050 ;
        RECT 1501.310 3517.320 1581.150 3518.050 ;
        RECT 1582.270 3517.320 1662.110 3518.050 ;
        RECT 1663.230 3517.320 1743.530 3518.050 ;
        RECT 1744.650 3517.320 1824.490 3518.050 ;
        RECT 1825.610 3517.320 1905.450 3518.050 ;
        RECT 1906.570 3517.320 1986.870 3518.050 ;
        RECT 1987.990 3517.320 2067.830 3518.050 ;
        RECT 2068.950 3517.320 2148.790 3518.050 ;
        RECT 2149.910 3517.320 2230.210 3518.050 ;
        RECT 2231.330 3517.320 2311.170 3518.050 ;
        RECT 2312.290 3517.320 2392.130 3518.050 ;
        RECT 2393.250 3517.320 2473.550 3518.050 ;
        RECT 2474.670 3517.320 2554.510 3518.050 ;
        RECT 2555.630 3517.320 2635.470 3518.050 ;
        RECT 2636.590 3517.320 2716.890 3518.050 ;
        RECT 2718.010 3517.320 2797.850 3518.050 ;
        RECT 2798.970 3517.320 2878.810 3518.050 ;
        RECT 2879.930 3517.320 2917.230 3518.050 ;
        RECT 2.850 2.680 2917.230 3517.320 ;
        RECT 3.550 1.630 7.950 2.680 ;
        RECT 9.070 1.630 13.930 2.680 ;
        RECT 15.050 1.630 19.910 2.680 ;
        RECT 21.030 1.630 25.890 2.680 ;
        RECT 27.010 1.630 31.870 2.680 ;
        RECT 32.990 1.630 37.850 2.680 ;
        RECT 38.970 1.630 43.370 2.680 ;
        RECT 44.490 1.630 49.350 2.680 ;
        RECT 50.470 1.630 55.330 2.680 ;
        RECT 56.450 1.630 61.310 2.680 ;
        RECT 62.430 1.630 67.290 2.680 ;
        RECT 68.410 1.630 73.270 2.680 ;
        RECT 74.390 1.630 79.250 2.680 ;
        RECT 80.370 1.630 84.770 2.680 ;
        RECT 85.890 1.630 90.750 2.680 ;
        RECT 91.870 1.630 96.730 2.680 ;
        RECT 97.850 1.630 102.710 2.680 ;
        RECT 103.830 1.630 108.690 2.680 ;
        RECT 109.810 1.630 114.670 2.680 ;
        RECT 115.790 1.630 120.650 2.680 ;
        RECT 121.770 1.630 126.170 2.680 ;
        RECT 127.290 1.630 132.150 2.680 ;
        RECT 133.270 1.630 138.130 2.680 ;
        RECT 139.250 1.630 144.110 2.680 ;
        RECT 145.230 1.630 150.090 2.680 ;
        RECT 151.210 1.630 156.070 2.680 ;
        RECT 157.190 1.630 161.590 2.680 ;
        RECT 162.710 1.630 167.570 2.680 ;
        RECT 168.690 1.630 173.550 2.680 ;
        RECT 174.670 1.630 179.530 2.680 ;
        RECT 180.650 1.630 185.510 2.680 ;
        RECT 186.630 1.630 191.490 2.680 ;
        RECT 192.610 1.630 197.470 2.680 ;
        RECT 198.590 1.630 202.990 2.680 ;
        RECT 204.110 1.630 208.970 2.680 ;
        RECT 210.090 1.630 214.950 2.680 ;
        RECT 216.070 1.630 220.930 2.680 ;
        RECT 222.050 1.630 226.910 2.680 ;
        RECT 228.030 1.630 232.890 2.680 ;
        RECT 234.010 1.630 238.870 2.680 ;
        RECT 239.990 1.630 244.390 2.680 ;
        RECT 245.510 1.630 250.370 2.680 ;
        RECT 251.490 1.630 256.350 2.680 ;
        RECT 257.470 1.630 262.330 2.680 ;
        RECT 263.450 1.630 268.310 2.680 ;
        RECT 269.430 1.630 274.290 2.680 ;
        RECT 275.410 1.630 279.810 2.680 ;
        RECT 280.930 1.630 285.790 2.680 ;
        RECT 286.910 1.630 291.770 2.680 ;
        RECT 292.890 1.630 297.750 2.680 ;
        RECT 298.870 1.630 303.730 2.680 ;
        RECT 304.850 1.630 309.710 2.680 ;
        RECT 310.830 1.630 315.690 2.680 ;
        RECT 316.810 1.630 321.210 2.680 ;
        RECT 322.330 1.630 327.190 2.680 ;
        RECT 328.310 1.630 333.170 2.680 ;
        RECT 334.290 1.630 339.150 2.680 ;
        RECT 340.270 1.630 345.130 2.680 ;
        RECT 346.250 1.630 351.110 2.680 ;
        RECT 352.230 1.630 357.090 2.680 ;
        RECT 358.210 1.630 362.610 2.680 ;
        RECT 363.730 1.630 368.590 2.680 ;
        RECT 369.710 1.630 374.570 2.680 ;
        RECT 375.690 1.630 380.550 2.680 ;
        RECT 381.670 1.630 386.530 2.680 ;
        RECT 387.650 1.630 392.510 2.680 ;
        RECT 393.630 1.630 398.030 2.680 ;
        RECT 399.150 1.630 404.010 2.680 ;
        RECT 405.130 1.630 409.990 2.680 ;
        RECT 411.110 1.630 415.970 2.680 ;
        RECT 417.090 1.630 421.950 2.680 ;
        RECT 423.070 1.630 427.930 2.680 ;
        RECT 429.050 1.630 433.910 2.680 ;
        RECT 435.030 1.630 439.430 2.680 ;
        RECT 440.550 1.630 445.410 2.680 ;
        RECT 446.530 1.630 451.390 2.680 ;
        RECT 452.510 1.630 457.370 2.680 ;
        RECT 458.490 1.630 463.350 2.680 ;
        RECT 464.470 1.630 469.330 2.680 ;
        RECT 470.450 1.630 475.310 2.680 ;
        RECT 476.430 1.630 480.830 2.680 ;
        RECT 481.950 1.630 486.810 2.680 ;
        RECT 487.930 1.630 492.790 2.680 ;
        RECT 493.910 1.630 498.770 2.680 ;
        RECT 499.890 1.630 504.750 2.680 ;
        RECT 505.870 1.630 510.730 2.680 ;
        RECT 511.850 1.630 516.250 2.680 ;
        RECT 517.370 1.630 522.230 2.680 ;
        RECT 523.350 1.630 528.210 2.680 ;
        RECT 529.330 1.630 534.190 2.680 ;
        RECT 535.310 1.630 540.170 2.680 ;
        RECT 541.290 1.630 546.150 2.680 ;
        RECT 547.270 1.630 552.130 2.680 ;
        RECT 553.250 1.630 557.650 2.680 ;
        RECT 558.770 1.630 563.630 2.680 ;
        RECT 564.750 1.630 569.610 2.680 ;
        RECT 570.730 1.630 575.590 2.680 ;
        RECT 576.710 1.630 581.570 2.680 ;
        RECT 582.690 1.630 587.550 2.680 ;
        RECT 588.670 1.630 593.530 2.680 ;
        RECT 594.650 1.630 599.050 2.680 ;
        RECT 600.170 1.630 605.030 2.680 ;
        RECT 606.150 1.630 611.010 2.680 ;
        RECT 612.130 1.630 616.990 2.680 ;
        RECT 618.110 1.630 622.970 2.680 ;
        RECT 624.090 1.630 628.950 2.680 ;
        RECT 630.070 1.630 634.470 2.680 ;
        RECT 635.590 1.630 640.450 2.680 ;
        RECT 641.570 1.630 646.430 2.680 ;
        RECT 647.550 1.630 652.410 2.680 ;
        RECT 653.530 1.630 658.390 2.680 ;
        RECT 659.510 1.630 664.370 2.680 ;
        RECT 665.490 1.630 670.350 2.680 ;
        RECT 671.470 1.630 675.870 2.680 ;
        RECT 676.990 1.630 681.850 2.680 ;
        RECT 682.970 1.630 687.830 2.680 ;
        RECT 688.950 1.630 693.810 2.680 ;
        RECT 694.930 1.630 699.790 2.680 ;
        RECT 700.910 1.630 705.770 2.680 ;
        RECT 706.890 1.630 711.750 2.680 ;
        RECT 712.870 1.630 717.270 2.680 ;
        RECT 718.390 1.630 723.250 2.680 ;
        RECT 724.370 1.630 729.230 2.680 ;
        RECT 730.350 1.630 735.210 2.680 ;
        RECT 736.330 1.630 741.190 2.680 ;
        RECT 742.310 1.630 747.170 2.680 ;
        RECT 748.290 1.630 752.690 2.680 ;
        RECT 753.810 1.630 758.670 2.680 ;
        RECT 759.790 1.630 764.650 2.680 ;
        RECT 765.770 1.630 770.630 2.680 ;
        RECT 771.750 1.630 776.610 2.680 ;
        RECT 777.730 1.630 782.590 2.680 ;
        RECT 783.710 1.630 788.570 2.680 ;
        RECT 789.690 1.630 794.090 2.680 ;
        RECT 795.210 1.630 800.070 2.680 ;
        RECT 801.190 1.630 806.050 2.680 ;
        RECT 807.170 1.630 812.030 2.680 ;
        RECT 813.150 1.630 818.010 2.680 ;
        RECT 819.130 1.630 823.990 2.680 ;
        RECT 825.110 1.630 829.970 2.680 ;
        RECT 831.090 1.630 835.490 2.680 ;
        RECT 836.610 1.630 841.470 2.680 ;
        RECT 842.590 1.630 847.450 2.680 ;
        RECT 848.570 1.630 853.430 2.680 ;
        RECT 854.550 1.630 859.410 2.680 ;
        RECT 860.530 1.630 865.390 2.680 ;
        RECT 866.510 1.630 870.910 2.680 ;
        RECT 872.030 1.630 876.890 2.680 ;
        RECT 878.010 1.630 882.870 2.680 ;
        RECT 883.990 1.630 888.850 2.680 ;
        RECT 889.970 1.630 894.830 2.680 ;
        RECT 895.950 1.630 900.810 2.680 ;
        RECT 901.930 1.630 906.790 2.680 ;
        RECT 907.910 1.630 912.310 2.680 ;
        RECT 913.430 1.630 918.290 2.680 ;
        RECT 919.410 1.630 924.270 2.680 ;
        RECT 925.390 1.630 930.250 2.680 ;
        RECT 931.370 1.630 936.230 2.680 ;
        RECT 937.350 1.630 942.210 2.680 ;
        RECT 943.330 1.630 948.190 2.680 ;
        RECT 949.310 1.630 953.710 2.680 ;
        RECT 954.830 1.630 959.690 2.680 ;
        RECT 960.810 1.630 965.670 2.680 ;
        RECT 966.790 1.630 971.650 2.680 ;
        RECT 972.770 1.630 977.630 2.680 ;
        RECT 978.750 1.630 983.610 2.680 ;
        RECT 984.730 1.630 989.130 2.680 ;
        RECT 990.250 1.630 995.110 2.680 ;
        RECT 996.230 1.630 1001.090 2.680 ;
        RECT 1002.210 1.630 1007.070 2.680 ;
        RECT 1008.190 1.630 1013.050 2.680 ;
        RECT 1014.170 1.630 1019.030 2.680 ;
        RECT 1020.150 1.630 1025.010 2.680 ;
        RECT 1026.130 1.630 1030.530 2.680 ;
        RECT 1031.650 1.630 1036.510 2.680 ;
        RECT 1037.630 1.630 1042.490 2.680 ;
        RECT 1043.610 1.630 1048.470 2.680 ;
        RECT 1049.590 1.630 1054.450 2.680 ;
        RECT 1055.570 1.630 1060.430 2.680 ;
        RECT 1061.550 1.630 1066.410 2.680 ;
        RECT 1067.530 1.630 1071.930 2.680 ;
        RECT 1073.050 1.630 1077.910 2.680 ;
        RECT 1079.030 1.630 1083.890 2.680 ;
        RECT 1085.010 1.630 1089.870 2.680 ;
        RECT 1090.990 1.630 1095.850 2.680 ;
        RECT 1096.970 1.630 1101.830 2.680 ;
        RECT 1102.950 1.630 1107.350 2.680 ;
        RECT 1108.470 1.630 1113.330 2.680 ;
        RECT 1114.450 1.630 1119.310 2.680 ;
        RECT 1120.430 1.630 1125.290 2.680 ;
        RECT 1126.410 1.630 1131.270 2.680 ;
        RECT 1132.390 1.630 1137.250 2.680 ;
        RECT 1138.370 1.630 1143.230 2.680 ;
        RECT 1144.350 1.630 1148.750 2.680 ;
        RECT 1149.870 1.630 1154.730 2.680 ;
        RECT 1155.850 1.630 1160.710 2.680 ;
        RECT 1161.830 1.630 1166.690 2.680 ;
        RECT 1167.810 1.630 1172.670 2.680 ;
        RECT 1173.790 1.630 1178.650 2.680 ;
        RECT 1179.770 1.630 1184.630 2.680 ;
        RECT 1185.750 1.630 1190.150 2.680 ;
        RECT 1191.270 1.630 1196.130 2.680 ;
        RECT 1197.250 1.630 1202.110 2.680 ;
        RECT 1203.230 1.630 1208.090 2.680 ;
        RECT 1209.210 1.630 1214.070 2.680 ;
        RECT 1215.190 1.630 1220.050 2.680 ;
        RECT 1221.170 1.630 1225.570 2.680 ;
        RECT 1226.690 1.630 1231.550 2.680 ;
        RECT 1232.670 1.630 1237.530 2.680 ;
        RECT 1238.650 1.630 1243.510 2.680 ;
        RECT 1244.630 1.630 1249.490 2.680 ;
        RECT 1250.610 1.630 1255.470 2.680 ;
        RECT 1256.590 1.630 1261.450 2.680 ;
        RECT 1262.570 1.630 1266.970 2.680 ;
        RECT 1268.090 1.630 1272.950 2.680 ;
        RECT 1274.070 1.630 1278.930 2.680 ;
        RECT 1280.050 1.630 1284.910 2.680 ;
        RECT 1286.030 1.630 1290.890 2.680 ;
        RECT 1292.010 1.630 1296.870 2.680 ;
        RECT 1297.990 1.630 1302.850 2.680 ;
        RECT 1303.970 1.630 1308.370 2.680 ;
        RECT 1309.490 1.630 1314.350 2.680 ;
        RECT 1315.470 1.630 1320.330 2.680 ;
        RECT 1321.450 1.630 1326.310 2.680 ;
        RECT 1327.430 1.630 1332.290 2.680 ;
        RECT 1333.410 1.630 1338.270 2.680 ;
        RECT 1339.390 1.630 1343.790 2.680 ;
        RECT 1344.910 1.630 1349.770 2.680 ;
        RECT 1350.890 1.630 1355.750 2.680 ;
        RECT 1356.870 1.630 1361.730 2.680 ;
        RECT 1362.850 1.630 1367.710 2.680 ;
        RECT 1368.830 1.630 1373.690 2.680 ;
        RECT 1374.810 1.630 1379.670 2.680 ;
        RECT 1380.790 1.630 1385.190 2.680 ;
        RECT 1386.310 1.630 1391.170 2.680 ;
        RECT 1392.290 1.630 1397.150 2.680 ;
        RECT 1398.270 1.630 1403.130 2.680 ;
        RECT 1404.250 1.630 1409.110 2.680 ;
        RECT 1410.230 1.630 1415.090 2.680 ;
        RECT 1416.210 1.630 1421.070 2.680 ;
        RECT 1422.190 1.630 1426.590 2.680 ;
        RECT 1427.710 1.630 1432.570 2.680 ;
        RECT 1433.690 1.630 1438.550 2.680 ;
        RECT 1439.670 1.630 1444.530 2.680 ;
        RECT 1445.650 1.630 1450.510 2.680 ;
        RECT 1451.630 1.630 1456.490 2.680 ;
        RECT 1457.610 1.630 1462.470 2.680 ;
        RECT 1463.590 1.630 1467.990 2.680 ;
        RECT 1469.110 1.630 1473.970 2.680 ;
        RECT 1475.090 1.630 1479.950 2.680 ;
        RECT 1481.070 1.630 1485.930 2.680 ;
        RECT 1487.050 1.630 1491.910 2.680 ;
        RECT 1493.030 1.630 1497.890 2.680 ;
        RECT 1499.010 1.630 1503.410 2.680 ;
        RECT 1504.530 1.630 1509.390 2.680 ;
        RECT 1510.510 1.630 1515.370 2.680 ;
        RECT 1516.490 1.630 1521.350 2.680 ;
        RECT 1522.470 1.630 1527.330 2.680 ;
        RECT 1528.450 1.630 1533.310 2.680 ;
        RECT 1534.430 1.630 1539.290 2.680 ;
        RECT 1540.410 1.630 1544.810 2.680 ;
        RECT 1545.930 1.630 1550.790 2.680 ;
        RECT 1551.910 1.630 1556.770 2.680 ;
        RECT 1557.890 1.630 1562.750 2.680 ;
        RECT 1563.870 1.630 1568.730 2.680 ;
        RECT 1569.850 1.630 1574.710 2.680 ;
        RECT 1575.830 1.630 1580.690 2.680 ;
        RECT 1581.810 1.630 1586.210 2.680 ;
        RECT 1587.330 1.630 1592.190 2.680 ;
        RECT 1593.310 1.630 1598.170 2.680 ;
        RECT 1599.290 1.630 1604.150 2.680 ;
        RECT 1605.270 1.630 1610.130 2.680 ;
        RECT 1611.250 1.630 1616.110 2.680 ;
        RECT 1617.230 1.630 1621.630 2.680 ;
        RECT 1622.750 1.630 1627.610 2.680 ;
        RECT 1628.730 1.630 1633.590 2.680 ;
        RECT 1634.710 1.630 1639.570 2.680 ;
        RECT 1640.690 1.630 1645.550 2.680 ;
        RECT 1646.670 1.630 1651.530 2.680 ;
        RECT 1652.650 1.630 1657.510 2.680 ;
        RECT 1658.630 1.630 1663.030 2.680 ;
        RECT 1664.150 1.630 1669.010 2.680 ;
        RECT 1670.130 1.630 1674.990 2.680 ;
        RECT 1676.110 1.630 1680.970 2.680 ;
        RECT 1682.090 1.630 1686.950 2.680 ;
        RECT 1688.070 1.630 1692.930 2.680 ;
        RECT 1694.050 1.630 1698.910 2.680 ;
        RECT 1700.030 1.630 1704.430 2.680 ;
        RECT 1705.550 1.630 1710.410 2.680 ;
        RECT 1711.530 1.630 1716.390 2.680 ;
        RECT 1717.510 1.630 1722.370 2.680 ;
        RECT 1723.490 1.630 1728.350 2.680 ;
        RECT 1729.470 1.630 1734.330 2.680 ;
        RECT 1735.450 1.630 1739.850 2.680 ;
        RECT 1740.970 1.630 1745.830 2.680 ;
        RECT 1746.950 1.630 1751.810 2.680 ;
        RECT 1752.930 1.630 1757.790 2.680 ;
        RECT 1758.910 1.630 1763.770 2.680 ;
        RECT 1764.890 1.630 1769.750 2.680 ;
        RECT 1770.870 1.630 1775.730 2.680 ;
        RECT 1776.850 1.630 1781.250 2.680 ;
        RECT 1782.370 1.630 1787.230 2.680 ;
        RECT 1788.350 1.630 1793.210 2.680 ;
        RECT 1794.330 1.630 1799.190 2.680 ;
        RECT 1800.310 1.630 1805.170 2.680 ;
        RECT 1806.290 1.630 1811.150 2.680 ;
        RECT 1812.270 1.630 1817.130 2.680 ;
        RECT 1818.250 1.630 1822.650 2.680 ;
        RECT 1823.770 1.630 1828.630 2.680 ;
        RECT 1829.750 1.630 1834.610 2.680 ;
        RECT 1835.730 1.630 1840.590 2.680 ;
        RECT 1841.710 1.630 1846.570 2.680 ;
        RECT 1847.690 1.630 1852.550 2.680 ;
        RECT 1853.670 1.630 1858.070 2.680 ;
        RECT 1859.190 1.630 1864.050 2.680 ;
        RECT 1865.170 1.630 1870.030 2.680 ;
        RECT 1871.150 1.630 1876.010 2.680 ;
        RECT 1877.130 1.630 1881.990 2.680 ;
        RECT 1883.110 1.630 1887.970 2.680 ;
        RECT 1889.090 1.630 1893.950 2.680 ;
        RECT 1895.070 1.630 1899.470 2.680 ;
        RECT 1900.590 1.630 1905.450 2.680 ;
        RECT 1906.570 1.630 1911.430 2.680 ;
        RECT 1912.550 1.630 1917.410 2.680 ;
        RECT 1918.530 1.630 1923.390 2.680 ;
        RECT 1924.510 1.630 1929.370 2.680 ;
        RECT 1930.490 1.630 1935.350 2.680 ;
        RECT 1936.470 1.630 1940.870 2.680 ;
        RECT 1941.990 1.630 1946.850 2.680 ;
        RECT 1947.970 1.630 1952.830 2.680 ;
        RECT 1953.950 1.630 1958.810 2.680 ;
        RECT 1959.930 1.630 1964.790 2.680 ;
        RECT 1965.910 1.630 1970.770 2.680 ;
        RECT 1971.890 1.630 1976.290 2.680 ;
        RECT 1977.410 1.630 1982.270 2.680 ;
        RECT 1983.390 1.630 1988.250 2.680 ;
        RECT 1989.370 1.630 1994.230 2.680 ;
        RECT 1995.350 1.630 2000.210 2.680 ;
        RECT 2001.330 1.630 2006.190 2.680 ;
        RECT 2007.310 1.630 2012.170 2.680 ;
        RECT 2013.290 1.630 2017.690 2.680 ;
        RECT 2018.810 1.630 2023.670 2.680 ;
        RECT 2024.790 1.630 2029.650 2.680 ;
        RECT 2030.770 1.630 2035.630 2.680 ;
        RECT 2036.750 1.630 2041.610 2.680 ;
        RECT 2042.730 1.630 2047.590 2.680 ;
        RECT 2048.710 1.630 2053.570 2.680 ;
        RECT 2054.690 1.630 2059.090 2.680 ;
        RECT 2060.210 1.630 2065.070 2.680 ;
        RECT 2066.190 1.630 2071.050 2.680 ;
        RECT 2072.170 1.630 2077.030 2.680 ;
        RECT 2078.150 1.630 2083.010 2.680 ;
        RECT 2084.130 1.630 2088.990 2.680 ;
        RECT 2090.110 1.630 2094.510 2.680 ;
        RECT 2095.630 1.630 2100.490 2.680 ;
        RECT 2101.610 1.630 2106.470 2.680 ;
        RECT 2107.590 1.630 2112.450 2.680 ;
        RECT 2113.570 1.630 2118.430 2.680 ;
        RECT 2119.550 1.630 2124.410 2.680 ;
        RECT 2125.530 1.630 2130.390 2.680 ;
        RECT 2131.510 1.630 2135.910 2.680 ;
        RECT 2137.030 1.630 2141.890 2.680 ;
        RECT 2143.010 1.630 2147.870 2.680 ;
        RECT 2148.990 1.630 2153.850 2.680 ;
        RECT 2154.970 1.630 2159.830 2.680 ;
        RECT 2160.950 1.630 2165.810 2.680 ;
        RECT 2166.930 1.630 2171.790 2.680 ;
        RECT 2172.910 1.630 2177.310 2.680 ;
        RECT 2178.430 1.630 2183.290 2.680 ;
        RECT 2184.410 1.630 2189.270 2.680 ;
        RECT 2190.390 1.630 2195.250 2.680 ;
        RECT 2196.370 1.630 2201.230 2.680 ;
        RECT 2202.350 1.630 2207.210 2.680 ;
        RECT 2208.330 1.630 2212.730 2.680 ;
        RECT 2213.850 1.630 2218.710 2.680 ;
        RECT 2219.830 1.630 2224.690 2.680 ;
        RECT 2225.810 1.630 2230.670 2.680 ;
        RECT 2231.790 1.630 2236.650 2.680 ;
        RECT 2237.770 1.630 2242.630 2.680 ;
        RECT 2243.750 1.630 2248.610 2.680 ;
        RECT 2249.730 1.630 2254.130 2.680 ;
        RECT 2255.250 1.630 2260.110 2.680 ;
        RECT 2261.230 1.630 2266.090 2.680 ;
        RECT 2267.210 1.630 2272.070 2.680 ;
        RECT 2273.190 1.630 2278.050 2.680 ;
        RECT 2279.170 1.630 2284.030 2.680 ;
        RECT 2285.150 1.630 2290.010 2.680 ;
        RECT 2291.130 1.630 2295.530 2.680 ;
        RECT 2296.650 1.630 2301.510 2.680 ;
        RECT 2302.630 1.630 2307.490 2.680 ;
        RECT 2308.610 1.630 2313.470 2.680 ;
        RECT 2314.590 1.630 2319.450 2.680 ;
        RECT 2320.570 1.630 2325.430 2.680 ;
        RECT 2326.550 1.630 2330.950 2.680 ;
        RECT 2332.070 1.630 2336.930 2.680 ;
        RECT 2338.050 1.630 2342.910 2.680 ;
        RECT 2344.030 1.630 2348.890 2.680 ;
        RECT 2350.010 1.630 2354.870 2.680 ;
        RECT 2355.990 1.630 2360.850 2.680 ;
        RECT 2361.970 1.630 2366.830 2.680 ;
        RECT 2367.950 1.630 2372.350 2.680 ;
        RECT 2373.470 1.630 2378.330 2.680 ;
        RECT 2379.450 1.630 2384.310 2.680 ;
        RECT 2385.430 1.630 2390.290 2.680 ;
        RECT 2391.410 1.630 2396.270 2.680 ;
        RECT 2397.390 1.630 2402.250 2.680 ;
        RECT 2403.370 1.630 2408.230 2.680 ;
        RECT 2409.350 1.630 2413.750 2.680 ;
        RECT 2414.870 1.630 2419.730 2.680 ;
        RECT 2420.850 1.630 2425.710 2.680 ;
        RECT 2426.830 1.630 2431.690 2.680 ;
        RECT 2432.810 1.630 2437.670 2.680 ;
        RECT 2438.790 1.630 2443.650 2.680 ;
        RECT 2444.770 1.630 2449.170 2.680 ;
        RECT 2450.290 1.630 2455.150 2.680 ;
        RECT 2456.270 1.630 2461.130 2.680 ;
        RECT 2462.250 1.630 2467.110 2.680 ;
        RECT 2468.230 1.630 2473.090 2.680 ;
        RECT 2474.210 1.630 2479.070 2.680 ;
        RECT 2480.190 1.630 2485.050 2.680 ;
        RECT 2486.170 1.630 2490.570 2.680 ;
        RECT 2491.690 1.630 2496.550 2.680 ;
        RECT 2497.670 1.630 2502.530 2.680 ;
        RECT 2503.650 1.630 2508.510 2.680 ;
        RECT 2509.630 1.630 2514.490 2.680 ;
        RECT 2515.610 1.630 2520.470 2.680 ;
        RECT 2521.590 1.630 2526.450 2.680 ;
        RECT 2527.570 1.630 2531.970 2.680 ;
        RECT 2533.090 1.630 2537.950 2.680 ;
        RECT 2539.070 1.630 2543.930 2.680 ;
        RECT 2545.050 1.630 2549.910 2.680 ;
        RECT 2551.030 1.630 2555.890 2.680 ;
        RECT 2557.010 1.630 2561.870 2.680 ;
        RECT 2562.990 1.630 2567.390 2.680 ;
        RECT 2568.510 1.630 2573.370 2.680 ;
        RECT 2574.490 1.630 2579.350 2.680 ;
        RECT 2580.470 1.630 2585.330 2.680 ;
        RECT 2586.450 1.630 2591.310 2.680 ;
        RECT 2592.430 1.630 2597.290 2.680 ;
        RECT 2598.410 1.630 2603.270 2.680 ;
        RECT 2604.390 1.630 2608.790 2.680 ;
        RECT 2609.910 1.630 2614.770 2.680 ;
        RECT 2615.890 1.630 2620.750 2.680 ;
        RECT 2621.870 1.630 2626.730 2.680 ;
        RECT 2627.850 1.630 2632.710 2.680 ;
        RECT 2633.830 1.630 2638.690 2.680 ;
        RECT 2639.810 1.630 2644.670 2.680 ;
        RECT 2645.790 1.630 2650.190 2.680 ;
        RECT 2651.310 1.630 2656.170 2.680 ;
        RECT 2657.290 1.630 2662.150 2.680 ;
        RECT 2663.270 1.630 2668.130 2.680 ;
        RECT 2669.250 1.630 2674.110 2.680 ;
        RECT 2675.230 1.630 2680.090 2.680 ;
        RECT 2681.210 1.630 2685.610 2.680 ;
        RECT 2686.730 1.630 2691.590 2.680 ;
        RECT 2692.710 1.630 2697.570 2.680 ;
        RECT 2698.690 1.630 2703.550 2.680 ;
        RECT 2704.670 1.630 2709.530 2.680 ;
        RECT 2710.650 1.630 2715.510 2.680 ;
        RECT 2716.630 1.630 2721.490 2.680 ;
        RECT 2722.610 1.630 2727.010 2.680 ;
        RECT 2728.130 1.630 2732.990 2.680 ;
        RECT 2734.110 1.630 2738.970 2.680 ;
        RECT 2740.090 1.630 2744.950 2.680 ;
        RECT 2746.070 1.630 2750.930 2.680 ;
        RECT 2752.050 1.630 2756.910 2.680 ;
        RECT 2758.030 1.630 2762.890 2.680 ;
        RECT 2764.010 1.630 2768.410 2.680 ;
        RECT 2769.530 1.630 2774.390 2.680 ;
        RECT 2775.510 1.630 2780.370 2.680 ;
        RECT 2781.490 1.630 2786.350 2.680 ;
        RECT 2787.470 1.630 2792.330 2.680 ;
        RECT 2793.450 1.630 2798.310 2.680 ;
        RECT 2799.430 1.630 2803.830 2.680 ;
        RECT 2804.950 1.630 2809.810 2.680 ;
        RECT 2810.930 1.630 2815.790 2.680 ;
        RECT 2816.910 1.630 2821.770 2.680 ;
        RECT 2822.890 1.630 2827.750 2.680 ;
        RECT 2828.870 1.630 2833.730 2.680 ;
        RECT 2834.850 1.630 2839.710 2.680 ;
        RECT 2840.830 1.630 2845.230 2.680 ;
        RECT 2846.350 1.630 2851.210 2.680 ;
        RECT 2852.330 1.630 2857.190 2.680 ;
        RECT 2858.310 1.630 2863.170 2.680 ;
        RECT 2864.290 1.630 2869.150 2.680 ;
        RECT 2870.270 1.630 2875.130 2.680 ;
        RECT 2876.250 1.630 2881.110 2.680 ;
        RECT 2882.230 1.630 2886.630 2.680 ;
        RECT 2887.750 1.630 2892.610 2.680 ;
        RECT 2893.730 1.630 2898.590 2.680 ;
        RECT 2899.710 1.630 2904.570 2.680 ;
        RECT 2905.690 1.630 2910.550 2.680 ;
        RECT 2911.670 1.630 2916.530 2.680 ;
      LAYER met3 ;
        RECT 2.400 3487.700 2917.600 3499.105 ;
        RECT 2.800 3487.020 2917.600 3487.700 ;
        RECT 2.800 3485.700 2917.200 3487.020 ;
        RECT 2.400 3485.020 2917.200 3485.700 ;
        RECT 2.400 3422.420 2917.600 3485.020 ;
        RECT 2.800 3420.420 2917.600 3422.420 ;
        RECT 2.400 3420.380 2917.600 3420.420 ;
        RECT 2.400 3418.380 2917.200 3420.380 ;
        RECT 2.400 3357.140 2917.600 3418.380 ;
        RECT 2.800 3355.140 2917.600 3357.140 ;
        RECT 2.400 3354.420 2917.600 3355.140 ;
        RECT 2.400 3352.420 2917.200 3354.420 ;
        RECT 2.400 3291.860 2917.600 3352.420 ;
        RECT 2.800 3289.860 2917.600 3291.860 ;
        RECT 2.400 3287.780 2917.600 3289.860 ;
        RECT 2.400 3285.780 2917.200 3287.780 ;
        RECT 2.400 3226.580 2917.600 3285.780 ;
        RECT 2.800 3224.580 2917.600 3226.580 ;
        RECT 2.400 3221.140 2917.600 3224.580 ;
        RECT 2.400 3219.140 2917.200 3221.140 ;
        RECT 2.400 3161.300 2917.600 3219.140 ;
        RECT 2.800 3159.300 2917.600 3161.300 ;
        RECT 2.400 3155.180 2917.600 3159.300 ;
        RECT 2.400 3153.180 2917.200 3155.180 ;
        RECT 2.400 3096.700 2917.600 3153.180 ;
        RECT 2.800 3094.700 2917.600 3096.700 ;
        RECT 2.400 3088.540 2917.600 3094.700 ;
        RECT 2.400 3086.540 2917.200 3088.540 ;
        RECT 2.400 3031.420 2917.600 3086.540 ;
        RECT 2.800 3029.420 2917.600 3031.420 ;
        RECT 2.400 3021.900 2917.600 3029.420 ;
        RECT 2.400 3019.900 2917.200 3021.900 ;
        RECT 2.400 2966.140 2917.600 3019.900 ;
        RECT 2.800 2964.140 2917.600 2966.140 ;
        RECT 2.400 2955.940 2917.600 2964.140 ;
        RECT 2.400 2953.940 2917.200 2955.940 ;
        RECT 2.400 2900.860 2917.600 2953.940 ;
        RECT 2.800 2898.860 2917.600 2900.860 ;
        RECT 2.400 2889.300 2917.600 2898.860 ;
        RECT 2.400 2887.300 2917.200 2889.300 ;
        RECT 2.400 2835.580 2917.600 2887.300 ;
        RECT 2.800 2833.580 2917.600 2835.580 ;
        RECT 2.400 2822.660 2917.600 2833.580 ;
        RECT 2.400 2820.660 2917.200 2822.660 ;
        RECT 2.400 2770.300 2917.600 2820.660 ;
        RECT 2.800 2768.300 2917.600 2770.300 ;
        RECT 2.400 2756.700 2917.600 2768.300 ;
        RECT 2.400 2754.700 2917.200 2756.700 ;
        RECT 2.400 2705.020 2917.600 2754.700 ;
        RECT 2.800 2703.020 2917.600 2705.020 ;
        RECT 2.400 2690.060 2917.600 2703.020 ;
        RECT 2.400 2688.060 2917.200 2690.060 ;
        RECT 2.400 2640.420 2917.600 2688.060 ;
        RECT 2.800 2638.420 2917.600 2640.420 ;
        RECT 2.400 2623.420 2917.600 2638.420 ;
        RECT 2.400 2621.420 2917.200 2623.420 ;
        RECT 2.400 2575.140 2917.600 2621.420 ;
        RECT 2.800 2573.140 2917.600 2575.140 ;
        RECT 2.400 2557.460 2917.600 2573.140 ;
        RECT 2.400 2555.460 2917.200 2557.460 ;
        RECT 2.400 2509.860 2917.600 2555.460 ;
        RECT 2.800 2507.860 2917.600 2509.860 ;
        RECT 2.400 2490.820 2917.600 2507.860 ;
        RECT 2.400 2488.820 2917.200 2490.820 ;
        RECT 2.400 2444.580 2917.600 2488.820 ;
        RECT 2.800 2442.580 2917.600 2444.580 ;
        RECT 2.400 2424.180 2917.600 2442.580 ;
        RECT 2.400 2422.180 2917.200 2424.180 ;
        RECT 2.400 2379.300 2917.600 2422.180 ;
        RECT 2.800 2377.300 2917.600 2379.300 ;
        RECT 2.400 2358.220 2917.600 2377.300 ;
        RECT 2.400 2356.220 2917.200 2358.220 ;
        RECT 2.400 2314.020 2917.600 2356.220 ;
        RECT 2.800 2312.020 2917.600 2314.020 ;
        RECT 2.400 2291.580 2917.600 2312.020 ;
        RECT 2.400 2289.580 2917.200 2291.580 ;
        RECT 2.400 2248.740 2917.600 2289.580 ;
        RECT 2.800 2246.740 2917.600 2248.740 ;
        RECT 2.400 2224.940 2917.600 2246.740 ;
        RECT 2.400 2222.940 2917.200 2224.940 ;
        RECT 2.400 2184.140 2917.600 2222.940 ;
        RECT 2.800 2182.140 2917.600 2184.140 ;
        RECT 2.400 2158.980 2917.600 2182.140 ;
        RECT 2.400 2156.980 2917.200 2158.980 ;
        RECT 2.400 2118.860 2917.600 2156.980 ;
        RECT 2.800 2116.860 2917.600 2118.860 ;
        RECT 2.400 2092.340 2917.600 2116.860 ;
        RECT 2.400 2090.340 2917.200 2092.340 ;
        RECT 2.400 2053.580 2917.600 2090.340 ;
        RECT 2.800 2051.580 2917.600 2053.580 ;
        RECT 2.400 2025.700 2917.600 2051.580 ;
        RECT 2.400 2023.700 2917.200 2025.700 ;
        RECT 2.400 1988.300 2917.600 2023.700 ;
        RECT 2.800 1986.300 2917.600 1988.300 ;
        RECT 2.400 1959.740 2917.600 1986.300 ;
        RECT 2.400 1957.740 2917.200 1959.740 ;
        RECT 2.400 1923.020 2917.600 1957.740 ;
        RECT 2.800 1921.020 2917.600 1923.020 ;
        RECT 2.400 1893.100 2917.600 1921.020 ;
        RECT 2.400 1891.100 2917.200 1893.100 ;
        RECT 2.400 1857.740 2917.600 1891.100 ;
        RECT 2.800 1855.740 2917.600 1857.740 ;
        RECT 2.400 1826.460 2917.600 1855.740 ;
        RECT 2.400 1824.460 2917.200 1826.460 ;
        RECT 2.400 1793.140 2917.600 1824.460 ;
        RECT 2.800 1791.140 2917.600 1793.140 ;
        RECT 2.400 1760.500 2917.600 1791.140 ;
        RECT 2.400 1758.500 2917.200 1760.500 ;
        RECT 2.400 1727.860 2917.600 1758.500 ;
        RECT 2.800 1725.860 2917.600 1727.860 ;
        RECT 2.400 1693.860 2917.600 1725.860 ;
        RECT 2.400 1691.860 2917.200 1693.860 ;
        RECT 2.400 1662.580 2917.600 1691.860 ;
        RECT 2.800 1660.580 2917.600 1662.580 ;
        RECT 2.400 1627.220 2917.600 1660.580 ;
        RECT 2.400 1625.220 2917.200 1627.220 ;
        RECT 2.400 1597.300 2917.600 1625.220 ;
        RECT 2.800 1595.300 2917.600 1597.300 ;
        RECT 2.400 1561.260 2917.600 1595.300 ;
        RECT 2.400 1559.260 2917.200 1561.260 ;
        RECT 2.400 1532.020 2917.600 1559.260 ;
        RECT 2.800 1530.020 2917.600 1532.020 ;
        RECT 2.400 1494.620 2917.600 1530.020 ;
        RECT 2.400 1492.620 2917.200 1494.620 ;
        RECT 2.400 1466.740 2917.600 1492.620 ;
        RECT 2.800 1464.740 2917.600 1466.740 ;
        RECT 2.400 1427.980 2917.600 1464.740 ;
        RECT 2.400 1425.980 2917.200 1427.980 ;
        RECT 2.400 1401.460 2917.600 1425.980 ;
        RECT 2.800 1399.460 2917.600 1401.460 ;
        RECT 2.400 1362.020 2917.600 1399.460 ;
        RECT 2.400 1360.020 2917.200 1362.020 ;
        RECT 2.400 1336.860 2917.600 1360.020 ;
        RECT 2.800 1334.860 2917.600 1336.860 ;
        RECT 2.400 1295.380 2917.600 1334.860 ;
        RECT 2.400 1293.380 2917.200 1295.380 ;
        RECT 2.400 1271.580 2917.600 1293.380 ;
        RECT 2.800 1269.580 2917.600 1271.580 ;
        RECT 2.400 1228.740 2917.600 1269.580 ;
        RECT 2.400 1226.740 2917.200 1228.740 ;
        RECT 2.400 1206.300 2917.600 1226.740 ;
        RECT 2.800 1204.300 2917.600 1206.300 ;
        RECT 2.400 1162.780 2917.600 1204.300 ;
        RECT 2.400 1160.780 2917.200 1162.780 ;
        RECT 2.400 1141.020 2917.600 1160.780 ;
        RECT 2.800 1139.020 2917.600 1141.020 ;
        RECT 2.400 1096.140 2917.600 1139.020 ;
        RECT 2.400 1094.140 2917.200 1096.140 ;
        RECT 2.400 1075.740 2917.600 1094.140 ;
        RECT 2.800 1073.740 2917.600 1075.740 ;
        RECT 2.400 1029.500 2917.600 1073.740 ;
        RECT 2.400 1027.500 2917.200 1029.500 ;
        RECT 2.400 1010.460 2917.600 1027.500 ;
        RECT 2.800 1008.460 2917.600 1010.460 ;
        RECT 2.400 963.540 2917.600 1008.460 ;
        RECT 2.400 961.540 2917.200 963.540 ;
        RECT 2.400 945.180 2917.600 961.540 ;
        RECT 2.800 943.180 2917.600 945.180 ;
        RECT 2.400 896.900 2917.600 943.180 ;
        RECT 2.400 894.900 2917.200 896.900 ;
        RECT 2.400 880.580 2917.600 894.900 ;
        RECT 2.800 878.580 2917.600 880.580 ;
        RECT 2.400 830.260 2917.600 878.580 ;
        RECT 2.400 828.260 2917.200 830.260 ;
        RECT 2.400 815.300 2917.600 828.260 ;
        RECT 2.800 813.300 2917.600 815.300 ;
        RECT 2.400 764.300 2917.600 813.300 ;
        RECT 2.400 762.300 2917.200 764.300 ;
        RECT 2.400 750.020 2917.600 762.300 ;
        RECT 2.800 748.020 2917.600 750.020 ;
        RECT 2.400 697.660 2917.600 748.020 ;
        RECT 2.400 695.660 2917.200 697.660 ;
        RECT 2.400 684.740 2917.600 695.660 ;
        RECT 2.800 682.740 2917.600 684.740 ;
        RECT 2.400 631.020 2917.600 682.740 ;
        RECT 2.400 629.020 2917.200 631.020 ;
        RECT 2.400 619.460 2917.600 629.020 ;
        RECT 2.800 617.460 2917.600 619.460 ;
        RECT 2.400 565.060 2917.600 617.460 ;
        RECT 2.400 563.060 2917.200 565.060 ;
        RECT 2.400 554.180 2917.600 563.060 ;
        RECT 2.800 552.180 2917.600 554.180 ;
        RECT 2.400 498.420 2917.600 552.180 ;
        RECT 2.400 496.420 2917.200 498.420 ;
        RECT 2.400 488.900 2917.600 496.420 ;
        RECT 2.800 486.900 2917.600 488.900 ;
        RECT 2.400 431.780 2917.600 486.900 ;
        RECT 2.400 429.780 2917.200 431.780 ;
        RECT 2.400 424.300 2917.600 429.780 ;
        RECT 2.800 422.300 2917.600 424.300 ;
        RECT 2.400 365.820 2917.600 422.300 ;
        RECT 2.400 363.820 2917.200 365.820 ;
        RECT 2.400 359.020 2917.600 363.820 ;
        RECT 2.800 357.020 2917.600 359.020 ;
        RECT 2.400 299.180 2917.600 357.020 ;
        RECT 2.400 297.180 2917.200 299.180 ;
        RECT 2.400 293.740 2917.600 297.180 ;
        RECT 2.800 291.740 2917.600 293.740 ;
        RECT 2.400 232.540 2917.600 291.740 ;
        RECT 2.400 230.540 2917.200 232.540 ;
        RECT 2.400 228.460 2917.600 230.540 ;
        RECT 2.800 226.460 2917.600 228.460 ;
        RECT 2.400 166.580 2917.600 226.460 ;
        RECT 2.400 164.580 2917.200 166.580 ;
        RECT 2.400 163.180 2917.600 164.580 ;
        RECT 2.800 161.180 2917.600 163.180 ;
        RECT 2.400 99.940 2917.600 161.180 ;
        RECT 2.400 97.940 2917.200 99.940 ;
        RECT 2.400 97.900 2917.600 97.940 ;
        RECT 2.800 95.900 2917.600 97.900 ;
        RECT 2.400 33.980 2917.600 95.900 ;
        RECT 2.400 33.300 2917.200 33.980 ;
        RECT 2.800 31.980 2917.200 33.300 ;
        RECT 2.800 31.300 2917.600 31.980 ;
        RECT 2.400 16.495 2917.600 31.300 ;
      LAYER met4 ;
        RECT 16.855 16.495 31.070 3499.105 ;
        RECT 34.970 16.495 53.570 3499.105 ;
        RECT 57.470 16.495 76.070 3499.105 ;
        RECT 79.970 16.495 98.570 3499.105 ;
        RECT 102.470 16.495 121.070 3499.105 ;
        RECT 124.970 16.495 143.570 3499.105 ;
        RECT 147.470 16.495 166.070 3499.105 ;
        RECT 169.970 16.495 188.570 3499.105 ;
        RECT 192.470 16.495 211.070 3499.105 ;
        RECT 214.970 1243.020 233.570 3499.105 ;
        RECT 237.470 1243.020 256.070 3499.105 ;
        RECT 259.970 1243.020 278.570 3499.105 ;
        RECT 282.470 1243.020 301.070 3499.105 ;
        RECT 304.970 1243.020 323.570 3499.105 ;
        RECT 327.470 1243.020 346.070 3499.105 ;
        RECT 349.970 1243.020 368.570 3499.105 ;
        RECT 372.470 1243.020 391.070 3499.105 ;
        RECT 394.970 1243.020 413.570 3499.105 ;
        RECT 417.470 1243.020 436.070 3499.105 ;
        RECT 439.970 1243.020 458.570 3499.105 ;
        RECT 462.470 1243.020 481.070 3499.105 ;
        RECT 484.970 1243.020 503.570 3499.105 ;
        RECT 507.470 1243.020 526.070 3499.105 ;
        RECT 529.970 1243.020 548.570 3499.105 ;
        RECT 552.470 1243.020 571.070 3499.105 ;
        RECT 574.970 1243.020 593.570 3499.105 ;
        RECT 597.470 1243.020 616.070 3499.105 ;
        RECT 619.970 1243.020 638.570 3499.105 ;
        RECT 642.470 1243.020 661.070 3499.105 ;
        RECT 664.970 1243.020 683.570 3499.105 ;
        RECT 687.470 1243.020 706.070 3499.105 ;
        RECT 709.970 1243.020 728.570 3499.105 ;
        RECT 732.470 1243.020 751.070 3499.105 ;
        RECT 754.970 1243.020 773.570 3499.105 ;
        RECT 777.470 1243.020 796.070 3499.105 ;
        RECT 799.970 1243.020 818.570 3499.105 ;
        RECT 822.470 1243.020 841.070 3499.105 ;
        RECT 844.970 1243.020 863.570 3499.105 ;
        RECT 867.470 1243.020 886.070 3499.105 ;
        RECT 889.970 1243.020 908.570 3499.105 ;
        RECT 912.470 1243.020 931.070 3499.105 ;
        RECT 934.970 1243.020 953.570 3499.105 ;
        RECT 957.470 1243.020 976.070 3499.105 ;
        RECT 979.970 1243.020 998.570 3499.105 ;
        RECT 1002.470 1243.020 1021.070 3499.105 ;
        RECT 1024.970 1243.020 1043.570 3499.105 ;
        RECT 1047.470 1243.020 1066.070 3499.105 ;
        RECT 1069.970 1243.020 1088.570 3499.105 ;
        RECT 1092.470 1243.020 1111.070 3499.105 ;
        RECT 1114.970 1243.020 1133.570 3499.105 ;
        RECT 1137.470 1243.020 1156.070 3499.105 ;
        RECT 1159.970 1243.020 1178.570 3499.105 ;
        RECT 1182.470 1243.020 1201.070 3499.105 ;
        RECT 1204.970 1243.020 1223.570 3499.105 ;
        RECT 1227.470 1243.020 1246.070 3499.105 ;
        RECT 1249.970 1243.020 1268.570 3499.105 ;
        RECT 1272.470 1243.020 1291.070 3499.105 ;
        RECT 1294.970 1243.020 1313.570 3499.105 ;
        RECT 1317.470 1243.020 1336.070 3499.105 ;
        RECT 1339.970 1243.020 1358.570 3499.105 ;
        RECT 1362.470 1243.020 1381.070 3499.105 ;
        RECT 1384.970 1243.020 1403.570 3499.105 ;
        RECT 1407.470 1243.020 1426.070 3499.105 ;
        RECT 1429.970 1243.020 1448.570 3499.105 ;
        RECT 1452.470 1243.020 1471.070 3499.105 ;
        RECT 1474.970 1243.020 1493.570 3499.105 ;
        RECT 1497.470 1243.020 1516.070 3499.105 ;
        RECT 1519.970 1243.020 1538.570 3499.105 ;
        RECT 1542.470 1243.020 1561.070 3499.105 ;
        RECT 1564.970 1243.020 1583.570 3499.105 ;
        RECT 1587.470 1243.020 1606.070 3499.105 ;
        RECT 1609.970 1243.020 1628.570 3499.105 ;
        RECT 1632.470 1243.020 1651.070 3499.105 ;
        RECT 1654.970 1243.020 1673.570 3499.105 ;
        RECT 1677.470 1243.020 1696.070 3499.105 ;
        RECT 1699.970 1243.020 1718.570 3499.105 ;
        RECT 1722.470 1243.020 1741.070 3499.105 ;
        RECT 1744.970 1243.020 1763.570 3499.105 ;
        RECT 1767.470 1243.020 1786.070 3499.105 ;
        RECT 1789.970 1243.020 1808.570 3499.105 ;
        RECT 1812.470 1243.020 1831.070 3499.105 ;
        RECT 1834.970 1243.020 1853.570 3499.105 ;
        RECT 1857.470 1243.020 1876.070 3499.105 ;
        RECT 1879.970 1243.020 1898.570 3499.105 ;
        RECT 1902.470 1243.020 1921.070 3499.105 ;
        RECT 1924.970 1243.020 1943.570 3499.105 ;
        RECT 1947.470 1243.020 1966.070 3499.105 ;
        RECT 1969.970 1243.020 1988.570 3499.105 ;
        RECT 1992.470 1243.020 2011.070 3499.105 ;
        RECT 214.970 1142.820 2011.070 1243.020 ;
        RECT 214.970 16.495 233.570 1142.820 ;
        RECT 237.470 16.495 256.070 1142.820 ;
        RECT 259.970 16.495 278.570 1142.820 ;
        RECT 282.470 16.495 301.070 1142.820 ;
        RECT 304.970 16.495 323.570 1142.820 ;
        RECT 327.470 16.495 346.070 1142.820 ;
        RECT 349.970 16.495 368.570 1142.820 ;
        RECT 372.470 16.495 391.070 1142.820 ;
        RECT 394.970 16.495 413.570 1142.820 ;
        RECT 417.470 16.495 436.070 1142.820 ;
        RECT 439.970 16.495 458.570 1142.820 ;
        RECT 462.470 16.495 481.070 1142.820 ;
        RECT 484.970 16.495 503.570 1142.820 ;
        RECT 507.470 16.495 526.070 1142.820 ;
        RECT 529.970 16.495 548.570 1142.820 ;
        RECT 552.470 684.600 571.070 1142.820 ;
        RECT 574.970 684.600 593.570 1142.820 ;
        RECT 597.470 684.600 616.070 1142.820 ;
        RECT 619.970 684.600 638.570 1142.820 ;
        RECT 642.470 684.600 661.070 1142.820 ;
        RECT 664.970 684.600 863.570 1142.820 ;
        RECT 867.470 684.600 886.070 1142.820 ;
        RECT 889.970 684.600 908.570 1142.820 ;
        RECT 552.470 365.400 908.570 684.600 ;
        RECT 552.470 16.495 571.070 365.400 ;
        RECT 574.970 16.495 593.570 365.400 ;
        RECT 597.470 16.495 616.070 365.400 ;
        RECT 619.970 16.495 638.570 365.400 ;
        RECT 642.470 16.495 661.070 365.400 ;
        RECT 664.970 16.495 683.570 365.400 ;
        RECT 687.470 16.495 706.070 365.400 ;
        RECT 709.970 16.495 728.570 365.400 ;
        RECT 732.470 16.495 751.070 365.400 ;
        RECT 754.970 16.495 773.570 365.400 ;
        RECT 777.470 16.495 796.070 365.400 ;
        RECT 799.970 16.495 818.570 365.400 ;
        RECT 822.470 16.495 841.070 365.400 ;
        RECT 844.970 16.495 863.570 365.400 ;
        RECT 867.470 16.495 886.070 365.400 ;
        RECT 889.970 16.495 908.570 365.400 ;
        RECT 912.470 16.495 931.070 1142.820 ;
        RECT 934.970 16.495 953.570 1142.820 ;
        RECT 957.470 16.495 976.070 1142.820 ;
        RECT 979.970 16.495 998.570 1142.820 ;
        RECT 1002.470 16.495 1021.070 1142.820 ;
        RECT 1024.970 16.495 1043.570 1142.820 ;
        RECT 1047.470 16.495 1066.070 1142.820 ;
        RECT 1069.970 16.495 1088.570 1142.820 ;
        RECT 1092.470 16.495 1111.070 1142.820 ;
        RECT 1114.970 16.495 1133.570 1142.820 ;
        RECT 1137.470 16.495 1156.070 1142.820 ;
        RECT 1159.970 16.495 1178.570 1142.820 ;
        RECT 1182.470 16.495 1201.070 1142.820 ;
        RECT 1204.970 16.495 1223.570 1142.820 ;
        RECT 1227.470 16.495 1246.070 1142.820 ;
        RECT 1249.970 16.495 1268.570 1142.820 ;
        RECT 1272.470 16.495 1291.070 1142.820 ;
        RECT 1294.970 16.495 1313.570 1142.820 ;
        RECT 1317.470 16.495 1336.070 1142.820 ;
        RECT 1339.970 16.495 1358.570 1142.820 ;
        RECT 1362.470 16.495 1381.070 1142.820 ;
        RECT 1384.970 16.495 1403.570 1142.820 ;
        RECT 1407.470 16.495 1426.070 1142.820 ;
        RECT 1429.970 16.495 1448.570 1142.820 ;
        RECT 1452.470 16.495 1471.070 1142.820 ;
        RECT 1474.970 16.495 1493.570 1142.820 ;
        RECT 1497.470 16.495 1516.070 1142.820 ;
        RECT 1519.970 16.495 1538.570 1142.820 ;
        RECT 1542.470 16.495 1561.070 1142.820 ;
        RECT 1564.970 16.495 1583.570 1142.820 ;
        RECT 1587.470 16.495 1606.070 1142.820 ;
        RECT 1609.970 16.495 1628.570 1142.820 ;
        RECT 1632.470 16.495 1651.070 1142.820 ;
        RECT 1654.970 16.495 1673.570 1142.820 ;
        RECT 1677.470 16.495 1696.070 1142.820 ;
        RECT 1699.970 16.495 1718.570 1142.820 ;
        RECT 1722.470 16.495 1741.070 1142.820 ;
        RECT 1744.970 16.495 1763.570 1142.820 ;
        RECT 1767.470 16.495 1786.070 1142.820 ;
        RECT 1789.970 16.495 1808.570 1142.820 ;
        RECT 1812.470 16.495 1831.070 1142.820 ;
        RECT 1834.970 16.495 1853.570 1142.820 ;
        RECT 1857.470 16.495 1876.070 1142.820 ;
        RECT 1879.970 16.495 1898.570 1142.820 ;
        RECT 1902.470 16.495 1921.070 1142.820 ;
        RECT 1924.970 16.495 1943.570 1142.820 ;
        RECT 1947.470 16.495 1966.070 1142.820 ;
        RECT 1969.970 16.495 1988.570 1142.820 ;
        RECT 1992.470 16.495 2011.070 1142.820 ;
        RECT 2014.970 16.495 2033.570 3499.105 ;
        RECT 2037.470 16.495 2056.070 3499.105 ;
        RECT 2059.970 16.495 2078.570 3499.105 ;
        RECT 2082.470 16.495 2101.070 3499.105 ;
        RECT 2104.970 16.495 2123.570 3499.105 ;
        RECT 2127.470 16.495 2146.070 3499.105 ;
        RECT 2149.970 16.495 2168.570 3499.105 ;
        RECT 2172.470 16.495 2191.070 3499.105 ;
        RECT 2194.970 16.495 2213.570 3499.105 ;
        RECT 2217.470 16.495 2236.070 3499.105 ;
        RECT 2239.970 16.495 2258.570 3499.105 ;
        RECT 2262.470 16.495 2281.070 3499.105 ;
        RECT 2284.970 16.495 2303.570 3499.105 ;
        RECT 2307.470 16.495 2326.070 3499.105 ;
        RECT 2329.970 16.495 2348.570 3499.105 ;
        RECT 2352.470 16.495 2371.070 3499.105 ;
        RECT 2374.970 16.495 2393.570 3499.105 ;
        RECT 2397.470 16.495 2416.070 3499.105 ;
        RECT 2419.970 16.495 2438.570 3499.105 ;
        RECT 2442.470 16.495 2461.070 3499.105 ;
        RECT 2464.970 16.495 2483.570 3499.105 ;
        RECT 2487.470 16.495 2506.070 3499.105 ;
        RECT 2509.970 16.495 2528.570 3499.105 ;
        RECT 2532.470 16.495 2551.070 3499.105 ;
        RECT 2554.970 16.495 2573.570 3499.105 ;
        RECT 2577.470 16.495 2596.070 3499.105 ;
        RECT 2599.970 16.495 2618.570 3499.105 ;
        RECT 2622.470 16.495 2641.070 3499.105 ;
        RECT 2644.970 16.495 2663.570 3499.105 ;
        RECT 2667.470 16.495 2686.070 3499.105 ;
        RECT 2689.970 1603.600 2708.570 3499.105 ;
        RECT 2712.470 1603.600 2731.070 3499.105 ;
        RECT 2734.970 1603.600 2753.570 3499.105 ;
        RECT 2757.470 1603.600 2776.070 3499.105 ;
        RECT 2779.970 1603.600 2798.570 3499.105 ;
        RECT 2802.470 1603.600 2821.070 3499.105 ;
        RECT 2824.970 1603.600 2843.570 3499.105 ;
        RECT 2847.470 1603.600 2866.070 3499.105 ;
        RECT 2689.970 1500.400 2866.070 1603.600 ;
        RECT 2689.970 16.495 2708.570 1500.400 ;
        RECT 2712.470 16.495 2731.070 1500.400 ;
        RECT 2734.970 16.495 2753.570 1500.400 ;
        RECT 2757.470 16.495 2776.070 1500.400 ;
        RECT 2779.970 16.495 2798.570 1500.400 ;
        RECT 2802.470 16.495 2821.070 1500.400 ;
        RECT 2824.970 16.495 2843.570 1500.400 ;
        RECT 2847.470 16.495 2866.070 1500.400 ;
        RECT 2869.970 16.495 2888.570 3499.105 ;
        RECT 2892.470 16.495 2901.385 3499.105 ;
  END
END user_project_wrapper
END LIBRARY

