magic
tech sky130B
magscale 1 2
timestamp 1668033750
<< metal1 >>
rect 201494 702992 201500 703044
rect 201552 703032 201558 703044
rect 202782 703032 202788 703044
rect 201552 703004 202788 703032
rect 201552 702992 201558 703004
rect 202782 702992 202788 703004
rect 202840 702992 202846 703044
rect 331214 702992 331220 703044
rect 331272 703032 331278 703044
rect 332502 703032 332508 703044
rect 331272 703004 332508 703032
rect 331272 702992 331278 703004
rect 332502 702992 332508 703004
rect 332560 702992 332566 703044
rect 207658 700612 207664 700664
rect 207716 700652 207722 700664
rect 218974 700652 218980 700664
rect 207716 700624 218980 700652
rect 207716 700612 207722 700624
rect 218974 700612 218980 700624
rect 219032 700612 219038 700664
rect 206278 700544 206284 700596
rect 206336 700584 206342 700596
rect 283834 700584 283840 700596
rect 206336 700556 283840 700584
rect 206336 700544 206342 700556
rect 283834 700544 283840 700556
rect 283892 700544 283898 700596
rect 203518 700476 203524 700528
rect 203576 700516 203582 700528
rect 348786 700516 348792 700528
rect 203576 700488 348792 700516
rect 203576 700476 203582 700488
rect 348786 700476 348792 700488
rect 348844 700476 348850 700528
rect 154114 700408 154120 700460
rect 154172 700448 154178 700460
rect 189074 700448 189080 700460
rect 154172 700420 189080 700448
rect 154172 700408 154178 700420
rect 189074 700408 189080 700420
rect 189132 700408 189138 700460
rect 200758 700408 200764 700460
rect 200816 700448 200822 700460
rect 413646 700448 413652 700460
rect 200816 700420 413652 700448
rect 200816 700408 200822 700420
rect 413646 700408 413652 700420
rect 413704 700408 413710 700460
rect 72970 700340 72976 700392
rect 73028 700380 73034 700392
rect 119338 700380 119344 700392
rect 73028 700352 119344 700380
rect 73028 700340 73034 700352
rect 119338 700340 119344 700352
rect 119396 700340 119402 700392
rect 137830 700340 137836 700392
rect 137888 700380 137894 700392
rect 189350 700380 189356 700392
rect 137888 700352 189356 700380
rect 137888 700340 137894 700352
rect 189350 700340 189356 700352
rect 189408 700340 189414 700392
rect 199378 700340 199384 700392
rect 199436 700380 199442 700392
rect 478506 700380 478512 700392
rect 199436 700352 478512 700380
rect 199436 700340 199442 700352
rect 478506 700340 478512 700352
rect 478564 700340 478570 700392
rect 24302 700272 24308 700324
rect 24360 700312 24366 700324
rect 189166 700312 189172 700324
rect 24360 700284 189172 700312
rect 24360 700272 24366 700284
rect 189166 700272 189172 700284
rect 189224 700272 189230 700324
rect 197998 700272 198004 700324
rect 198056 700312 198062 700324
rect 543458 700312 543464 700324
rect 198056 700284 543464 700312
rect 198056 700272 198062 700284
rect 543458 700272 543464 700284
rect 543516 700272 543522 700324
rect 105446 699660 105452 699712
rect 105504 699700 105510 699712
rect 106918 699700 106924 699712
rect 105504 699672 106924 699700
rect 105504 699660 105510 699672
rect 106918 699660 106924 699672
rect 106976 699660 106982 699712
rect 266354 697552 266360 697604
rect 266412 697592 266418 697604
rect 267642 697592 267648 697604
rect 266412 697564 267648 697592
rect 266412 697552 266418 697564
rect 267642 697552 267648 697564
rect 267700 697552 267706 697604
rect 2774 683612 2780 683664
rect 2832 683652 2838 683664
rect 6178 683652 6184 683664
rect 2832 683624 6184 683652
rect 2832 683612 2838 683624
rect 6178 683612 6184 683624
rect 6236 683612 6242 683664
rect 196618 683136 196624 683188
rect 196676 683176 196682 683188
rect 579614 683176 579620 683188
rect 196676 683148 579620 683176
rect 196676 683136 196682 683148
rect 579614 683136 579620 683148
rect 579672 683136 579678 683188
rect 3418 670760 3424 670812
rect 3476 670800 3482 670812
rect 189258 670800 189264 670812
rect 3476 670772 189264 670800
rect 3476 670760 3482 670772
rect 189258 670760 189264 670772
rect 189316 670760 189322 670812
rect 120718 670692 120724 670744
rect 120776 670732 120782 670744
rect 580166 670732 580172 670744
rect 120776 670704 580172 670732
rect 120776 670692 120782 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 191098 643084 191104 643136
rect 191156 643124 191162 643136
rect 580166 643124 580172 643136
rect 191156 643096 580172 643124
rect 191156 643084 191162 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 2774 632068 2780 632120
rect 2832 632108 2838 632120
rect 4798 632108 4804 632120
rect 2832 632080 4804 632108
rect 2832 632068 2838 632080
rect 4798 632068 4804 632080
rect 4856 632068 4862 632120
rect 193858 630640 193864 630692
rect 193916 630680 193922 630692
rect 579982 630680 579988 630692
rect 193916 630652 579988 630680
rect 193916 630640 193922 630652
rect 579982 630640 579988 630652
rect 580040 630640 580046 630692
rect 3510 618264 3516 618316
rect 3568 618304 3574 618316
rect 190454 618304 190460 618316
rect 3568 618276 190460 618304
rect 3568 618264 3574 618276
rect 190454 618264 190460 618276
rect 190512 618264 190518 618316
rect 118694 616836 118700 616888
rect 118752 616876 118758 616888
rect 580166 616876 580172 616888
rect 118752 616848 580172 616876
rect 118752 616836 118758 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 192478 590656 192484 590708
rect 192536 590696 192542 590708
rect 580166 590696 580172 590708
rect 192536 590668 580172 590696
rect 192536 590656 192542 590668
rect 580166 590656 580172 590668
rect 580224 590656 580230 590708
rect 3142 579776 3148 579828
rect 3200 579816 3206 579828
rect 7558 579816 7564 579828
rect 3200 579788 7564 579816
rect 3200 579776 3206 579788
rect 7558 579776 7564 579788
rect 7616 579776 7622 579828
rect 193950 576852 193956 576904
rect 194008 576892 194014 576904
rect 580166 576892 580172 576904
rect 194008 576864 580172 576892
rect 194008 576852 194014 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 3050 565836 3056 565888
rect 3108 565876 3114 565888
rect 191834 565876 191840 565888
rect 3108 565848 191840 565876
rect 3108 565836 3114 565848
rect 191834 565836 191840 565848
rect 191892 565836 191898 565888
rect 120810 563048 120816 563100
rect 120868 563088 120874 563100
rect 580166 563088 580172 563100
rect 120868 563060 580172 563088
rect 120868 563048 120874 563060
rect 580166 563048 580172 563060
rect 580224 563048 580230 563100
rect 3326 553392 3332 553444
rect 3384 553432 3390 553444
rect 116578 553432 116584 553444
rect 3384 553404 116584 553432
rect 3384 553392 3390 553404
rect 116578 553392 116584 553404
rect 116636 553392 116642 553444
rect 192570 536800 192576 536852
rect 192628 536840 192634 536852
rect 579890 536840 579896 536852
rect 192628 536812 579896 536840
rect 192628 536800 192634 536812
rect 579890 536800 579896 536812
rect 579948 536800 579954 536852
rect 2958 527144 2964 527196
rect 3016 527184 3022 527196
rect 15838 527184 15844 527196
rect 3016 527156 15844 527184
rect 3016 527144 3022 527156
rect 15838 527144 15844 527156
rect 15896 527144 15902 527196
rect 194042 524424 194048 524476
rect 194100 524464 194106 524476
rect 580166 524464 580172 524476
rect 194100 524436 580172 524464
rect 194100 524424 194106 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 120902 510620 120908 510672
rect 120960 510660 120966 510672
rect 580166 510660 580172 510672
rect 120960 510632 580172 510660
rect 120960 510620 120966 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 3326 474716 3332 474768
rect 3384 474756 3390 474768
rect 19978 474756 19984 474768
rect 3384 474728 19984 474756
rect 3384 474716 3390 474728
rect 19978 474716 19984 474728
rect 20036 474716 20042 474768
rect 120994 456764 121000 456816
rect 121052 456804 121058 456816
rect 579614 456804 579620 456816
rect 121052 456776 579620 456804
rect 121052 456764 121058 456776
rect 579614 456764 579620 456776
rect 579672 456764 579678 456816
rect 2958 422288 2964 422340
rect 3016 422328 3022 422340
rect 22738 422328 22744 422340
rect 3016 422300 22744 422328
rect 3016 422288 3022 422300
rect 22738 422288 22744 422300
rect 22796 422288 22802 422340
rect 192662 418140 192668 418192
rect 192720 418180 192726 418192
rect 579706 418180 579712 418192
rect 192720 418152 579712 418180
rect 192720 418140 192726 418152
rect 579706 418140 579712 418152
rect 579764 418140 579770 418192
rect 3326 409844 3332 409896
rect 3384 409884 3390 409896
rect 189442 409884 189448 409896
rect 3384 409856 189448 409884
rect 3384 409844 3390 409856
rect 189442 409844 189448 409856
rect 189500 409844 189506 409896
rect 118602 404336 118608 404388
rect 118660 404376 118666 404388
rect 580166 404376 580172 404388
rect 118660 404348 580172 404376
rect 118660 404336 118666 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 192754 378156 192760 378208
rect 192812 378196 192818 378208
rect 580166 378196 580172 378208
rect 192812 378168 580172 378196
rect 192812 378156 192818 378168
rect 580166 378156 580172 378168
rect 580224 378156 580230 378208
rect 3326 371220 3332 371272
rect 3384 371260 3390 371272
rect 22830 371260 22836 371272
rect 3384 371232 22836 371260
rect 3384 371220 3390 371232
rect 22830 371220 22836 371232
rect 22888 371220 22894 371272
rect 366358 364352 366364 364404
rect 366416 364392 366422 364404
rect 580166 364392 580172 364404
rect 366416 364364 580172 364392
rect 366416 364352 366422 364364
rect 580166 364352 580172 364364
rect 580224 364352 580230 364404
rect 3326 357416 3332 357468
rect 3384 357456 3390 357468
rect 190546 357456 190552 357468
rect 3384 357428 190552 357456
rect 3384 357416 3390 357428
rect 190546 357416 190552 357428
rect 190604 357416 190610 357468
rect 118510 351908 118516 351960
rect 118568 351948 118574 351960
rect 580166 351948 580172 351960
rect 118568 351920 580172 351948
rect 118568 351908 118574 351920
rect 580166 351908 580172 351920
rect 580224 351908 580230 351960
rect 3326 345040 3332 345092
rect 3384 345080 3390 345092
rect 116670 345080 116676 345092
rect 3384 345052 116676 345080
rect 3384 345040 3390 345052
rect 116670 345040 116676 345052
rect 116728 345040 116734 345092
rect 2774 319064 2780 319116
rect 2832 319104 2838 319116
rect 4890 319104 4896 319116
rect 2832 319076 4896 319104
rect 2832 319064 2838 319076
rect 4890 319064 4896 319076
rect 4948 319064 4954 319116
rect 362218 311856 362224 311908
rect 362276 311896 362282 311908
rect 580166 311896 580172 311908
rect 362276 311868 580172 311896
rect 362276 311856 362282 311868
rect 580166 311856 580172 311868
rect 580224 311856 580230 311908
rect 2866 304988 2872 305040
rect 2924 305028 2930 305040
rect 188338 305028 188344 305040
rect 2924 305000 188344 305028
rect 2924 304988 2930 305000
rect 188338 304988 188344 305000
rect 188396 304988 188402 305040
rect 280798 298120 280804 298172
rect 280856 298160 280862 298172
rect 580166 298160 580172 298172
rect 280856 298132 580172 298160
rect 280856 298120 280862 298132
rect 580166 298120 580172 298132
rect 580224 298120 580230 298172
rect 3326 292544 3332 292596
rect 3384 292584 3390 292596
rect 79318 292584 79324 292596
rect 3384 292556 79324 292584
rect 3384 292544 3390 292556
rect 79318 292544 79324 292556
rect 79376 292544 79382 292596
rect 118786 275272 118792 275324
rect 118844 275312 118850 275324
rect 234614 275312 234620 275324
rect 118844 275284 234620 275312
rect 118844 275272 118850 275284
rect 234614 275272 234620 275284
rect 234672 275272 234678 275324
rect 192846 271872 192852 271924
rect 192904 271912 192910 271924
rect 580166 271912 580172 271924
rect 192904 271884 580172 271912
rect 192904 271872 192910 271884
rect 580166 271872 580172 271884
rect 580224 271872 580230 271924
rect 3234 266364 3240 266416
rect 3292 266404 3298 266416
rect 22922 266404 22928 266416
rect 3292 266376 22928 266404
rect 3292 266364 3298 266376
rect 22922 266364 22928 266376
rect 22980 266364 22986 266416
rect 531958 258068 531964 258120
rect 532016 258108 532022 258120
rect 579614 258108 579620 258120
rect 532016 258080 579620 258108
rect 532016 258068 532022 258080
rect 579614 258068 579620 258080
rect 579672 258068 579678 258120
rect 2866 253920 2872 253972
rect 2924 253960 2930 253972
rect 188430 253960 188436 253972
rect 2924 253932 188436 253960
rect 2924 253920 2930 253932
rect 188430 253920 188436 253932
rect 188488 253920 188494 253972
rect 360838 244264 360844 244316
rect 360896 244304 360902 244316
rect 580166 244304 580172 244316
rect 360896 244276 580172 244304
rect 360896 244264 360902 244276
rect 580166 244264 580172 244276
rect 580224 244264 580230 244316
rect 3234 240116 3240 240168
rect 3292 240156 3298 240168
rect 119430 240156 119436 240168
rect 3292 240128 119436 240156
rect 3292 240116 3298 240128
rect 119430 240116 119436 240128
rect 119488 240116 119494 240168
rect 118418 239368 118424 239420
rect 118476 239408 118482 239420
rect 280798 239408 280804 239420
rect 118476 239380 280804 239408
rect 118476 239368 118482 239380
rect 280798 239368 280804 239380
rect 280856 239368 280862 239420
rect 532050 218016 532056 218068
rect 532108 218056 532114 218068
rect 580166 218056 580172 218068
rect 532108 218028 580172 218056
rect 532108 218016 532114 218028
rect 580166 218016 580172 218028
rect 580224 218016 580230 218068
rect 3326 213936 3332 213988
rect 3384 213976 3390 213988
rect 24118 213976 24124 213988
rect 3384 213948 24124 213976
rect 3384 213936 3390 213948
rect 24118 213936 24124 213948
rect 24176 213936 24182 213988
rect 280798 205640 280804 205692
rect 280856 205680 280862 205692
rect 580166 205680 580172 205692
rect 280856 205652 580172 205680
rect 280856 205640 280862 205652
rect 580166 205640 580172 205652
rect 580224 205640 580230 205692
rect 118326 202104 118332 202156
rect 118384 202144 118390 202156
rect 360838 202144 360844 202156
rect 118384 202116 360844 202144
rect 118384 202104 118390 202116
rect 360838 202104 360844 202116
rect 360896 202104 360902 202156
rect 3326 201492 3332 201544
rect 3384 201532 3390 201544
rect 190730 201532 190736 201544
rect 3384 201504 190736 201532
rect 3384 201492 3390 201504
rect 190730 201492 190736 201504
rect 190788 201492 190794 201544
rect 196710 191836 196716 191888
rect 196768 191876 196774 191888
rect 580166 191876 580172 191888
rect 196768 191848 580172 191876
rect 196768 191836 196774 191848
rect 580166 191836 580172 191848
rect 580224 191836 580230 191888
rect 358078 178032 358084 178084
rect 358136 178072 358142 178084
rect 580166 178072 580172 178084
rect 358136 178044 580172 178072
rect 358136 178032 358142 178044
rect 580166 178032 580172 178044
rect 580224 178032 580230 178084
rect 122098 165588 122104 165640
rect 122156 165628 122162 165640
rect 579614 165628 579620 165640
rect 122156 165600 579620 165628
rect 122156 165588 122162 165600
rect 579614 165588 579620 165600
rect 579672 165588 579678 165640
rect 3326 162868 3332 162920
rect 3384 162908 3390 162920
rect 29638 162908 29644 162920
rect 3384 162880 29644 162908
rect 3384 162868 3390 162880
rect 29638 162868 29644 162880
rect 29696 162868 29702 162920
rect 196894 151784 196900 151836
rect 196952 151824 196958 151836
rect 579982 151824 579988 151836
rect 196952 151796 579988 151824
rect 196952 151784 196958 151796
rect 579982 151784 579988 151796
rect 580040 151784 580046 151836
rect 118878 149676 118884 149728
rect 118936 149716 118942 149728
rect 299474 149716 299480 149728
rect 118936 149688 299480 149716
rect 118936 149676 118942 149688
rect 299474 149676 299480 149688
rect 299532 149676 299538 149728
rect 3326 149064 3332 149116
rect 3384 149104 3390 149116
rect 189718 149104 189724 149116
rect 3384 149076 189724 149104
rect 3384 149064 3390 149076
rect 189718 149064 189724 149076
rect 189776 149064 189782 149116
rect 3970 148316 3976 148368
rect 4028 148356 4034 148368
rect 189626 148356 189632 148368
rect 4028 148328 189632 148356
rect 4028 148316 4034 148328
rect 189626 148316 189632 148328
rect 189684 148316 189690 148368
rect 3694 144168 3700 144220
rect 3752 144208 3758 144220
rect 190914 144208 190920 144220
rect 3752 144180 190920 144208
rect 3752 144168 3758 144180
rect 190914 144168 190920 144180
rect 190972 144168 190978 144220
rect 88334 142876 88340 142928
rect 88392 142916 88398 142928
rect 190822 142916 190828 142928
rect 88392 142888 190828 142916
rect 88392 142876 88398 142888
rect 190822 142876 190828 142888
rect 190880 142876 190886 142928
rect 118234 142808 118240 142860
rect 118292 142848 118298 142860
rect 280798 142848 280804 142860
rect 118292 142820 280804 142848
rect 118292 142808 118298 142820
rect 280798 142808 280804 142820
rect 280856 142808 280862 142860
rect 118050 141448 118056 141500
rect 118108 141488 118114 141500
rect 169754 141488 169760 141500
rect 118108 141460 169760 141488
rect 118108 141448 118114 141460
rect 169754 141448 169760 141460
rect 169812 141448 169818 141500
rect 119154 141380 119160 141432
rect 119212 141420 119218 141432
rect 429194 141420 429200 141432
rect 119212 141392 429200 141420
rect 119212 141380 119218 141392
rect 429194 141380 429200 141392
rect 429252 141380 429258 141432
rect 119246 140156 119252 140208
rect 119304 140196 119310 140208
rect 364334 140196 364340 140208
rect 119304 140168 364340 140196
rect 119304 140156 119310 140168
rect 364334 140156 364340 140168
rect 364392 140156 364398 140208
rect 119062 140088 119068 140140
rect 119120 140128 119126 140140
rect 494054 140128 494060 140140
rect 119120 140100 494060 140128
rect 119120 140088 119126 140100
rect 494054 140088 494060 140100
rect 494112 140088 494118 140140
rect 118970 140020 118976 140072
rect 119028 140060 119034 140072
rect 558914 140060 558920 140072
rect 119028 140032 558920 140060
rect 119028 140020 119034 140032
rect 558914 140020 558920 140032
rect 558972 140020 558978 140072
rect 118142 139408 118148 139460
rect 118200 139448 118206 139460
rect 122098 139448 122104 139460
rect 118200 139420 122104 139448
rect 118200 139408 118206 139420
rect 122098 139408 122104 139420
rect 122156 139408 122162 139460
rect 188338 139340 188344 139392
rect 188396 139380 188402 139392
rect 191926 139380 191932 139392
rect 188396 139352 191932 139380
rect 188396 139340 188402 139352
rect 191926 139340 191932 139352
rect 191984 139340 191990 139392
rect 188430 139272 188436 139324
rect 188488 139312 188494 139324
rect 192018 139312 192024 139324
rect 188488 139284 192024 139312
rect 188488 139272 188494 139284
rect 192018 139272 192024 139284
rect 192076 139272 192082 139324
rect 3694 137980 3700 138032
rect 3752 138020 3758 138032
rect 190638 138020 190644 138032
rect 3752 137992 190644 138020
rect 3752 137980 3758 137992
rect 190638 137980 190644 137992
rect 190696 137980 190702 138032
rect 2774 136688 2780 136740
rect 2832 136728 2838 136740
rect 4982 136728 4988 136740
rect 2832 136700 4988 136728
rect 2832 136688 2838 136700
rect 4982 136688 4988 136700
rect 5040 136688 5046 136740
rect 23014 136620 23020 136672
rect 23072 136660 23078 136672
rect 117314 136660 117320 136672
rect 23072 136632 117320 136660
rect 23072 136620 23078 136632
rect 117314 136620 117320 136632
rect 117372 136620 117378 136672
rect 24210 135260 24216 135312
rect 24268 135300 24274 135312
rect 117314 135300 117320 135312
rect 24268 135272 117320 135300
rect 24268 135260 24274 135272
rect 117314 135260 117320 135272
rect 117372 135260 117378 135312
rect 190638 134444 190644 134496
rect 190696 134484 190702 134496
rect 191006 134484 191012 134496
rect 190696 134456 191012 134484
rect 190696 134444 190702 134456
rect 191006 134444 191012 134456
rect 191064 134444 191070 134496
rect 21358 133900 21364 133952
rect 21416 133940 21422 133952
rect 117314 133940 117320 133952
rect 21416 133912 117320 133940
rect 21416 133900 21422 133912
rect 117314 133900 117320 133912
rect 117372 133900 117378 133952
rect 29638 133832 29644 133884
rect 29696 133872 29702 133884
rect 117406 133872 117412 133884
rect 29696 133844 117412 133872
rect 29696 133832 29702 133844
rect 117406 133832 117412 133844
rect 117464 133832 117470 133884
rect 24118 132404 24124 132456
rect 24176 132444 24182 132456
rect 117314 132444 117320 132456
rect 24176 132416 117320 132444
rect 24176 132404 24182 132416
rect 117314 132404 117320 132416
rect 117372 132404 117378 132456
rect 22922 131044 22928 131096
rect 22980 131084 22986 131096
rect 117314 131084 117320 131096
rect 22980 131056 117320 131084
rect 22980 131044 22986 131056
rect 117314 131044 117320 131056
rect 117372 131044 117378 131096
rect 4890 129684 4896 129736
rect 4948 129724 4954 129736
rect 117314 129724 117320 129736
rect 4948 129696 117320 129724
rect 4948 129684 4954 129696
rect 117314 129684 117320 129696
rect 117372 129684 117378 129736
rect 22830 128256 22836 128308
rect 22888 128296 22894 128308
rect 117314 128296 117320 128308
rect 22888 128268 117320 128296
rect 22888 128256 22894 128268
rect 117314 128256 117320 128268
rect 117372 128256 117378 128308
rect 22738 126896 22744 126948
rect 22796 126936 22802 126948
rect 117314 126936 117320 126948
rect 22796 126908 117320 126936
rect 22796 126896 22802 126908
rect 117314 126896 117320 126908
rect 117372 126896 117378 126948
rect 19978 124108 19984 124160
rect 20036 124148 20042 124160
rect 117314 124148 117320 124160
rect 20036 124120 117320 124148
rect 20036 124108 20042 124120
rect 117314 124108 117320 124120
rect 117372 124108 117378 124160
rect 15838 122748 15844 122800
rect 15896 122788 15902 122800
rect 117314 122788 117320 122800
rect 15896 122760 117320 122788
rect 15896 122748 15902 122760
rect 117314 122748 117320 122760
rect 117372 122748 117378 122800
rect 7558 121388 7564 121440
rect 7616 121428 7622 121440
rect 117314 121428 117320 121440
rect 7616 121400 117320 121428
rect 7616 121388 7622 121400
rect 117314 121388 117320 121400
rect 117372 121388 117378 121440
rect 4798 120028 4804 120080
rect 4856 120068 4862 120080
rect 117314 120068 117320 120080
rect 4856 120040 117320 120068
rect 4856 120028 4862 120040
rect 117314 120028 117320 120040
rect 117372 120028 117378 120080
rect 6178 118600 6184 118652
rect 6236 118640 6242 118652
rect 117314 118640 117320 118652
rect 6236 118612 117320 118640
rect 6236 118600 6242 118612
rect 117314 118600 117320 118612
rect 117372 118600 117378 118652
rect 189258 118600 189264 118652
rect 189316 118640 189322 118652
rect 189442 118640 189448 118652
rect 189316 118612 189448 118640
rect 189316 118600 189322 118612
rect 189442 118600 189448 118612
rect 189500 118600 189506 118652
rect 40034 117240 40040 117292
rect 40092 117280 40098 117292
rect 117314 117280 117320 117292
rect 40092 117252 117320 117280
rect 40092 117240 40098 117252
rect 117314 117240 117320 117252
rect 117372 117240 117378 117292
rect 189166 117240 189172 117292
rect 189224 117280 189230 117292
rect 189442 117280 189448 117292
rect 189224 117252 189448 117280
rect 189224 117240 189230 117252
rect 189442 117240 189448 117252
rect 189500 117240 189506 117292
rect 106918 115880 106924 115932
rect 106976 115920 106982 115932
rect 117314 115920 117320 115932
rect 106976 115892 117320 115920
rect 106976 115880 106982 115892
rect 117314 115880 117320 115892
rect 117372 115880 117378 115932
rect 189074 114452 189080 114504
rect 189132 114492 189138 114504
rect 189442 114492 189448 114504
rect 189132 114464 189448 114492
rect 189132 114452 189138 114464
rect 189442 114452 189448 114464
rect 189500 114452 189506 114504
rect 193122 113092 193128 113144
rect 193180 113132 193186 113144
rect 207658 113132 207664 113144
rect 193180 113104 207664 113132
rect 193180 113092 193186 113104
rect 207658 113092 207664 113104
rect 207716 113092 207722 113144
rect 189718 111800 189724 111852
rect 189776 111840 189782 111852
rect 580074 111840 580080 111852
rect 189776 111812 580080 111840
rect 189776 111800 189782 111812
rect 580074 111800 580080 111812
rect 580132 111800 580138 111852
rect 3326 111732 3332 111784
rect 3384 111772 3390 111784
rect 21358 111772 21364 111784
rect 3384 111744 21364 111772
rect 3384 111732 3390 111744
rect 21358 111732 21364 111744
rect 21416 111732 21422 111784
rect 193122 111732 193128 111784
rect 193180 111772 193186 111784
rect 206278 111772 206284 111784
rect 193180 111744 206284 111772
rect 193180 111732 193186 111744
rect 206278 111732 206284 111744
rect 206336 111732 206342 111784
rect 193030 110372 193036 110424
rect 193088 110412 193094 110424
rect 203518 110412 203524 110424
rect 193088 110384 203524 110412
rect 193088 110372 193094 110384
rect 203518 110372 203524 110384
rect 203576 110372 203582 110424
rect 193030 108944 193036 108996
rect 193088 108984 193094 108996
rect 200758 108984 200764 108996
rect 193088 108956 200764 108984
rect 193088 108944 193094 108956
rect 200758 108944 200764 108956
rect 200816 108944 200822 108996
rect 193122 106156 193128 106208
rect 193180 106196 193186 106208
rect 199378 106196 199384 106208
rect 193180 106168 199384 106196
rect 193180 106156 193186 106168
rect 199378 106156 199384 106168
rect 199436 106156 199442 106208
rect 193122 104660 193128 104712
rect 193180 104700 193186 104712
rect 197998 104700 198004 104712
rect 193180 104672 198004 104700
rect 193180 104660 193186 104672
rect 197998 104660 198004 104672
rect 198056 104660 198062 104712
rect 193122 103164 193128 103216
rect 193180 103204 193186 103216
rect 196618 103204 196624 103216
rect 193180 103176 196624 103204
rect 193180 103164 193186 103176
rect 196618 103164 196624 103176
rect 196676 103164 196682 103216
rect 192202 101736 192208 101788
rect 192260 101776 192266 101788
rect 193858 101776 193864 101788
rect 192260 101748 193864 101776
rect 192260 101736 192266 101748
rect 193858 101736 193864 101748
rect 193916 101736 193922 101788
rect 192202 100376 192208 100428
rect 192260 100416 192266 100428
rect 193950 100416 193956 100428
rect 192260 100388 193956 100416
rect 192260 100376 192266 100388
rect 193950 100376 193956 100388
rect 194008 100376 194014 100428
rect 192202 98812 192208 98864
rect 192260 98852 192266 98864
rect 194042 98852 194048 98864
rect 192260 98824 194048 98852
rect 192260 98812 192266 98824
rect 194042 98812 194048 98824
rect 194100 98812 194106 98864
rect 193122 97928 193128 97980
rect 193180 97968 193186 97980
rect 580442 97968 580448 97980
rect 193180 97940 580448 97968
rect 193180 97928 193186 97940
rect 580442 97928 580448 97940
rect 580500 97928 580506 97980
rect 193122 95140 193128 95192
rect 193180 95180 193186 95192
rect 366358 95180 366364 95192
rect 193180 95152 366364 95180
rect 193180 95140 193186 95152
rect 366358 95140 366364 95152
rect 366416 95140 366422 95192
rect 193122 93780 193128 93832
rect 193180 93820 193186 93832
rect 362218 93820 362224 93832
rect 193180 93792 362224 93820
rect 193180 93780 193186 93792
rect 362218 93780 362224 93792
rect 362276 93780 362282 93832
rect 193122 92420 193128 92472
rect 193180 92460 193186 92472
rect 531958 92460 531964 92472
rect 193180 92432 531964 92460
rect 193180 92420 193186 92432
rect 531958 92420 531964 92432
rect 532016 92420 532022 92472
rect 193122 89632 193128 89684
rect 193180 89672 193186 89684
rect 532050 89672 532056 89684
rect 193180 89644 532056 89672
rect 193180 89632 193186 89644
rect 532050 89632 532056 89644
rect 532108 89632 532114 89684
rect 193122 88272 193128 88324
rect 193180 88312 193186 88324
rect 358078 88312 358084 88324
rect 193180 88284 358084 88312
rect 193180 88272 193186 88284
rect 358078 88272 358084 88284
rect 358136 88272 358142 88324
rect 193122 86912 193128 86964
rect 193180 86952 193186 86964
rect 580718 86952 580724 86964
rect 193180 86924 580724 86952
rect 193180 86912 193186 86924
rect 580718 86912 580724 86924
rect 580776 86912 580782 86964
rect 193122 85484 193128 85536
rect 193180 85524 193186 85536
rect 580902 85524 580908 85536
rect 193180 85496 580908 85524
rect 193180 85484 193186 85496
rect 580902 85484 580908 85496
rect 580960 85484 580966 85536
rect 192846 81404 192852 81456
rect 192904 81444 192910 81456
rect 347038 81444 347044 81456
rect 192904 81416 347044 81444
rect 192904 81404 192910 81416
rect 347038 81404 347044 81416
rect 347096 81404 347102 81456
rect 118602 80928 118608 80980
rect 118660 80968 118666 80980
rect 579982 80968 579988 80980
rect 118660 80940 579988 80968
rect 118660 80928 118666 80940
rect 579982 80928 579988 80940
rect 580040 80928 580046 80980
rect 4982 80792 4988 80844
rect 5040 80832 5046 80844
rect 5040 80804 172514 80832
rect 5040 80792 5046 80804
rect 3694 80656 3700 80708
rect 3752 80696 3758 80708
rect 172486 80696 172514 80804
rect 176718 80804 179736 80832
rect 176718 80764 176746 80804
rect 176626 80736 176746 80764
rect 176626 80696 176654 80736
rect 3752 80668 157334 80696
rect 172486 80668 176654 80696
rect 179708 80696 179736 80804
rect 179782 80696 179788 80708
rect 179708 80668 179788 80696
rect 3752 80656 3758 80668
rect 157306 80628 157334 80668
rect 179782 80656 179788 80668
rect 179840 80656 179846 80708
rect 179506 80628 179512 80640
rect 157306 80600 179512 80628
rect 179506 80588 179512 80600
rect 179564 80588 179570 80640
rect 180242 80560 180248 80572
rect 137986 80532 147674 80560
rect 127802 80384 127808 80436
rect 127860 80424 127866 80436
rect 137986 80424 138014 80532
rect 127860 80396 138014 80424
rect 127860 80384 127866 80396
rect 129366 80248 129372 80300
rect 129424 80288 129430 80300
rect 129424 80260 133966 80288
rect 129424 80248 129430 80260
rect 129274 80112 129280 80164
rect 129332 80152 129338 80164
rect 129332 80124 132126 80152
rect 129332 80112 129338 80124
rect 130470 80016 130476 80028
rect 125566 79988 130476 80016
rect 116578 79772 116584 79824
rect 116636 79812 116642 79824
rect 125566 79812 125594 79988
rect 130470 79976 130476 79988
rect 130528 79976 130534 80028
rect 132098 79960 132126 80124
rect 133938 79960 133966 80260
rect 147646 80220 147674 80532
rect 164206 80532 180248 80560
rect 147646 80192 157886 80220
rect 136238 79988 136634 80016
rect 136238 79960 136266 79988
rect 130700 79908 130706 79960
rect 130758 79908 130764 79960
rect 130792 79908 130798 79960
rect 130850 79908 130856 79960
rect 131344 79948 131350 79960
rect 131178 79920 131350 79948
rect 130718 79880 130746 79908
rect 130672 79852 130746 79880
rect 130672 79824 130700 79852
rect 130810 79824 130838 79908
rect 116636 79784 125594 79812
rect 116636 79772 116642 79784
rect 130654 79772 130660 79824
rect 130712 79772 130718 79824
rect 130746 79772 130752 79824
rect 130804 79784 130838 79824
rect 131178 79812 131206 79920
rect 131344 79908 131350 79920
rect 131402 79908 131408 79960
rect 131804 79908 131810 79960
rect 131862 79908 131868 79960
rect 132080 79908 132086 79960
rect 132138 79908 132144 79960
rect 132172 79908 132178 79960
rect 132230 79908 132236 79960
rect 132264 79908 132270 79960
rect 132322 79908 132328 79960
rect 132356 79908 132362 79960
rect 132414 79908 132420 79960
rect 132632 79908 132638 79960
rect 132690 79908 132696 79960
rect 133368 79908 133374 79960
rect 133426 79908 133432 79960
rect 133828 79948 133834 79960
rect 133478 79920 133834 79948
rect 131436 79880 131442 79892
rect 131040 79784 131206 79812
rect 131316 79852 131442 79880
rect 130804 79772 130810 79784
rect 130562 79704 130568 79756
rect 130620 79744 130626 79756
rect 131040 79744 131068 79784
rect 130620 79716 131068 79744
rect 130620 79704 130626 79716
rect 131316 79688 131344 79852
rect 131436 79840 131442 79852
rect 131494 79840 131500 79892
rect 131822 79756 131850 79908
rect 132190 79812 132218 79908
rect 132144 79784 132218 79812
rect 132144 79756 132172 79784
rect 132282 79756 132310 79908
rect 131758 79704 131764 79756
rect 131816 79716 131850 79756
rect 131816 79704 131822 79716
rect 132126 79704 132132 79756
rect 132184 79704 132190 79756
rect 132218 79704 132224 79756
rect 132276 79716 132310 79756
rect 132276 79704 132282 79716
rect 132374 79688 132402 79908
rect 131298 79636 131304 79688
rect 131356 79636 131362 79688
rect 132310 79636 132316 79688
rect 132368 79648 132402 79688
rect 132368 79636 132374 79648
rect 132494 79636 132500 79688
rect 132552 79676 132558 79688
rect 132650 79676 132678 79908
rect 133000 79840 133006 79892
rect 133058 79840 133064 79892
rect 132552 79648 132678 79676
rect 132552 79636 132558 79648
rect 132770 79636 132776 79688
rect 132828 79676 132834 79688
rect 133018 79676 133046 79840
rect 132828 79648 133046 79676
rect 132828 79636 132834 79648
rect 133230 79636 133236 79688
rect 133288 79676 133294 79688
rect 133386 79676 133414 79908
rect 133288 79648 133414 79676
rect 133478 79688 133506 79920
rect 133828 79908 133834 79920
rect 133886 79908 133892 79960
rect 133920 79908 133926 79960
rect 133978 79908 133984 79960
rect 135116 79908 135122 79960
rect 135174 79908 135180 79960
rect 135208 79908 135214 79960
rect 135266 79908 135272 79960
rect 135392 79908 135398 79960
rect 135450 79908 135456 79960
rect 135576 79908 135582 79960
rect 135634 79908 135640 79960
rect 136220 79908 136226 79960
rect 136278 79908 136284 79960
rect 136496 79908 136502 79960
rect 136554 79908 136560 79960
rect 133552 79840 133558 79892
rect 133610 79880 133616 79892
rect 133610 79852 134012 79880
rect 133610 79840 133616 79852
rect 133984 79824 134012 79852
rect 134472 79840 134478 79892
rect 134530 79840 134536 79892
rect 134932 79840 134938 79892
rect 134990 79840 134996 79892
rect 133966 79772 133972 79824
rect 134024 79772 134030 79824
rect 133478 79648 133512 79688
rect 133288 79636 133294 79648
rect 133506 79636 133512 79648
rect 133564 79636 133570 79688
rect 134490 79676 134518 79840
rect 134564 79772 134570 79824
rect 134622 79772 134628 79824
rect 134656 79772 134662 79824
rect 134714 79772 134720 79824
rect 134444 79648 134518 79676
rect 116670 79500 116676 79552
rect 116728 79540 116734 79552
rect 127802 79540 127808 79552
rect 116728 79512 127808 79540
rect 116728 79500 116734 79512
rect 127802 79500 127808 79512
rect 127860 79500 127866 79552
rect 79318 79432 79324 79484
rect 79376 79472 79382 79484
rect 131666 79472 131672 79484
rect 79376 79444 131672 79472
rect 79376 79432 79382 79444
rect 131666 79432 131672 79444
rect 131724 79432 131730 79484
rect 4062 79364 4068 79416
rect 4120 79404 4126 79416
rect 4120 79376 125594 79404
rect 4120 79364 4126 79376
rect 3878 79296 3884 79348
rect 3936 79336 3942 79348
rect 125566 79336 125594 79376
rect 134058 79364 134064 79416
rect 134116 79404 134122 79416
rect 134444 79404 134472 79648
rect 134582 79552 134610 79772
rect 134518 79500 134524 79552
rect 134576 79512 134610 79552
rect 134576 79500 134582 79512
rect 134674 79484 134702 79772
rect 134674 79444 134708 79484
rect 134702 79432 134708 79444
rect 134760 79432 134766 79484
rect 134116 79376 134472 79404
rect 134116 79364 134122 79376
rect 134610 79364 134616 79416
rect 134668 79404 134674 79416
rect 134950 79404 134978 79840
rect 135134 79688 135162 79908
rect 135070 79636 135076 79688
rect 135128 79648 135162 79688
rect 135128 79636 135134 79648
rect 135226 79620 135254 79908
rect 135410 79744 135438 79908
rect 135364 79716 135438 79744
rect 135364 79688 135392 79716
rect 135346 79636 135352 79688
rect 135404 79636 135410 79688
rect 135162 79568 135168 79620
rect 135220 79580 135254 79620
rect 135594 79620 135622 79908
rect 135760 79880 135766 79892
rect 135732 79840 135766 79880
rect 135818 79840 135824 79892
rect 135852 79840 135858 79892
rect 135910 79840 135916 79892
rect 135944 79840 135950 79892
rect 136002 79840 136008 79892
rect 136036 79840 136042 79892
rect 136094 79840 136100 79892
rect 135732 79756 135760 79840
rect 135870 79756 135898 79840
rect 135714 79704 135720 79756
rect 135772 79704 135778 79756
rect 135806 79704 135812 79756
rect 135864 79716 135898 79756
rect 135864 79704 135870 79716
rect 135594 79580 135628 79620
rect 135220 79568 135226 79580
rect 135622 79568 135628 79580
rect 135680 79568 135686 79620
rect 135962 79552 135990 79840
rect 136054 79620 136082 79840
rect 136514 79824 136542 79908
rect 136312 79772 136318 79824
rect 136370 79772 136376 79824
rect 136450 79772 136456 79824
rect 136508 79784 136542 79824
rect 136508 79772 136514 79784
rect 136054 79580 136088 79620
rect 136082 79568 136088 79580
rect 136140 79568 136146 79620
rect 135962 79512 135996 79552
rect 135990 79500 135996 79512
rect 136048 79500 136054 79552
rect 136330 79540 136358 79772
rect 136606 79608 136634 79988
rect 137158 79988 137554 80016
rect 136864 79948 136870 79960
rect 136100 79512 136358 79540
rect 136422 79580 136634 79608
rect 136698 79920 136870 79948
rect 135530 79432 135536 79484
rect 135588 79472 135594 79484
rect 136100 79472 136128 79512
rect 135588 79444 136128 79472
rect 135588 79432 135594 79444
rect 136266 79432 136272 79484
rect 136324 79472 136330 79484
rect 136422 79472 136450 79580
rect 136698 79552 136726 79920
rect 136864 79908 136870 79920
rect 136922 79908 136928 79960
rect 137048 79908 137054 79960
rect 137106 79908 137112 79960
rect 137066 79552 137094 79908
rect 137158 79688 137186 79988
rect 137526 79960 137554 79988
rect 139826 79988 140222 80016
rect 137232 79908 137238 79960
rect 137290 79948 137296 79960
rect 137290 79908 137324 79948
rect 137508 79908 137514 79960
rect 137566 79908 137572 79960
rect 137968 79908 137974 79960
rect 138026 79908 138032 79960
rect 138060 79908 138066 79960
rect 138118 79908 138124 79960
rect 138152 79908 138158 79960
rect 138210 79908 138216 79960
rect 138428 79908 138434 79960
rect 138486 79908 138492 79960
rect 138520 79908 138526 79960
rect 138578 79908 138584 79960
rect 138888 79948 138894 79960
rect 138630 79920 138894 79948
rect 137158 79648 137192 79688
rect 137186 79636 137192 79648
rect 137244 79636 137250 79688
rect 136634 79500 136640 79552
rect 136692 79512 136726 79552
rect 136692 79500 136698 79512
rect 137002 79500 137008 79552
rect 137060 79512 137094 79552
rect 137060 79500 137066 79512
rect 136324 79444 136450 79472
rect 137296 79472 137324 79908
rect 137416 79840 137422 79892
rect 137474 79840 137480 79892
rect 137434 79552 137462 79840
rect 137986 79812 138014 79908
rect 137848 79784 138014 79812
rect 137848 79608 137876 79784
rect 138078 79744 138106 79908
rect 137940 79716 138106 79744
rect 137940 79688 137968 79716
rect 138170 79688 138198 79908
rect 138446 79824 138474 79908
rect 138428 79772 138434 79824
rect 138486 79772 138492 79824
rect 137922 79636 137928 79688
rect 137980 79636 137986 79688
rect 138106 79636 138112 79688
rect 138164 79648 138198 79688
rect 138538 79676 138566 79908
rect 138308 79648 138566 79676
rect 138164 79636 138170 79648
rect 138014 79608 138020 79620
rect 137848 79580 138020 79608
rect 138014 79568 138020 79580
rect 138072 79568 138078 79620
rect 137370 79500 137376 79552
rect 137428 79512 137462 79552
rect 137428 79500 137434 79512
rect 137646 79472 137652 79484
rect 137296 79444 137652 79472
rect 136324 79432 136330 79444
rect 137646 79432 137652 79444
rect 137704 79432 137710 79484
rect 138198 79432 138204 79484
rect 138256 79472 138262 79484
rect 138308 79472 138336 79648
rect 138474 79568 138480 79620
rect 138532 79608 138538 79620
rect 138630 79608 138658 79920
rect 138888 79908 138894 79920
rect 138946 79908 138952 79960
rect 138980 79908 138986 79960
rect 139038 79908 139044 79960
rect 139256 79908 139262 79960
rect 139314 79908 139320 79960
rect 139348 79908 139354 79960
rect 139406 79908 139412 79960
rect 138704 79840 138710 79892
rect 138762 79840 138768 79892
rect 138532 79580 138658 79608
rect 138532 79568 138538 79580
rect 138722 79552 138750 79840
rect 138998 79688 139026 79908
rect 139274 79744 139302 79908
rect 139228 79716 139302 79744
rect 139228 79688 139256 79716
rect 139366 79688 139394 79908
rect 139532 79840 139538 79892
rect 139590 79840 139596 79892
rect 139550 79688 139578 79840
rect 139624 79772 139630 79824
rect 139682 79772 139688 79824
rect 138934 79636 138940 79688
rect 138992 79648 139026 79688
rect 138992 79636 138998 79648
rect 139210 79636 139216 79688
rect 139268 79636 139274 79688
rect 139302 79636 139308 79688
rect 139360 79648 139394 79688
rect 139360 79636 139366 79648
rect 139486 79636 139492 79688
rect 139544 79648 139578 79688
rect 139544 79636 139550 79648
rect 138658 79500 138664 79552
rect 138716 79512 138750 79552
rect 138716 79500 138722 79512
rect 139486 79500 139492 79552
rect 139544 79540 139550 79552
rect 139642 79540 139670 79772
rect 139826 79608 139854 79988
rect 140194 79960 140222 79988
rect 150866 79988 151170 80016
rect 150866 79960 150894 79988
rect 139992 79908 139998 79960
rect 140050 79908 140056 79960
rect 140084 79908 140090 79960
rect 140142 79908 140148 79960
rect 140176 79908 140182 79960
rect 140234 79908 140240 79960
rect 141832 79948 141838 79960
rect 141804 79908 141838 79948
rect 141890 79908 141896 79960
rect 142384 79908 142390 79960
rect 142442 79908 142448 79960
rect 142844 79908 142850 79960
rect 142902 79908 142908 79960
rect 143212 79908 143218 79960
rect 143270 79908 143276 79960
rect 144316 79908 144322 79960
rect 144374 79948 144380 79960
rect 144374 79920 144592 79948
rect 144374 79908 144380 79920
rect 140010 79688 140038 79908
rect 139946 79636 139952 79688
rect 140004 79648 140038 79688
rect 140004 79636 140010 79648
rect 139544 79512 139670 79540
rect 139780 79580 139854 79608
rect 139544 79500 139550 79512
rect 138256 79444 138336 79472
rect 138256 79432 138262 79444
rect 139780 79416 139808 79580
rect 134668 79376 134978 79404
rect 134668 79364 134674 79376
rect 136910 79364 136916 79416
rect 136968 79404 136974 79416
rect 137462 79404 137468 79416
rect 136968 79376 137468 79404
rect 136968 79364 136974 79376
rect 137462 79364 137468 79376
rect 137520 79364 137526 79416
rect 138842 79364 138848 79416
rect 138900 79404 138906 79416
rect 139118 79404 139124 79416
rect 138900 79376 139124 79404
rect 138900 79364 138906 79376
rect 139118 79364 139124 79376
rect 139176 79364 139182 79416
rect 139762 79364 139768 79416
rect 139820 79364 139826 79416
rect 139946 79364 139952 79416
rect 140004 79404 140010 79416
rect 140102 79404 140130 79908
rect 140452 79840 140458 79892
rect 140510 79840 140516 79892
rect 140728 79840 140734 79892
rect 140786 79840 140792 79892
rect 140912 79840 140918 79892
rect 140970 79840 140976 79892
rect 141004 79840 141010 79892
rect 141062 79840 141068 79892
rect 141464 79840 141470 79892
rect 141522 79840 141528 79892
rect 141648 79880 141654 79892
rect 141620 79840 141654 79880
rect 141706 79840 141712 79892
rect 140360 79812 140366 79824
rect 140240 79784 140366 79812
rect 140240 79756 140268 79784
rect 140360 79772 140366 79784
rect 140418 79772 140424 79824
rect 140222 79704 140228 79756
rect 140280 79704 140286 79756
rect 140470 79688 140498 79840
rect 140406 79636 140412 79688
rect 140464 79648 140498 79688
rect 140464 79636 140470 79648
rect 140746 79620 140774 79840
rect 140746 79580 140780 79620
rect 140774 79568 140780 79580
rect 140832 79568 140838 79620
rect 140930 79552 140958 79840
rect 141022 79620 141050 79840
rect 141096 79772 141102 79824
rect 141154 79772 141160 79824
rect 141280 79772 141286 79824
rect 141338 79812 141344 79824
rect 141338 79784 141418 79812
rect 141338 79772 141344 79784
rect 141114 79676 141142 79772
rect 141390 79756 141418 79784
rect 141372 79704 141378 79756
rect 141430 79704 141436 79756
rect 141114 79648 141188 79676
rect 141022 79580 141056 79620
rect 141050 79568 141056 79580
rect 141108 79568 141114 79620
rect 140930 79512 140964 79552
rect 140958 79500 140964 79512
rect 141016 79500 141022 79552
rect 140590 79432 140596 79484
rect 140648 79472 140654 79484
rect 141160 79472 141188 79648
rect 140648 79444 141188 79472
rect 140648 79432 140654 79444
rect 140004 79376 140130 79404
rect 140004 79364 140010 79376
rect 141142 79364 141148 79416
rect 141200 79404 141206 79416
rect 141482 79404 141510 79840
rect 141620 79620 141648 79840
rect 141804 79756 141832 79908
rect 142402 79880 142430 79908
rect 141896 79852 142430 79880
rect 141896 79756 141924 79852
rect 141786 79704 141792 79756
rect 141844 79704 141850 79756
rect 141878 79704 141884 79756
rect 141936 79704 141942 79756
rect 142246 79636 142252 79688
rect 142304 79676 142310 79688
rect 142862 79676 142890 79908
rect 142936 79840 142942 79892
rect 142994 79840 143000 79892
rect 142954 79744 142982 79840
rect 142954 79716 143120 79744
rect 143092 79688 143120 79716
rect 143230 79688 143258 79908
rect 143856 79840 143862 79892
rect 143914 79840 143920 79892
rect 144224 79840 144230 79892
rect 144282 79840 144288 79892
rect 142304 79648 142890 79676
rect 142304 79636 142310 79648
rect 143074 79636 143080 79688
rect 143132 79636 143138 79688
rect 143166 79636 143172 79688
rect 143224 79648 143258 79688
rect 143874 79676 143902 79840
rect 144242 79688 144270 79840
rect 143994 79676 144000 79688
rect 143874 79648 144000 79676
rect 143224 79636 143230 79648
rect 143994 79636 144000 79648
rect 144052 79636 144058 79688
rect 144242 79648 144276 79688
rect 144270 79636 144276 79648
rect 144328 79636 144334 79688
rect 144564 79620 144592 79920
rect 144684 79908 144690 79960
rect 144742 79908 144748 79960
rect 144868 79908 144874 79960
rect 144926 79908 144932 79960
rect 145788 79948 145794 79960
rect 145116 79920 145794 79948
rect 144702 79688 144730 79908
rect 144638 79636 144644 79688
rect 144696 79648 144730 79688
rect 144696 79636 144702 79648
rect 144886 79620 144914 79908
rect 145116 79620 145144 79920
rect 145788 79908 145794 79920
rect 145846 79908 145852 79960
rect 145972 79948 145978 79960
rect 145944 79908 145978 79948
rect 146030 79908 146036 79960
rect 146708 79948 146714 79960
rect 146312 79920 146714 79948
rect 145328 79840 145334 79892
rect 145386 79880 145392 79892
rect 145386 79852 145788 79880
rect 145386 79840 145392 79852
rect 145512 79772 145518 79824
rect 145570 79812 145576 79824
rect 145570 79784 145696 79812
rect 145570 79772 145576 79784
rect 145668 79688 145696 79784
rect 145760 79688 145788 79852
rect 145944 79688 145972 79908
rect 146156 79880 146162 79892
rect 146036 79852 146162 79880
rect 145650 79636 145656 79688
rect 145708 79636 145714 79688
rect 145742 79636 145748 79688
rect 145800 79636 145806 79688
rect 145926 79636 145932 79688
rect 145984 79636 145990 79688
rect 141602 79568 141608 79620
rect 141660 79568 141666 79620
rect 144546 79568 144552 79620
rect 144604 79568 144610 79620
rect 144822 79568 144828 79620
rect 144880 79580 144914 79620
rect 144880 79568 144886 79580
rect 145006 79568 145012 79620
rect 145064 79568 145070 79620
rect 145098 79568 145104 79620
rect 145156 79568 145162 79620
rect 145466 79568 145472 79620
rect 145524 79608 145530 79620
rect 146036 79608 146064 79852
rect 146156 79840 146162 79852
rect 146214 79840 146220 79892
rect 146312 79688 146340 79920
rect 146708 79908 146714 79920
rect 146766 79908 146772 79960
rect 147352 79908 147358 79960
rect 147410 79908 147416 79960
rect 148272 79908 148278 79960
rect 148330 79908 148336 79960
rect 148364 79908 148370 79960
rect 148422 79908 148428 79960
rect 148456 79908 148462 79960
rect 148514 79908 148520 79960
rect 148548 79908 148554 79960
rect 148606 79908 148612 79960
rect 148916 79948 148922 79960
rect 148888 79908 148922 79948
rect 148974 79908 148980 79960
rect 149192 79908 149198 79960
rect 149250 79908 149256 79960
rect 150848 79908 150854 79960
rect 150906 79908 150912 79960
rect 151032 79908 151038 79960
rect 151090 79908 151096 79960
rect 146524 79840 146530 79892
rect 146582 79880 146588 79892
rect 146800 79880 146806 79892
rect 146582 79840 146616 79880
rect 146588 79688 146616 79840
rect 146680 79852 146806 79880
rect 146680 79688 146708 79852
rect 146800 79840 146806 79852
rect 146858 79840 146864 79892
rect 146984 79840 146990 79892
rect 147042 79840 147048 79892
rect 147002 79744 147030 79840
rect 147370 79824 147398 79908
rect 148290 79824 148318 79908
rect 147306 79772 147312 79824
rect 147364 79784 147398 79824
rect 147364 79772 147370 79784
rect 147536 79772 147542 79824
rect 147594 79772 147600 79824
rect 147720 79772 147726 79824
rect 147778 79772 147784 79824
rect 148088 79772 148094 79824
rect 148146 79772 148152 79824
rect 148226 79772 148232 79824
rect 148284 79784 148318 79824
rect 148284 79772 148290 79784
rect 146772 79716 147030 79744
rect 146294 79636 146300 79688
rect 146352 79636 146358 79688
rect 146570 79636 146576 79688
rect 146628 79636 146634 79688
rect 146662 79636 146668 79688
rect 146720 79636 146726 79688
rect 145524 79580 146064 79608
rect 145524 79568 145530 79580
rect 146386 79568 146392 79620
rect 146444 79608 146450 79620
rect 146772 79608 146800 79716
rect 147554 79676 147582 79772
rect 146956 79648 147582 79676
rect 146956 79620 146984 79648
rect 146444 79580 146800 79608
rect 146444 79568 146450 79580
rect 146938 79568 146944 79620
rect 146996 79568 147002 79620
rect 147738 79608 147766 79772
rect 147738 79580 147996 79608
rect 145024 79540 145052 79568
rect 147968 79552 147996 79580
rect 147858 79540 147864 79552
rect 145024 79512 147864 79540
rect 147858 79500 147864 79512
rect 147916 79500 147922 79552
rect 147950 79500 147956 79552
rect 148008 79500 148014 79552
rect 148106 79540 148134 79772
rect 148382 79756 148410 79908
rect 148474 79812 148502 79908
rect 148566 79880 148594 79908
rect 148566 79852 148640 79880
rect 148474 79784 148548 79812
rect 148520 79756 148548 79784
rect 148382 79716 148416 79756
rect 148410 79704 148416 79716
rect 148468 79704 148474 79756
rect 148502 79704 148508 79756
rect 148560 79704 148566 79756
rect 148612 79688 148640 79852
rect 148732 79840 148738 79892
rect 148790 79840 148796 79892
rect 148594 79636 148600 79688
rect 148652 79636 148658 79688
rect 148750 79620 148778 79840
rect 148888 79688 148916 79908
rect 149210 79756 149238 79908
rect 149376 79880 149382 79892
rect 149348 79840 149382 79880
rect 149434 79840 149440 79892
rect 149468 79840 149474 79892
rect 149526 79840 149532 79892
rect 149560 79840 149566 79892
rect 149618 79840 149624 79892
rect 151050 79880 151078 79908
rect 151004 79852 151078 79880
rect 149348 79756 149376 79840
rect 149210 79716 149244 79756
rect 149238 79704 149244 79716
rect 149296 79704 149302 79756
rect 149330 79704 149336 79756
rect 149388 79704 149394 79756
rect 149486 79744 149514 79840
rect 149440 79716 149514 79744
rect 148870 79636 148876 79688
rect 148928 79636 148934 79688
rect 149440 79620 149468 79716
rect 149578 79688 149606 79840
rect 150296 79772 150302 79824
rect 150354 79772 150360 79824
rect 150480 79772 150486 79824
rect 150538 79772 150544 79824
rect 150664 79772 150670 79824
rect 150722 79772 150728 79824
rect 149514 79636 149520 79688
rect 149572 79648 149606 79688
rect 149572 79636 149578 79648
rect 150158 79636 150164 79688
rect 150216 79676 150222 79688
rect 150314 79676 150342 79772
rect 150216 79648 150342 79676
rect 150216 79636 150222 79648
rect 148686 79568 148692 79620
rect 148744 79580 148778 79620
rect 148744 79568 148750 79580
rect 149422 79568 149428 79620
rect 149480 79568 149486 79620
rect 150498 79608 150526 79772
rect 150682 79688 150710 79772
rect 151004 79756 151032 79852
rect 151142 79824 151170 79988
rect 153902 79988 154206 80016
rect 153902 79960 153930 79988
rect 151860 79908 151866 79960
rect 151918 79908 151924 79960
rect 152412 79908 152418 79960
rect 152470 79908 152476 79960
rect 152872 79908 152878 79960
rect 152930 79908 152936 79960
rect 152964 79908 152970 79960
rect 153022 79948 153028 79960
rect 153022 79920 153148 79948
rect 153022 79908 153028 79920
rect 151078 79772 151084 79824
rect 151136 79784 151170 79824
rect 151136 79772 151142 79784
rect 150986 79704 150992 79756
rect 151044 79704 151050 79756
rect 150682 79648 150716 79688
rect 150710 79636 150716 79648
rect 150768 79636 150774 79688
rect 150618 79608 150624 79620
rect 150498 79580 150624 79608
rect 150618 79568 150624 79580
rect 150676 79568 150682 79620
rect 151538 79568 151544 79620
rect 151596 79608 151602 79620
rect 151878 79608 151906 79908
rect 152320 79840 152326 79892
rect 152378 79840 152384 79892
rect 152338 79688 152366 79840
rect 152430 79824 152458 79908
rect 152890 79880 152918 79908
rect 152890 79852 153056 79880
rect 153028 79824 153056 79852
rect 152412 79772 152418 79824
rect 152470 79772 152476 79824
rect 153010 79772 153016 79824
rect 153068 79772 153074 79824
rect 152338 79648 152372 79688
rect 152366 79636 152372 79648
rect 152424 79636 152430 79688
rect 151596 79580 151906 79608
rect 151596 79568 151602 79580
rect 148778 79540 148784 79552
rect 148106 79512 148784 79540
rect 148778 79500 148784 79512
rect 148836 79500 148842 79552
rect 153120 79540 153148 79920
rect 153424 79908 153430 79960
rect 153482 79908 153488 79960
rect 153608 79908 153614 79960
rect 153666 79948 153672 79960
rect 153666 79920 153746 79948
rect 153666 79908 153672 79920
rect 153286 79540 153292 79552
rect 153120 79512 153292 79540
rect 153286 79500 153292 79512
rect 153344 79500 153350 79552
rect 153442 79540 153470 79908
rect 153718 79688 153746 79920
rect 153884 79908 153890 79960
rect 153942 79908 153948 79960
rect 153976 79908 153982 79960
rect 154034 79908 154040 79960
rect 154068 79908 154074 79960
rect 154126 79908 154132 79960
rect 153792 79840 153798 79892
rect 153850 79880 153856 79892
rect 153850 79840 153884 79880
rect 153856 79756 153884 79840
rect 153838 79704 153844 79756
rect 153896 79704 153902 79756
rect 153718 79648 153752 79688
rect 153746 79636 153752 79648
rect 153804 79636 153810 79688
rect 153562 79568 153568 79620
rect 153620 79608 153626 79620
rect 153994 79608 154022 79908
rect 153620 79580 154022 79608
rect 153620 79568 153626 79580
rect 153654 79540 153660 79552
rect 153442 79512 153660 79540
rect 153654 79500 153660 79512
rect 153712 79500 153718 79552
rect 154086 79540 154114 79908
rect 154178 79824 154206 79988
rect 154344 79908 154350 79960
rect 154402 79948 154408 79960
rect 154804 79948 154810 79960
rect 154402 79920 154574 79948
rect 154402 79908 154408 79920
rect 154160 79772 154166 79824
rect 154218 79772 154224 79824
rect 154252 79772 154258 79824
rect 154310 79772 154316 79824
rect 154270 79688 154298 79772
rect 154206 79636 154212 79688
rect 154264 79648 154298 79688
rect 154546 79676 154574 79920
rect 154500 79648 154574 79676
rect 154638 79920 154810 79948
rect 154264 79636 154270 79648
rect 154500 79552 154528 79648
rect 154638 79620 154666 79920
rect 154804 79908 154810 79920
rect 154862 79908 154868 79960
rect 155264 79908 155270 79960
rect 155322 79908 155328 79960
rect 156092 79908 156098 79960
rect 156150 79908 156156 79960
rect 156368 79908 156374 79960
rect 156426 79908 156432 79960
rect 156828 79948 156834 79960
rect 156570 79920 156834 79948
rect 154712 79840 154718 79892
rect 154770 79840 154776 79892
rect 154730 79688 154758 79840
rect 155282 79688 155310 79908
rect 155448 79772 155454 79824
rect 155506 79772 155512 79824
rect 154730 79648 154764 79688
rect 154758 79636 154764 79648
rect 154816 79636 154822 79688
rect 155282 79648 155316 79688
rect 155310 79636 155316 79648
rect 155368 79636 155374 79688
rect 154574 79568 154580 79620
rect 154632 79580 154666 79620
rect 154632 79568 154638 79580
rect 154390 79540 154396 79552
rect 154086 79512 154396 79540
rect 154390 79500 154396 79512
rect 154448 79500 154454 79552
rect 154482 79500 154488 79552
rect 154540 79500 154546 79552
rect 154666 79500 154672 79552
rect 154724 79540 154730 79552
rect 155466 79540 155494 79772
rect 156110 79744 156138 79908
rect 156386 79824 156414 79908
rect 156460 79840 156466 79892
rect 156518 79840 156524 79892
rect 156368 79772 156374 79824
rect 156426 79772 156432 79824
rect 154724 79512 155494 79540
rect 155972 79716 156138 79744
rect 155972 79540 156000 79716
rect 156478 79676 156506 79840
rect 156064 79648 156506 79676
rect 156064 79620 156092 79648
rect 156046 79568 156052 79620
rect 156104 79568 156110 79620
rect 156138 79568 156144 79620
rect 156196 79608 156202 79620
rect 156570 79608 156598 79920
rect 156828 79908 156834 79920
rect 156886 79908 156892 79960
rect 156920 79908 156926 79960
rect 156978 79908 156984 79960
rect 157656 79908 157662 79960
rect 157714 79908 157720 79960
rect 156736 79840 156742 79892
rect 156794 79880 156800 79892
rect 156794 79840 156828 79880
rect 156800 79756 156828 79840
rect 156782 79704 156788 79756
rect 156840 79704 156846 79756
rect 156196 79580 156598 79608
rect 156196 79568 156202 79580
rect 156230 79540 156236 79552
rect 155972 79512 156236 79540
rect 154724 79500 154730 79512
rect 156230 79500 156236 79512
rect 156288 79500 156294 79552
rect 156690 79500 156696 79552
rect 156748 79540 156754 79552
rect 156938 79540 156966 79908
rect 157288 79840 157294 79892
rect 157346 79840 157352 79892
rect 157150 79568 157156 79620
rect 157208 79608 157214 79620
rect 157306 79608 157334 79840
rect 157208 79580 157334 79608
rect 157208 79568 157214 79580
rect 156748 79512 156966 79540
rect 157674 79540 157702 79908
rect 157858 79620 157886 80192
rect 164206 80152 164234 80532
rect 180242 80520 180248 80532
rect 180300 80520 180306 80572
rect 159698 80124 164234 80152
rect 167472 80464 182174 80492
rect 159698 79960 159726 80124
rect 160066 80056 166580 80084
rect 158024 79908 158030 79960
rect 158082 79908 158088 79960
rect 158484 79948 158490 79960
rect 158318 79920 158490 79948
rect 157794 79568 157800 79620
rect 157852 79580 157886 79620
rect 158042 79620 158070 79908
rect 158208 79840 158214 79892
rect 158266 79840 158272 79892
rect 158042 79580 158076 79620
rect 157852 79568 157858 79580
rect 158070 79568 158076 79580
rect 158128 79568 158134 79620
rect 158226 79608 158254 79840
rect 158318 79756 158346 79920
rect 158484 79908 158490 79920
rect 158542 79908 158548 79960
rect 158760 79908 158766 79960
rect 158818 79908 158824 79960
rect 158852 79908 158858 79960
rect 158910 79948 158916 79960
rect 158910 79920 159634 79948
rect 158910 79908 158916 79920
rect 158392 79840 158398 79892
rect 158450 79880 158456 79892
rect 158450 79852 158668 79880
rect 158450 79840 158456 79852
rect 158318 79716 158352 79756
rect 158346 79704 158352 79716
rect 158404 79704 158410 79756
rect 158640 79620 158668 79852
rect 158778 79756 158806 79908
rect 159128 79840 159134 79892
rect 159186 79840 159192 79892
rect 159496 79840 159502 79892
rect 159554 79840 159560 79892
rect 159606 79880 159634 79920
rect 159680 79908 159686 79960
rect 159738 79908 159744 79960
rect 160066 79880 160094 80056
rect 160802 79988 161198 80016
rect 160802 79960 160830 79988
rect 160784 79908 160790 79960
rect 160842 79908 160848 79960
rect 161060 79948 161066 79960
rect 161032 79908 161066 79948
rect 161118 79908 161124 79960
rect 159606 79852 160094 79880
rect 160140 79840 160146 79892
rect 160198 79840 160204 79892
rect 160416 79880 160422 79892
rect 160388 79840 160422 79880
rect 160474 79840 160480 79892
rect 160692 79840 160698 79892
rect 160750 79880 160756 79892
rect 160876 79880 160882 79892
rect 160750 79840 160784 79880
rect 158778 79716 158812 79756
rect 158806 79704 158812 79716
rect 158864 79704 158870 79756
rect 158530 79608 158536 79620
rect 158226 79580 158536 79608
rect 158530 79568 158536 79580
rect 158588 79568 158594 79620
rect 158622 79568 158628 79620
rect 158680 79568 158686 79620
rect 159146 79608 159174 79840
rect 159514 79688 159542 79840
rect 159514 79648 159548 79688
rect 159542 79636 159548 79648
rect 159600 79636 159606 79688
rect 159266 79608 159272 79620
rect 159146 79580 159272 79608
rect 159266 79568 159272 79580
rect 159324 79568 159330 79620
rect 160158 79608 160186 79840
rect 160278 79608 160284 79620
rect 160158 79580 160284 79608
rect 160278 79568 160284 79580
rect 160336 79568 160342 79620
rect 160388 79608 160416 79840
rect 160756 79756 160784 79840
rect 160848 79840 160882 79880
rect 160934 79840 160940 79892
rect 160848 79756 160876 79840
rect 160738 79704 160744 79756
rect 160796 79704 160802 79756
rect 160830 79704 160836 79756
rect 160888 79704 160894 79756
rect 161032 79620 161060 79908
rect 161170 79620 161198 79988
rect 163010 79988 163820 80016
rect 163010 79960 163038 79988
rect 161336 79948 161342 79960
rect 161308 79908 161342 79948
rect 161394 79908 161400 79960
rect 161428 79908 161434 79960
rect 161486 79908 161492 79960
rect 162532 79948 162538 79960
rect 161584 79920 161934 79948
rect 161308 79620 161336 79908
rect 161446 79880 161474 79908
rect 161446 79852 161520 79880
rect 161492 79756 161520 79852
rect 161474 79704 161480 79756
rect 161532 79704 161538 79756
rect 161584 79688 161612 79920
rect 161906 79892 161934 79920
rect 162504 79908 162538 79948
rect 162590 79908 162596 79960
rect 162624 79908 162630 79960
rect 162682 79908 162688 79960
rect 162808 79948 162814 79960
rect 162734 79920 162814 79948
rect 161704 79840 161710 79892
rect 161762 79880 161768 79892
rect 161762 79840 161796 79880
rect 161888 79840 161894 79892
rect 161946 79840 161952 79892
rect 162348 79840 162354 79892
rect 162406 79840 162412 79892
rect 161566 79636 161572 79688
rect 161624 79636 161630 79688
rect 160388 79580 160968 79608
rect 158438 79540 158444 79552
rect 157674 79512 158444 79540
rect 156748 79500 156754 79512
rect 158438 79500 158444 79512
rect 158496 79500 158502 79552
rect 160370 79500 160376 79552
rect 160428 79540 160434 79552
rect 160646 79540 160652 79552
rect 160428 79512 160652 79540
rect 160428 79500 160434 79512
rect 160646 79500 160652 79512
rect 160704 79500 160710 79552
rect 160940 79540 160968 79580
rect 161014 79568 161020 79620
rect 161072 79568 161078 79620
rect 161106 79568 161112 79620
rect 161164 79580 161198 79620
rect 161164 79568 161170 79580
rect 161290 79568 161296 79620
rect 161348 79568 161354 79620
rect 161198 79540 161204 79552
rect 160940 79512 161204 79540
rect 161198 79500 161204 79512
rect 161256 79500 161262 79552
rect 161474 79500 161480 79552
rect 161532 79540 161538 79552
rect 161768 79540 161796 79840
rect 162366 79620 162394 79840
rect 162504 79620 162532 79908
rect 162642 79880 162670 79908
rect 162596 79852 162670 79880
rect 162596 79824 162624 79852
rect 162578 79772 162584 79824
rect 162636 79772 162642 79824
rect 162734 79620 162762 79920
rect 162808 79908 162814 79920
rect 162866 79908 162872 79960
rect 162992 79908 162998 79960
rect 163050 79908 163056 79960
rect 163084 79840 163090 79892
rect 163142 79840 163148 79892
rect 163176 79840 163182 79892
rect 163234 79840 163240 79892
rect 163360 79840 163366 79892
rect 163418 79840 163424 79892
rect 163102 79688 163130 79840
rect 163038 79636 163044 79688
rect 163096 79648 163130 79688
rect 163194 79688 163222 79840
rect 163194 79648 163228 79688
rect 163096 79636 163102 79648
rect 163222 79636 163228 79648
rect 163280 79636 163286 79688
rect 162302 79568 162308 79620
rect 162360 79580 162394 79620
rect 162360 79568 162366 79580
rect 162486 79568 162492 79620
rect 162544 79568 162550 79620
rect 162670 79568 162676 79620
rect 162728 79580 162762 79620
rect 162728 79568 162734 79580
rect 162854 79568 162860 79620
rect 162912 79608 162918 79620
rect 163378 79608 163406 79840
rect 163636 79772 163642 79824
rect 163694 79772 163700 79824
rect 162912 79580 163406 79608
rect 163654 79620 163682 79772
rect 163792 79688 163820 79988
rect 163912 79908 163918 79960
rect 163970 79908 163976 79960
rect 164648 79948 164654 79960
rect 164482 79920 164654 79948
rect 163774 79636 163780 79688
rect 163832 79636 163838 79688
rect 163654 79580 163688 79620
rect 162912 79568 162918 79580
rect 163682 79568 163688 79580
rect 163740 79568 163746 79620
rect 163930 79608 163958 79908
rect 164096 79840 164102 79892
rect 164154 79840 164160 79892
rect 164114 79688 164142 79840
rect 164050 79636 164056 79688
rect 164108 79648 164142 79688
rect 164108 79636 164114 79648
rect 164142 79608 164148 79620
rect 163930 79580 164148 79608
rect 164142 79568 164148 79580
rect 164200 79568 164206 79620
rect 161532 79512 161796 79540
rect 161532 79500 161538 79512
rect 162118 79500 162124 79552
rect 162176 79540 162182 79552
rect 164326 79540 164332 79552
rect 162176 79512 164332 79540
rect 162176 79500 162182 79512
rect 164326 79500 164332 79512
rect 164384 79500 164390 79552
rect 164482 79540 164510 79920
rect 164648 79908 164654 79920
rect 164706 79908 164712 79960
rect 165200 79908 165206 79960
rect 165258 79908 165264 79960
rect 165660 79908 165666 79960
rect 165718 79908 165724 79960
rect 165752 79908 165758 79960
rect 165810 79908 165816 79960
rect 164556 79840 164562 79892
rect 164614 79840 164620 79892
rect 164740 79840 164746 79892
rect 164798 79840 164804 79892
rect 164574 79620 164602 79840
rect 164574 79580 164608 79620
rect 164602 79568 164608 79580
rect 164660 79568 164666 79620
rect 164758 79608 164786 79840
rect 165218 79756 165246 79908
rect 165292 79840 165298 79892
rect 165350 79880 165356 79892
rect 165350 79852 165568 79880
rect 165350 79840 165356 79852
rect 165384 79772 165390 79824
rect 165442 79772 165448 79824
rect 165218 79716 165252 79756
rect 165246 79704 165252 79716
rect 165304 79704 165310 79756
rect 165402 79620 165430 79772
rect 165540 79620 165568 79852
rect 165678 79620 165706 79908
rect 165770 79688 165798 79908
rect 165844 79840 165850 79892
rect 165902 79880 165908 79892
rect 166028 79880 166034 79892
rect 165902 79840 165936 79880
rect 165908 79756 165936 79840
rect 166000 79840 166034 79880
rect 166086 79840 166092 79892
rect 166304 79840 166310 79892
rect 166362 79840 166368 79892
rect 166396 79840 166402 79892
rect 166454 79840 166460 79892
rect 166000 79756 166028 79840
rect 166212 79772 166218 79824
rect 166270 79772 166276 79824
rect 165890 79704 165896 79756
rect 165948 79704 165954 79756
rect 165982 79704 165988 79756
rect 166040 79704 166046 79756
rect 166230 79688 166258 79772
rect 165770 79648 165804 79688
rect 165798 79636 165804 79648
rect 165856 79636 165862 79688
rect 166166 79636 166172 79688
rect 166224 79648 166258 79688
rect 166224 79636 166230 79648
rect 164758 79580 165016 79608
rect 165402 79580 165436 79620
rect 164988 79552 165016 79580
rect 165430 79568 165436 79580
rect 165488 79568 165494 79620
rect 165522 79568 165528 79620
rect 165580 79568 165586 79620
rect 165678 79580 165712 79620
rect 165706 79568 165712 79580
rect 165764 79568 165770 79620
rect 166322 79608 166350 79840
rect 165816 79580 166350 79608
rect 164786 79540 164792 79552
rect 164482 79512 164792 79540
rect 164786 79500 164792 79512
rect 164844 79500 164850 79552
rect 164970 79500 164976 79552
rect 165028 79500 165034 79552
rect 165338 79500 165344 79552
rect 165396 79540 165402 79552
rect 165816 79540 165844 79580
rect 165396 79512 165844 79540
rect 165396 79500 165402 79512
rect 166166 79500 166172 79552
rect 166224 79540 166230 79552
rect 166414 79540 166442 79840
rect 166224 79512 166442 79540
rect 166224 79500 166230 79512
rect 141200 79376 141510 79404
rect 145576 79444 153424 79472
rect 141200 79364 141206 79376
rect 145576 79336 145604 79444
rect 147674 79364 147680 79416
rect 147732 79404 147738 79416
rect 153396 79404 153424 79444
rect 153470 79432 153476 79484
rect 153528 79472 153534 79484
rect 166552 79472 166580 80056
rect 167472 80016 167500 80464
rect 179690 80424 179696 80436
rect 175246 80396 179696 80424
rect 175246 80356 175274 80396
rect 179690 80384 179696 80396
rect 179748 80384 179754 80436
rect 182146 80424 182174 80464
rect 182146 80396 183554 80424
rect 169036 80328 175274 80356
rect 183526 80356 183554 80396
rect 183526 80328 186314 80356
rect 169036 80152 169064 80328
rect 186286 80288 186314 80328
rect 292574 80288 292580 80300
rect 172394 80260 183554 80288
rect 186286 80260 292580 80288
rect 172394 80152 172422 80260
rect 179966 80220 179972 80232
rect 176028 80192 179972 80220
rect 176028 80152 176056 80192
rect 179966 80180 179972 80192
rect 180024 80180 180030 80232
rect 183526 80220 183554 80260
rect 292574 80248 292580 80260
rect 292632 80248 292638 80300
rect 316034 80220 316040 80232
rect 183526 80192 316040 80220
rect 316034 80180 316040 80192
rect 316092 80180 316098 80232
rect 179598 80152 179604 80164
rect 166966 79988 167500 80016
rect 167886 80124 169064 80152
rect 171290 80124 172422 80152
rect 172486 80124 176056 80152
rect 176626 80124 179604 80152
rect 166856 79948 166862 79960
rect 166690 79920 166862 79948
rect 166690 79552 166718 79920
rect 166856 79908 166862 79920
rect 166914 79908 166920 79960
rect 166764 79840 166770 79892
rect 166822 79840 166828 79892
rect 166782 79756 166810 79840
rect 166782 79716 166816 79756
rect 166810 79704 166816 79716
rect 166868 79704 166874 79756
rect 166810 79568 166816 79620
rect 166868 79608 166874 79620
rect 166966 79608 166994 79988
rect 167408 79908 167414 79960
rect 167466 79908 167472 79960
rect 167500 79908 167506 79960
rect 167558 79908 167564 79960
rect 167886 79948 167914 80124
rect 167610 79920 167914 79948
rect 167978 80056 170490 80084
rect 167132 79840 167138 79892
rect 167190 79840 167196 79892
rect 166868 79580 166994 79608
rect 167150 79608 167178 79840
rect 167426 79824 167454 79908
rect 167362 79772 167368 79824
rect 167420 79784 167454 79824
rect 167420 79772 167426 79784
rect 167518 79688 167546 79908
rect 167454 79636 167460 79688
rect 167512 79648 167546 79688
rect 167512 79636 167518 79648
rect 167270 79608 167276 79620
rect 167150 79580 167276 79608
rect 166868 79568 166874 79580
rect 167270 79568 167276 79580
rect 167328 79568 167334 79620
rect 166626 79500 166632 79552
rect 166684 79512 166718 79552
rect 166684 79500 166690 79512
rect 167610 79472 167638 79920
rect 167868 79840 167874 79892
rect 167926 79840 167932 79892
rect 167886 79620 167914 79840
rect 167978 79824 168006 80056
rect 168070 79988 168466 80016
rect 167960 79772 167966 79824
rect 168018 79772 168024 79824
rect 168070 79676 168098 79988
rect 168328 79908 168334 79960
rect 168386 79908 168392 79960
rect 168144 79840 168150 79892
rect 168202 79840 168208 79892
rect 168162 79812 168190 79840
rect 168162 79784 168236 79812
rect 168208 79756 168236 79784
rect 168190 79704 168196 79756
rect 168248 79704 168254 79756
rect 168346 79688 168374 79908
rect 168438 79892 168466 79988
rect 169156 79948 169162 79960
rect 169128 79908 169162 79948
rect 169214 79908 169220 79960
rect 169340 79908 169346 79960
rect 169398 79908 169404 79960
rect 169432 79908 169438 79960
rect 169490 79908 169496 79960
rect 170352 79908 170358 79960
rect 170410 79908 170416 79960
rect 168420 79840 168426 79892
rect 168478 79840 168484 79892
rect 168604 79840 168610 79892
rect 168662 79880 168668 79892
rect 168662 79852 168972 79880
rect 168662 79840 168668 79852
rect 168512 79812 168518 79824
rect 168024 79648 168098 79676
rect 167886 79580 167920 79620
rect 167914 79568 167920 79580
rect 167972 79568 167978 79620
rect 168024 79540 168052 79648
rect 168282 79636 168288 79688
rect 168340 79648 168374 79688
rect 168438 79784 168518 79812
rect 168340 79636 168346 79648
rect 168098 79568 168104 79620
rect 168156 79608 168162 79620
rect 168438 79608 168466 79784
rect 168512 79772 168518 79784
rect 168570 79772 168576 79824
rect 168696 79772 168702 79824
rect 168754 79772 168760 79824
rect 168156 79580 168466 79608
rect 168156 79568 168162 79580
rect 168558 79568 168564 79620
rect 168616 79608 168622 79620
rect 168714 79608 168742 79772
rect 168944 79688 168972 79852
rect 169128 79688 169156 79908
rect 169248 79880 169254 79892
rect 169220 79840 169254 79880
rect 169306 79840 169312 79892
rect 169220 79756 169248 79840
rect 169358 79756 169386 79908
rect 169202 79704 169208 79756
rect 169260 79704 169266 79756
rect 169294 79704 169300 79756
rect 169352 79716 169386 79756
rect 169450 79756 169478 79908
rect 169616 79840 169622 79892
rect 169674 79840 169680 79892
rect 169892 79840 169898 79892
rect 169950 79840 169956 79892
rect 169984 79840 169990 79892
rect 170042 79840 170048 79892
rect 169450 79716 169484 79756
rect 169352 79704 169358 79716
rect 169478 79704 169484 79716
rect 169536 79704 169542 79756
rect 168926 79636 168932 79688
rect 168984 79636 168990 79688
rect 169110 79636 169116 79688
rect 169168 79636 169174 79688
rect 168616 79580 168742 79608
rect 168616 79568 168622 79580
rect 168374 79540 168380 79552
rect 168024 79512 168380 79540
rect 168374 79500 168380 79512
rect 168432 79500 168438 79552
rect 169386 79500 169392 79552
rect 169444 79540 169450 79552
rect 169634 79540 169662 79840
rect 169754 79568 169760 79620
rect 169812 79608 169818 79620
rect 169910 79608 169938 79840
rect 169812 79580 169938 79608
rect 169812 79568 169818 79580
rect 170002 79552 170030 79840
rect 170076 79772 170082 79824
rect 170134 79812 170140 79824
rect 170134 79772 170168 79812
rect 170140 79688 170168 79772
rect 170122 79636 170128 79688
rect 170180 79636 170186 79688
rect 169444 79512 169662 79540
rect 169444 79500 169450 79512
rect 169938 79500 169944 79552
rect 169996 79512 170030 79552
rect 169996 79500 170002 79512
rect 170122 79500 170128 79552
rect 170180 79540 170186 79552
rect 170370 79540 170398 79908
rect 170462 79812 170490 80056
rect 170628 79908 170634 79960
rect 170686 79908 170692 79960
rect 170812 79908 170818 79960
rect 170870 79908 170876 79960
rect 170996 79908 171002 79960
rect 171054 79908 171060 79960
rect 170646 79880 170674 79908
rect 170646 79852 170720 79880
rect 170582 79812 170588 79824
rect 170462 79784 170588 79812
rect 170582 79772 170588 79784
rect 170640 79772 170646 79824
rect 170490 79704 170496 79756
rect 170548 79704 170554 79756
rect 170508 79552 170536 79704
rect 170582 79568 170588 79620
rect 170640 79608 170646 79620
rect 170692 79608 170720 79852
rect 170640 79580 170720 79608
rect 170640 79568 170646 79580
rect 170180 79512 170398 79540
rect 170180 79500 170186 79512
rect 170490 79500 170496 79552
rect 170548 79500 170554 79552
rect 170674 79500 170680 79552
rect 170732 79540 170738 79552
rect 170830 79540 170858 79908
rect 171014 79824 171042 79908
rect 171014 79784 171048 79824
rect 171042 79772 171048 79784
rect 171100 79772 171106 79824
rect 170950 79636 170956 79688
rect 171008 79676 171014 79688
rect 171290 79676 171318 80124
rect 171364 79908 171370 79960
rect 171422 79948 171428 79960
rect 172486 79948 172514 80124
rect 173268 80056 174722 80084
rect 173268 79960 173296 80056
rect 171422 79920 172514 79948
rect 171422 79908 171428 79920
rect 172560 79908 172566 79960
rect 172618 79908 172624 79960
rect 173020 79908 173026 79960
rect 173078 79908 173084 79960
rect 173204 79908 173210 79960
rect 173262 79920 173296 79960
rect 173262 79908 173268 79920
rect 171824 79880 171830 79892
rect 171796 79840 171830 79880
rect 171882 79840 171888 79892
rect 172578 79880 172606 79908
rect 172486 79852 172606 79880
rect 171796 79756 171824 79840
rect 172008 79772 172014 79824
rect 172066 79772 172072 79824
rect 172192 79772 172198 79824
rect 172250 79772 172256 79824
rect 172284 79772 172290 79824
rect 172342 79772 172348 79824
rect 171778 79704 171784 79756
rect 171836 79704 171842 79756
rect 172026 79744 172054 79772
rect 171980 79716 172054 79744
rect 171008 79648 171318 79676
rect 171008 79636 171014 79648
rect 171980 79620 172008 79716
rect 171962 79568 171968 79620
rect 172020 79568 172026 79620
rect 172210 79608 172238 79772
rect 172164 79580 172238 79608
rect 172164 79552 172192 79580
rect 172302 79552 172330 79772
rect 172486 79620 172514 79852
rect 172836 79840 172842 79892
rect 172894 79840 172900 79892
rect 172854 79744 172882 79840
rect 172422 79568 172428 79620
rect 172480 79580 172514 79620
rect 172624 79716 172882 79744
rect 172480 79568 172486 79580
rect 170732 79512 170858 79540
rect 170732 79500 170738 79512
rect 172146 79500 172152 79552
rect 172204 79500 172210 79552
rect 172238 79500 172244 79552
rect 172296 79512 172330 79552
rect 172624 79540 172652 79716
rect 172882 79636 172888 79688
rect 172940 79676 172946 79688
rect 173038 79676 173066 79908
rect 173480 79840 173486 79892
rect 173538 79840 173544 79892
rect 173848 79840 173854 79892
rect 173906 79840 173912 79892
rect 174216 79880 174222 79892
rect 174188 79840 174222 79880
rect 174274 79840 174280 79892
rect 174308 79840 174314 79892
rect 174366 79880 174372 79892
rect 174366 79840 174400 79880
rect 172940 79648 173066 79676
rect 172940 79636 172946 79648
rect 173158 79636 173164 79688
rect 173216 79676 173222 79688
rect 173498 79676 173526 79840
rect 173866 79688 173894 79840
rect 174188 79688 174216 79840
rect 174372 79688 174400 79840
rect 174492 79812 174498 79824
rect 174464 79772 174498 79812
rect 174550 79772 174556 79824
rect 174464 79688 174492 79772
rect 173216 79648 173526 79676
rect 173216 79636 173222 79648
rect 173848 79636 173854 79688
rect 173906 79636 173912 79688
rect 174170 79636 174176 79688
rect 174228 79636 174234 79688
rect 174354 79636 174360 79688
rect 174412 79636 174418 79688
rect 174446 79636 174452 79688
rect 174504 79636 174510 79688
rect 174694 79608 174722 80056
rect 176626 79960 176654 80124
rect 179598 80112 179604 80124
rect 179656 80112 179662 80164
rect 180150 80152 180156 80164
rect 179800 80124 180156 80152
rect 179800 80084 179828 80124
rect 180150 80112 180156 80124
rect 180208 80112 180214 80164
rect 180242 80112 180248 80164
rect 180300 80152 180306 80164
rect 373994 80152 374000 80164
rect 180300 80124 374000 80152
rect 180300 80112 180306 80124
rect 373994 80112 374000 80124
rect 374052 80112 374058 80164
rect 176718 80056 179828 80084
rect 176718 79960 176746 80056
rect 179874 80044 179880 80096
rect 179932 80084 179938 80096
rect 547966 80084 547972 80096
rect 179932 80056 547972 80084
rect 179932 80044 179938 80056
rect 547966 80044 547972 80056
rect 548024 80044 548030 80096
rect 179690 79976 179696 80028
rect 179748 80016 179754 80028
rect 179748 79988 186314 80016
rect 179748 79976 179754 79988
rect 174768 79908 174774 79960
rect 174826 79908 174832 79960
rect 175136 79908 175142 79960
rect 175194 79908 175200 79960
rect 175412 79908 175418 79960
rect 175470 79908 175476 79960
rect 175596 79908 175602 79960
rect 175654 79908 175660 79960
rect 175964 79908 175970 79960
rect 176022 79948 176028 79960
rect 176022 79920 176378 79948
rect 176022 79908 176028 79920
rect 174786 79676 174814 79908
rect 174906 79676 174912 79688
rect 174786 79648 174912 79676
rect 174906 79636 174912 79648
rect 174964 79636 174970 79688
rect 174998 79636 175004 79688
rect 175056 79676 175062 79688
rect 175154 79676 175182 79908
rect 175320 79840 175326 79892
rect 175378 79840 175384 79892
rect 175056 79648 175182 79676
rect 175056 79636 175062 79648
rect 175338 79620 175366 79840
rect 175430 79756 175458 79908
rect 175614 79756 175642 79908
rect 175872 79840 175878 79892
rect 175930 79840 175936 79892
rect 176056 79880 176062 79892
rect 175982 79852 176062 79880
rect 175430 79716 175464 79756
rect 175458 79704 175464 79716
rect 175516 79704 175522 79756
rect 175550 79704 175556 79756
rect 175608 79716 175642 79756
rect 175608 79704 175614 79716
rect 175890 79620 175918 79840
rect 175982 79676 176010 79852
rect 176056 79840 176062 79852
rect 176114 79840 176120 79892
rect 176240 79840 176246 79892
rect 176298 79840 176304 79892
rect 176148 79772 176154 79824
rect 176206 79772 176212 79824
rect 176056 79676 176062 79688
rect 175982 79648 176062 79676
rect 176056 79636 176062 79648
rect 176114 79636 176120 79688
rect 175182 79608 175188 79620
rect 174694 79580 175188 79608
rect 175182 79568 175188 79580
rect 175240 79568 175246 79620
rect 175338 79580 175372 79620
rect 175366 79568 175372 79580
rect 175424 79568 175430 79620
rect 175890 79580 175924 79620
rect 175918 79568 175924 79580
rect 175976 79568 175982 79620
rect 173158 79540 173164 79552
rect 172624 79512 173164 79540
rect 172296 79500 172302 79512
rect 173158 79500 173164 79512
rect 173216 79500 173222 79552
rect 176166 79540 176194 79772
rect 176258 79676 176286 79840
rect 176350 79744 176378 79920
rect 176608 79908 176614 79960
rect 176666 79908 176672 79960
rect 176700 79908 176706 79960
rect 176758 79908 176764 79960
rect 177068 79908 177074 79960
rect 177126 79908 177132 79960
rect 177160 79908 177166 79960
rect 177218 79908 177224 79960
rect 177528 79908 177534 79960
rect 177586 79908 177592 79960
rect 177620 79908 177626 79960
rect 177678 79948 177684 79960
rect 177896 79948 177902 79960
rect 177678 79920 177804 79948
rect 177678 79908 177684 79920
rect 176424 79840 176430 79892
rect 176482 79840 176488 79892
rect 176442 79812 176470 79840
rect 176746 79812 176752 79824
rect 176442 79784 176752 79812
rect 176746 79772 176752 79784
rect 176804 79772 176810 79824
rect 176562 79744 176568 79756
rect 176350 79716 176568 79744
rect 176562 79704 176568 79716
rect 176620 79704 176626 79756
rect 176654 79676 176660 79688
rect 176258 79648 176660 79676
rect 176654 79636 176660 79648
rect 176712 79636 176718 79688
rect 177086 79620 177114 79908
rect 177178 79676 177206 79908
rect 177252 79840 177258 79892
rect 177310 79840 177316 79892
rect 177546 79880 177574 79908
rect 177546 79852 177712 79880
rect 177270 79812 177298 79840
rect 177574 79812 177580 79824
rect 177270 79784 177580 79812
rect 177574 79772 177580 79784
rect 177632 79772 177638 79824
rect 177684 79688 177712 79852
rect 177776 79688 177804 79920
rect 177868 79908 177902 79948
rect 177954 79908 177960 79960
rect 178080 79908 178086 79960
rect 178138 79908 178144 79960
rect 178724 79908 178730 79960
rect 178782 79908 178788 79960
rect 179184 79908 179190 79960
rect 179242 79948 179248 79960
rect 179506 79948 179512 79960
rect 179242 79920 179512 79948
rect 179242 79908 179248 79920
rect 179506 79908 179512 79920
rect 179564 79908 179570 79960
rect 177868 79756 177896 79908
rect 178098 79824 178126 79908
rect 178172 79840 178178 79892
rect 178230 79840 178236 79892
rect 178540 79840 178546 79892
rect 178598 79840 178604 79892
rect 178080 79772 178086 79824
rect 178138 79772 178144 79824
rect 177850 79704 177856 79756
rect 177908 79704 177914 79756
rect 177298 79676 177304 79688
rect 177178 79648 177304 79676
rect 177298 79636 177304 79648
rect 177356 79636 177362 79688
rect 177666 79636 177672 79688
rect 177724 79636 177730 79688
rect 177758 79636 177764 79688
rect 177816 79636 177822 79688
rect 177086 79580 177120 79620
rect 177114 79568 177120 79580
rect 177172 79568 177178 79620
rect 177206 79568 177212 79620
rect 177264 79608 177270 79620
rect 177942 79608 177948 79620
rect 177264 79580 177948 79608
rect 177264 79568 177270 79580
rect 177942 79568 177948 79580
rect 178000 79568 178006 79620
rect 178034 79568 178040 79620
rect 178092 79608 178098 79620
rect 178190 79608 178218 79840
rect 178402 79636 178408 79688
rect 178460 79676 178466 79688
rect 178558 79676 178586 79840
rect 178460 79648 178586 79676
rect 178460 79636 178466 79648
rect 178092 79580 178218 79608
rect 178092 79568 178098 79580
rect 178494 79568 178500 79620
rect 178552 79608 178558 79620
rect 178742 79608 178770 79908
rect 178908 79840 178914 79892
rect 178966 79880 178972 79892
rect 179690 79880 179696 79892
rect 178966 79852 179696 79880
rect 178966 79840 178972 79852
rect 179690 79840 179696 79852
rect 179748 79840 179754 79892
rect 179000 79772 179006 79824
rect 179058 79772 179064 79824
rect 186286 79812 186314 79988
rect 362954 79812 362960 79824
rect 186286 79784 362960 79812
rect 362954 79772 362960 79784
rect 363012 79772 363018 79824
rect 178552 79580 178770 79608
rect 179018 79608 179046 79772
rect 179138 79704 179144 79756
rect 179196 79744 179202 79756
rect 179782 79744 179788 79756
rect 179196 79716 179788 79744
rect 179196 79704 179202 79716
rect 179782 79704 179788 79716
rect 179840 79704 179846 79756
rect 179966 79636 179972 79688
rect 180024 79676 180030 79688
rect 523126 79676 523132 79688
rect 180024 79648 523132 79676
rect 180024 79636 180030 79648
rect 523126 79636 523132 79648
rect 523184 79636 523190 79688
rect 179138 79608 179144 79620
rect 179018 79580 179144 79608
rect 178552 79568 178558 79580
rect 179138 79568 179144 79580
rect 179196 79568 179202 79620
rect 189718 79540 189724 79552
rect 176166 79512 189724 79540
rect 189718 79500 189724 79512
rect 189776 79500 189782 79552
rect 153528 79444 164740 79472
rect 166552 79444 167638 79472
rect 153528 79432 153534 79444
rect 164326 79404 164332 79416
rect 147732 79376 149928 79404
rect 153396 79376 164332 79404
rect 147732 79364 147738 79376
rect 149606 79336 149612 79348
rect 3936 79308 118694 79336
rect 125566 79308 126974 79336
rect 3936 79296 3942 79308
rect 118666 79200 118694 79308
rect 126946 79268 126974 79308
rect 134076 79308 145604 79336
rect 145668 79308 149612 79336
rect 134076 79268 134104 79308
rect 126946 79240 134104 79268
rect 134242 79228 134248 79280
rect 134300 79268 134306 79280
rect 145668 79268 145696 79308
rect 149606 79296 149612 79308
rect 149664 79296 149670 79348
rect 149900 79268 149928 79376
rect 164326 79364 164332 79376
rect 164384 79364 164390 79416
rect 164712 79336 164740 79444
rect 167730 79432 167736 79484
rect 167788 79472 167794 79484
rect 167788 79444 171548 79472
rect 167788 79432 167794 79444
rect 165614 79404 165620 79416
rect 164896 79376 165620 79404
rect 164896 79336 164924 79376
rect 165614 79364 165620 79376
rect 165672 79364 165678 79416
rect 168282 79364 168288 79416
rect 168340 79404 168346 79416
rect 171410 79404 171416 79416
rect 168340 79376 171416 79404
rect 168340 79364 168346 79376
rect 171410 79364 171416 79376
rect 171468 79364 171474 79416
rect 171520 79404 171548 79444
rect 171594 79432 171600 79484
rect 171652 79472 171658 79484
rect 171870 79472 171876 79484
rect 171652 79444 171876 79472
rect 171652 79432 171658 79444
rect 171870 79432 171876 79444
rect 171928 79432 171934 79484
rect 172054 79432 172060 79484
rect 172112 79472 172118 79484
rect 178218 79472 178224 79484
rect 172112 79444 178224 79472
rect 172112 79432 172118 79444
rect 178218 79432 178224 79444
rect 178276 79432 178282 79484
rect 178862 79404 178868 79416
rect 171520 79376 178868 79404
rect 178862 79364 178868 79376
rect 178920 79364 178926 79416
rect 155052 79308 164234 79336
rect 164712 79308 164924 79336
rect 164988 79308 172514 79336
rect 153470 79268 153476 79280
rect 134300 79240 145696 79268
rect 145760 79240 149054 79268
rect 149900 79240 153476 79268
rect 134300 79228 134306 79240
rect 118666 79172 126974 79200
rect 126946 79132 126974 79172
rect 138290 79160 138296 79212
rect 138348 79200 138354 79212
rect 138750 79200 138756 79212
rect 138348 79172 138756 79200
rect 138348 79160 138354 79172
rect 138750 79160 138756 79172
rect 138808 79160 138814 79212
rect 139118 79160 139124 79212
rect 139176 79200 139182 79212
rect 141326 79200 141332 79212
rect 139176 79172 141332 79200
rect 139176 79160 139182 79172
rect 141326 79160 141332 79172
rect 141384 79160 141390 79212
rect 145760 79132 145788 79240
rect 149026 79200 149054 79240
rect 153470 79228 153476 79240
rect 153528 79228 153534 79280
rect 155052 79200 155080 79308
rect 157794 79228 157800 79280
rect 157852 79268 157858 79280
rect 162762 79268 162768 79280
rect 157852 79240 162768 79268
rect 157852 79228 157858 79240
rect 162762 79228 162768 79240
rect 162820 79228 162826 79280
rect 149026 79172 155080 79200
rect 159174 79160 159180 79212
rect 159232 79200 159238 79212
rect 161290 79200 161296 79212
rect 159232 79172 161296 79200
rect 159232 79160 159238 79172
rect 161290 79160 161296 79172
rect 161348 79160 161354 79212
rect 162026 79160 162032 79212
rect 162084 79200 162090 79212
rect 162394 79200 162400 79212
rect 162084 79172 162400 79200
rect 162084 79160 162090 79172
rect 162394 79160 162400 79172
rect 162452 79160 162458 79212
rect 164206 79200 164234 79308
rect 164988 79200 165016 79308
rect 165614 79228 165620 79280
rect 165672 79268 165678 79280
rect 167730 79268 167736 79280
rect 165672 79240 167736 79268
rect 165672 79228 165678 79240
rect 167730 79228 167736 79240
rect 167788 79228 167794 79280
rect 168558 79228 168564 79280
rect 168616 79268 168622 79280
rect 171870 79268 171876 79280
rect 168616 79240 171876 79268
rect 168616 79228 168622 79240
rect 171870 79228 171876 79240
rect 171928 79228 171934 79280
rect 172486 79268 172514 79308
rect 175274 79296 175280 79348
rect 175332 79336 175338 79348
rect 176194 79336 176200 79348
rect 175332 79308 176200 79336
rect 175332 79296 175338 79308
rect 176194 79296 176200 79308
rect 176252 79296 176258 79348
rect 176286 79296 176292 79348
rect 176344 79336 176350 79348
rect 178126 79336 178132 79348
rect 176344 79308 178132 79336
rect 176344 79296 176350 79308
rect 178126 79296 178132 79308
rect 178184 79296 178190 79348
rect 179782 79296 179788 79348
rect 179840 79336 179846 79348
rect 527174 79336 527180 79348
rect 179840 79308 527180 79336
rect 179840 79296 179846 79308
rect 527174 79296 527180 79308
rect 527232 79296 527238 79348
rect 178678 79268 178684 79280
rect 172486 79240 178684 79268
rect 178678 79228 178684 79240
rect 178736 79228 178742 79280
rect 180150 79228 180156 79280
rect 180208 79268 180214 79280
rect 192754 79268 192760 79280
rect 180208 79240 192760 79268
rect 180208 79228 180214 79240
rect 192754 79228 192760 79240
rect 192812 79228 192818 79280
rect 164206 79172 165016 79200
rect 166902 79160 166908 79212
rect 166960 79200 166966 79212
rect 170950 79200 170956 79212
rect 166960 79172 170956 79200
rect 166960 79160 166966 79172
rect 170950 79160 170956 79172
rect 171008 79160 171014 79212
rect 171410 79160 171416 79212
rect 171468 79200 171474 79212
rect 175642 79200 175648 79212
rect 171468 79172 175648 79200
rect 171468 79160 171474 79172
rect 175642 79160 175648 79172
rect 175700 79160 175706 79212
rect 176194 79160 176200 79212
rect 176252 79200 176258 79212
rect 178310 79200 178316 79212
rect 176252 79172 178316 79200
rect 176252 79160 176258 79172
rect 178310 79160 178316 79172
rect 178368 79160 178374 79212
rect 180058 79160 180064 79212
rect 180116 79200 180122 79212
rect 192938 79200 192944 79212
rect 180116 79172 192944 79200
rect 180116 79160 180122 79172
rect 192938 79160 192944 79172
rect 192996 79160 193002 79212
rect 150526 79132 150532 79144
rect 126946 79104 145788 79132
rect 150406 79104 150532 79132
rect 130470 79024 130476 79076
rect 130528 79064 130534 79076
rect 134242 79064 134248 79076
rect 130528 79036 134248 79064
rect 130528 79024 130534 79036
rect 134242 79024 134248 79036
rect 134300 79024 134306 79076
rect 135254 79024 135260 79076
rect 135312 79064 135318 79076
rect 137094 79064 137100 79076
rect 135312 79036 137100 79064
rect 135312 79024 135318 79036
rect 137094 79024 137100 79036
rect 137152 79024 137158 79076
rect 139854 79024 139860 79076
rect 139912 79064 139918 79076
rect 140130 79064 140136 79076
rect 139912 79036 140136 79064
rect 139912 79024 139918 79036
rect 140130 79024 140136 79036
rect 140188 79024 140194 79076
rect 144914 79024 144920 79076
rect 144972 79064 144978 79076
rect 147674 79064 147680 79076
rect 144972 79036 147680 79064
rect 144972 79024 144978 79036
rect 147674 79024 147680 79036
rect 147732 79024 147738 79076
rect 3786 78956 3792 79008
rect 3844 78996 3850 79008
rect 133874 78996 133880 79008
rect 3844 78968 133880 78996
rect 3844 78956 3850 78968
rect 133874 78956 133880 78968
rect 133932 78956 133938 79008
rect 138658 78956 138664 79008
rect 138716 78996 138722 79008
rect 138716 78968 145604 78996
rect 138716 78956 138722 78968
rect 131666 78888 131672 78940
rect 131724 78928 131730 78940
rect 144914 78928 144920 78940
rect 131724 78900 144920 78928
rect 131724 78888 131730 78900
rect 144914 78888 144920 78900
rect 144972 78888 144978 78940
rect 145576 78928 145604 78968
rect 147214 78956 147220 79008
rect 147272 78996 147278 79008
rect 150406 78996 150434 79104
rect 150526 79092 150532 79104
rect 150584 79092 150590 79144
rect 164326 79092 164332 79144
rect 164384 79132 164390 79144
rect 168282 79132 168288 79144
rect 164384 79104 168288 79132
rect 164384 79092 164390 79104
rect 168282 79092 168288 79104
rect 168340 79092 168346 79144
rect 169386 79092 169392 79144
rect 169444 79132 169450 79144
rect 169444 79104 172192 79132
rect 169444 79092 169450 79104
rect 158778 79036 168696 79064
rect 147272 78968 150434 78996
rect 147272 78956 147278 78968
rect 156230 78956 156236 79008
rect 156288 78996 156294 79008
rect 158778 78996 158806 79036
rect 156288 78968 158806 78996
rect 156288 78956 156294 78968
rect 159910 78956 159916 79008
rect 159968 78996 159974 79008
rect 162118 78996 162124 79008
rect 159968 78968 162124 78996
rect 159968 78956 159974 78968
rect 162118 78956 162124 78968
rect 162176 78956 162182 79008
rect 162210 78956 162216 79008
rect 162268 78996 162274 79008
rect 162394 78996 162400 79008
rect 162268 78968 162400 78996
rect 162268 78956 162274 78968
rect 162394 78956 162400 78968
rect 162452 78956 162458 79008
rect 162762 78956 162768 79008
rect 162820 78996 162826 79008
rect 168558 78996 168564 79008
rect 162820 78968 168564 78996
rect 162820 78956 162826 78968
rect 168558 78956 168564 78968
rect 168616 78956 168622 79008
rect 168668 78996 168696 79036
rect 169662 79024 169668 79076
rect 169720 79064 169726 79076
rect 172054 79064 172060 79076
rect 169720 79036 172060 79064
rect 169720 79024 169726 79036
rect 172054 79024 172060 79036
rect 172112 79024 172118 79076
rect 172164 79064 172192 79104
rect 172606 79092 172612 79144
rect 172664 79132 172670 79144
rect 176746 79132 176752 79144
rect 172664 79104 176752 79132
rect 172664 79092 172670 79104
rect 176746 79092 176752 79104
rect 176804 79092 176810 79144
rect 180702 79092 180708 79144
rect 180760 79132 180766 79144
rect 201494 79132 201500 79144
rect 180760 79104 201500 79132
rect 180760 79092 180766 79104
rect 201494 79092 201500 79104
rect 201552 79092 201558 79144
rect 274634 79064 274640 79076
rect 172164 79036 274640 79064
rect 274634 79024 274640 79036
rect 274692 79024 274698 79076
rect 171134 78996 171140 79008
rect 168668 78968 171140 78996
rect 171134 78956 171140 78968
rect 171192 78956 171198 79008
rect 171502 78956 171508 79008
rect 171560 78956 171566 79008
rect 173250 78956 173256 79008
rect 173308 78996 173314 79008
rect 178586 78996 178592 79008
rect 173308 78968 178592 78996
rect 173308 78956 173314 78968
rect 178586 78956 178592 78968
rect 178644 78956 178650 79008
rect 145576 78900 151814 78928
rect 3510 78820 3516 78872
rect 3568 78860 3574 78872
rect 147214 78860 147220 78872
rect 3568 78832 147220 78860
rect 3568 78820 3574 78832
rect 147214 78820 147220 78832
rect 147272 78820 147278 78872
rect 151786 78860 151814 78900
rect 151878 78900 169156 78928
rect 151878 78860 151906 78900
rect 151786 78832 151906 78860
rect 157702 78820 157708 78872
rect 157760 78860 157766 78872
rect 157978 78860 157984 78872
rect 157760 78832 157984 78860
rect 157760 78820 157766 78832
rect 157978 78820 157984 78832
rect 158036 78820 158042 78872
rect 158254 78820 158260 78872
rect 158312 78860 158318 78872
rect 169128 78860 169156 78900
rect 171042 78888 171048 78940
rect 171100 78928 171106 78940
rect 171520 78928 171548 78956
rect 171100 78900 171548 78928
rect 171100 78888 171106 78900
rect 172606 78888 172612 78940
rect 172664 78928 172670 78940
rect 313274 78928 313280 78940
rect 172664 78900 313280 78928
rect 172664 78888 172670 78900
rect 313274 78888 313280 78900
rect 313332 78888 313338 78940
rect 158312 78832 169064 78860
rect 169128 78832 171502 78860
rect 158312 78820 158318 78832
rect 133874 78752 133880 78804
rect 133932 78792 133938 78804
rect 138658 78792 138664 78804
rect 133932 78764 138664 78792
rect 133932 78752 133938 78764
rect 138658 78752 138664 78764
rect 138716 78752 138722 78804
rect 150526 78752 150532 78804
rect 150584 78792 150590 78804
rect 165614 78792 165620 78804
rect 150584 78764 165620 78792
rect 150584 78752 150590 78764
rect 165614 78752 165620 78764
rect 165672 78752 165678 78804
rect 169036 78792 169064 78832
rect 169662 78792 169668 78804
rect 169036 78764 169668 78792
rect 169662 78752 169668 78764
rect 169720 78752 169726 78804
rect 171474 78792 171502 78832
rect 171870 78820 171876 78872
rect 171928 78860 171934 78872
rect 178494 78860 178500 78872
rect 171928 78832 178500 78860
rect 171928 78820 171934 78832
rect 178494 78820 178500 78832
rect 178552 78820 178558 78872
rect 178402 78792 178408 78804
rect 171474 78764 178408 78792
rect 178402 78752 178408 78764
rect 178460 78752 178466 78804
rect 178586 78752 178592 78804
rect 178644 78792 178650 78804
rect 179230 78792 179236 78804
rect 178644 78764 179236 78792
rect 178644 78752 178650 78764
rect 179230 78752 179236 78764
rect 179288 78752 179294 78804
rect 126238 78684 126244 78736
rect 126296 78724 126302 78736
rect 132678 78724 132684 78736
rect 126296 78696 132684 78724
rect 126296 78684 126302 78696
rect 132678 78684 132684 78696
rect 132736 78684 132742 78736
rect 157058 78684 157064 78736
rect 157116 78724 157122 78736
rect 157978 78724 157984 78736
rect 157116 78696 157984 78724
rect 157116 78684 157122 78696
rect 157978 78684 157984 78696
rect 158036 78684 158042 78736
rect 168282 78684 168288 78736
rect 168340 78724 168346 78736
rect 177850 78724 177856 78736
rect 168340 78696 169524 78724
rect 168340 78684 168346 78696
rect 126330 78616 126336 78668
rect 126388 78656 126394 78668
rect 133230 78656 133236 78668
rect 126388 78628 133236 78656
rect 126388 78616 126394 78628
rect 133230 78616 133236 78628
rect 133288 78616 133294 78668
rect 133322 78616 133328 78668
rect 133380 78656 133386 78668
rect 133874 78656 133880 78668
rect 133380 78628 133880 78656
rect 133380 78616 133386 78628
rect 133874 78616 133880 78628
rect 133932 78616 133938 78668
rect 137094 78616 137100 78668
rect 137152 78656 137158 78668
rect 138014 78656 138020 78668
rect 137152 78628 138020 78656
rect 137152 78616 137158 78628
rect 138014 78616 138020 78628
rect 138072 78616 138078 78668
rect 151906 78616 151912 78668
rect 151964 78656 151970 78668
rect 169386 78656 169392 78668
rect 151964 78628 169392 78656
rect 151964 78616 151970 78628
rect 169386 78616 169392 78628
rect 169444 78616 169450 78668
rect 169496 78656 169524 78696
rect 173866 78696 177856 78724
rect 173866 78656 173894 78696
rect 177850 78684 177856 78696
rect 177908 78684 177914 78736
rect 169496 78628 173894 78656
rect 174630 78616 174636 78668
rect 174688 78656 174694 78668
rect 174814 78656 174820 78668
rect 174688 78628 174820 78656
rect 174688 78616 174694 78628
rect 174814 78616 174820 78628
rect 174872 78616 174878 78668
rect 174906 78616 174912 78668
rect 174964 78656 174970 78668
rect 175182 78656 175188 78668
rect 174964 78628 175188 78656
rect 174964 78616 174970 78628
rect 175182 78616 175188 78628
rect 175240 78616 175246 78668
rect 176194 78616 176200 78668
rect 176252 78656 176258 78668
rect 176562 78656 176568 78668
rect 176252 78628 176568 78656
rect 176252 78616 176258 78628
rect 176562 78616 176568 78628
rect 176620 78616 176626 78668
rect 127618 78548 127624 78600
rect 127676 78588 127682 78600
rect 140314 78588 140320 78600
rect 127676 78560 140320 78588
rect 127676 78548 127682 78560
rect 140314 78548 140320 78560
rect 140372 78548 140378 78600
rect 149698 78548 149704 78600
rect 149756 78588 149762 78600
rect 156690 78588 156696 78600
rect 149756 78560 156696 78588
rect 149756 78548 149762 78560
rect 156690 78548 156696 78560
rect 156748 78548 156754 78600
rect 168098 78548 168104 78600
rect 168156 78588 168162 78600
rect 176470 78588 176476 78600
rect 168156 78560 176476 78588
rect 168156 78548 168162 78560
rect 176470 78548 176476 78560
rect 176528 78548 176534 78600
rect 177114 78548 177120 78600
rect 177172 78588 177178 78600
rect 192478 78588 192484 78600
rect 177172 78560 192484 78588
rect 177172 78548 177178 78560
rect 192478 78548 192484 78560
rect 192536 78548 192542 78600
rect 143718 78480 143724 78532
rect 143776 78520 143782 78532
rect 144178 78520 144184 78532
rect 143776 78492 144184 78520
rect 143776 78480 143782 78492
rect 144178 78480 144184 78492
rect 144236 78480 144242 78532
rect 153378 78480 153384 78532
rect 153436 78520 153442 78532
rect 166810 78520 166816 78532
rect 153436 78492 166816 78520
rect 153436 78480 153442 78492
rect 166810 78480 166816 78492
rect 166868 78480 166874 78532
rect 170950 78480 170956 78532
rect 171008 78520 171014 78532
rect 171502 78520 171508 78532
rect 171008 78492 171508 78520
rect 171008 78480 171014 78492
rect 171502 78480 171508 78492
rect 171560 78480 171566 78532
rect 177022 78480 177028 78532
rect 177080 78520 177086 78532
rect 192570 78520 192576 78532
rect 177080 78492 192576 78520
rect 177080 78480 177086 78492
rect 192570 78480 192576 78492
rect 192628 78480 192634 78532
rect 129090 78412 129096 78464
rect 129148 78452 129154 78464
rect 138842 78452 138848 78464
rect 129148 78424 138848 78452
rect 129148 78412 129154 78424
rect 138842 78412 138848 78424
rect 138900 78412 138906 78464
rect 162578 78412 162584 78464
rect 162636 78452 162642 78464
rect 177666 78452 177672 78464
rect 162636 78424 177672 78452
rect 162636 78412 162642 78424
rect 177666 78412 177672 78424
rect 177724 78412 177730 78464
rect 177942 78412 177948 78464
rect 178000 78452 178006 78464
rect 189350 78452 189356 78464
rect 178000 78424 189356 78452
rect 178000 78412 178006 78424
rect 189350 78412 189356 78424
rect 189408 78412 189414 78464
rect 130010 78344 130016 78396
rect 130068 78384 130074 78396
rect 131114 78384 131120 78396
rect 130068 78356 131120 78384
rect 130068 78344 130074 78356
rect 131114 78344 131120 78356
rect 131172 78344 131178 78396
rect 134058 78344 134064 78396
rect 134116 78384 134122 78396
rect 134610 78384 134616 78396
rect 134116 78356 134616 78384
rect 134116 78344 134122 78356
rect 134610 78344 134616 78356
rect 134668 78344 134674 78396
rect 170030 78344 170036 78396
rect 170088 78384 170094 78396
rect 170398 78384 170404 78396
rect 170088 78356 170404 78384
rect 170088 78344 170094 78356
rect 170398 78344 170404 78356
rect 170456 78344 170462 78396
rect 171318 78344 171324 78396
rect 171376 78384 171382 78396
rect 171594 78384 171600 78396
rect 171376 78356 171600 78384
rect 171376 78344 171382 78356
rect 171594 78344 171600 78356
rect 171652 78344 171658 78396
rect 175734 78344 175740 78396
rect 175792 78384 175798 78396
rect 187602 78384 187608 78396
rect 175792 78356 187608 78384
rect 175792 78344 175798 78356
rect 187602 78344 187608 78356
rect 187660 78344 187666 78396
rect 118666 78288 129596 78316
rect 96614 78208 96620 78260
rect 96672 78248 96678 78260
rect 118666 78248 118694 78288
rect 96672 78220 118694 78248
rect 129568 78248 129596 78288
rect 129642 78276 129648 78328
rect 129700 78316 129706 78328
rect 145742 78316 145748 78328
rect 129700 78288 145748 78316
rect 129700 78276 129706 78288
rect 145742 78276 145748 78288
rect 145800 78276 145806 78328
rect 155770 78276 155776 78328
rect 155828 78316 155834 78328
rect 177482 78316 177488 78328
rect 155828 78288 177488 78316
rect 155828 78276 155834 78288
rect 177482 78276 177488 78288
rect 177540 78276 177546 78328
rect 181364 78288 181576 78316
rect 138106 78248 138112 78260
rect 129568 78220 138112 78248
rect 96672 78208 96678 78220
rect 138106 78208 138112 78220
rect 138164 78208 138170 78260
rect 143902 78208 143908 78260
rect 143960 78248 143966 78260
rect 144086 78248 144092 78260
rect 143960 78220 144092 78248
rect 143960 78208 143966 78220
rect 144086 78208 144092 78220
rect 144144 78208 144150 78260
rect 155310 78208 155316 78260
rect 155368 78248 155374 78260
rect 166902 78248 166908 78260
rect 155368 78220 166908 78248
rect 155368 78208 155374 78220
rect 166902 78208 166908 78220
rect 166960 78208 166966 78260
rect 167086 78208 167092 78260
rect 167144 78248 167150 78260
rect 181364 78248 181392 78288
rect 167144 78220 181392 78248
rect 181548 78248 181576 78288
rect 186130 78248 186136 78260
rect 181548 78220 186136 78248
rect 167144 78208 167150 78220
rect 186130 78208 186136 78220
rect 186188 78208 186194 78260
rect 186406 78208 186412 78260
rect 186464 78248 186470 78260
rect 268378 78248 268384 78260
rect 186464 78220 268384 78248
rect 186464 78208 186470 78220
rect 268378 78208 268384 78220
rect 268436 78208 268442 78260
rect 78674 78140 78680 78192
rect 78732 78180 78738 78192
rect 136726 78180 136732 78192
rect 78732 78152 136732 78180
rect 78732 78140 78738 78152
rect 136726 78140 136732 78152
rect 136784 78140 136790 78192
rect 161750 78140 161756 78192
rect 161808 78180 161814 78192
rect 162026 78180 162032 78192
rect 161808 78152 162032 78180
rect 161808 78140 161814 78152
rect 162026 78140 162032 78152
rect 162084 78140 162090 78192
rect 164326 78140 164332 78192
rect 164384 78180 164390 78192
rect 164602 78180 164608 78192
rect 164384 78152 164608 78180
rect 164384 78140 164390 78152
rect 164602 78140 164608 78152
rect 164660 78140 164666 78192
rect 164878 78140 164884 78192
rect 164936 78180 164942 78192
rect 180150 78180 180156 78192
rect 164936 78152 180156 78180
rect 164936 78140 164942 78152
rect 180150 78140 180156 78152
rect 180208 78140 180214 78192
rect 187602 78140 187608 78192
rect 187660 78180 187666 78192
rect 337378 78180 337384 78192
rect 187660 78152 337384 78180
rect 187660 78140 187666 78152
rect 337378 78140 337384 78152
rect 337436 78140 337442 78192
rect 10318 78072 10324 78124
rect 10376 78112 10382 78124
rect 130930 78112 130936 78124
rect 10376 78084 130936 78112
rect 10376 78072 10382 78084
rect 130930 78072 130936 78084
rect 130988 78072 130994 78124
rect 131114 78072 131120 78124
rect 131172 78112 131178 78124
rect 133966 78112 133972 78124
rect 131172 78084 133972 78112
rect 131172 78072 131178 78084
rect 133966 78072 133972 78084
rect 134024 78072 134030 78124
rect 144270 78112 144276 78124
rect 144196 78084 144276 78112
rect 43438 78004 43444 78056
rect 43496 78044 43502 78056
rect 132126 78044 132132 78056
rect 43496 78016 132132 78044
rect 43496 78004 43502 78016
rect 132126 78004 132132 78016
rect 132184 78004 132190 78056
rect 137002 78004 137008 78056
rect 137060 78044 137066 78056
rect 137370 78044 137376 78056
rect 137060 78016 137376 78044
rect 137060 78004 137066 78016
rect 137370 78004 137376 78016
rect 137428 78004 137434 78056
rect 2774 77936 2780 77988
rect 2832 77976 2838 77988
rect 130838 77976 130844 77988
rect 2832 77948 130844 77976
rect 2832 77936 2838 77948
rect 130838 77936 130844 77948
rect 130896 77936 130902 77988
rect 130930 77936 130936 77988
rect 130988 77976 130994 77988
rect 138566 77976 138572 77988
rect 130988 77948 138572 77976
rect 130988 77936 130994 77948
rect 138566 77936 138572 77948
rect 138624 77936 138630 77988
rect 131206 77732 131212 77784
rect 131264 77772 131270 77784
rect 131574 77772 131580 77784
rect 131264 77744 131580 77772
rect 131264 77732 131270 77744
rect 131574 77732 131580 77744
rect 131632 77732 131638 77784
rect 139394 77732 139400 77784
rect 139452 77772 139458 77784
rect 140590 77772 140596 77784
rect 139452 77744 140596 77772
rect 139452 77732 139458 77744
rect 140590 77732 140596 77744
rect 140648 77732 140654 77784
rect 144196 77772 144224 78084
rect 144270 78072 144276 78084
rect 144328 78072 144334 78124
rect 151354 78072 151360 78124
rect 151412 78112 151418 78124
rect 155310 78112 155316 78124
rect 151412 78084 155316 78112
rect 151412 78072 151418 78084
rect 155310 78072 155316 78084
rect 155368 78072 155374 78124
rect 158806 78072 158812 78124
rect 158864 78112 158870 78124
rect 166902 78112 166908 78124
rect 158864 78084 166908 78112
rect 158864 78072 158870 78084
rect 166902 78072 166908 78084
rect 166960 78072 166966 78124
rect 169018 78072 169024 78124
rect 169076 78112 169082 78124
rect 169662 78112 169668 78124
rect 169076 78084 169668 78112
rect 169076 78072 169082 78084
rect 169662 78072 169668 78084
rect 169720 78072 169726 78124
rect 170214 78072 170220 78124
rect 170272 78112 170278 78124
rect 170674 78112 170680 78124
rect 170272 78084 170680 78112
rect 170272 78072 170278 78084
rect 170674 78072 170680 78084
rect 170732 78072 170738 78124
rect 175918 78072 175924 78124
rect 175976 78112 175982 78124
rect 349798 78112 349804 78124
rect 175976 78084 349804 78112
rect 175976 78072 175982 78084
rect 349798 78072 349804 78084
rect 349856 78072 349862 78124
rect 161198 78004 161204 78056
rect 161256 78044 161262 78056
rect 164878 78044 164884 78056
rect 161256 78016 164884 78044
rect 161256 78004 161262 78016
rect 164878 78004 164884 78016
rect 164936 78004 164942 78056
rect 167546 78004 167552 78056
rect 167604 78044 167610 78056
rect 431218 78044 431224 78056
rect 167604 78016 431224 78044
rect 167604 78004 167610 78016
rect 431218 78004 431224 78016
rect 431276 78004 431282 78056
rect 146478 77936 146484 77988
rect 146536 77976 146542 77988
rect 151354 77976 151360 77988
rect 146536 77948 151360 77976
rect 146536 77936 146542 77948
rect 151354 77936 151360 77948
rect 151412 77936 151418 77988
rect 154942 77936 154948 77988
rect 155000 77976 155006 77988
rect 155000 77948 164234 77976
rect 155000 77936 155006 77948
rect 161658 77868 161664 77920
rect 161716 77908 161722 77920
rect 162394 77908 162400 77920
rect 161716 77880 162400 77908
rect 161716 77868 161722 77880
rect 162394 77868 162400 77880
rect 162452 77868 162458 77920
rect 164206 77908 164234 77948
rect 164602 77936 164608 77988
rect 164660 77976 164666 77988
rect 164970 77976 164976 77988
rect 164660 77948 164976 77976
rect 164660 77936 164666 77948
rect 164970 77936 164976 77948
rect 165028 77936 165034 77988
rect 168742 77936 168748 77988
rect 168800 77976 168806 77988
rect 489914 77976 489920 77988
rect 168800 77948 489920 77976
rect 168800 77936 168806 77948
rect 489914 77936 489920 77948
rect 489972 77936 489978 77988
rect 172606 77908 172612 77920
rect 164206 77880 172612 77908
rect 172606 77868 172612 77880
rect 172664 77868 172670 77920
rect 177390 77908 177396 77920
rect 176626 77880 177396 77908
rect 151630 77800 151636 77852
rect 151688 77840 151694 77852
rect 162118 77840 162124 77852
rect 151688 77812 162124 77840
rect 151688 77800 151694 77812
rect 162118 77800 162124 77812
rect 162176 77800 162182 77852
rect 165798 77800 165804 77852
rect 165856 77840 165862 77852
rect 166442 77840 166448 77852
rect 165856 77812 166448 77840
rect 165856 77800 165862 77812
rect 166442 77800 166448 77812
rect 166500 77800 166506 77852
rect 167362 77800 167368 77852
rect 167420 77840 167426 77852
rect 167546 77840 167552 77852
rect 167420 77812 167552 77840
rect 167420 77800 167426 77812
rect 167546 77800 167552 77812
rect 167604 77800 167610 77852
rect 169938 77800 169944 77852
rect 169996 77840 170002 77852
rect 170122 77840 170128 77852
rect 169996 77812 170128 77840
rect 169996 77800 170002 77812
rect 170122 77800 170128 77812
rect 170180 77800 170186 77852
rect 170582 77800 170588 77852
rect 170640 77840 170646 77852
rect 170858 77840 170864 77852
rect 170640 77812 170864 77840
rect 170640 77800 170646 77812
rect 170858 77800 170864 77812
rect 170916 77800 170922 77852
rect 171042 77800 171048 77852
rect 171100 77840 171106 77852
rect 171686 77840 171692 77852
rect 171100 77812 171692 77840
rect 171100 77800 171106 77812
rect 171686 77800 171692 77812
rect 171744 77800 171750 77852
rect 144362 77772 144368 77784
rect 144196 77744 144368 77772
rect 144362 77732 144368 77744
rect 144420 77732 144426 77784
rect 150802 77732 150808 77784
rect 150860 77772 150866 77784
rect 162394 77772 162400 77784
rect 150860 77744 162400 77772
rect 150860 77732 150866 77744
rect 162394 77732 162400 77744
rect 162452 77732 162458 77784
rect 164234 77732 164240 77784
rect 164292 77772 164298 77784
rect 164292 77744 169110 77772
rect 164292 77732 164298 77744
rect 130562 77664 130568 77716
rect 130620 77704 130626 77716
rect 138382 77704 138388 77716
rect 130620 77676 138388 77704
rect 130620 77664 130626 77676
rect 138382 77664 138388 77676
rect 138440 77664 138446 77716
rect 147858 77664 147864 77716
rect 147916 77704 147922 77716
rect 147916 77676 162164 77704
rect 147916 77664 147922 77676
rect 129182 77596 129188 77648
rect 129240 77636 129246 77648
rect 139670 77636 139676 77648
rect 129240 77608 139676 77636
rect 129240 77596 129246 77608
rect 139670 77596 139676 77608
rect 139728 77596 139734 77648
rect 145282 77596 145288 77648
rect 145340 77636 145346 77648
rect 145340 77608 153194 77636
rect 145340 77596 145346 77608
rect 134518 77528 134524 77580
rect 134576 77568 134582 77580
rect 136358 77568 136364 77580
rect 134576 77540 136364 77568
rect 134576 77528 134582 77540
rect 136358 77528 136364 77540
rect 136416 77528 136422 77580
rect 153166 77568 153194 77608
rect 159818 77596 159824 77648
rect 159876 77636 159882 77648
rect 162136 77636 162164 77676
rect 165798 77664 165804 77716
rect 165856 77704 165862 77716
rect 165982 77704 165988 77716
rect 165856 77676 165988 77704
rect 165856 77664 165862 77676
rect 165982 77664 165988 77676
rect 166040 77664 166046 77716
rect 169082 77704 169110 77744
rect 169662 77732 169668 77784
rect 169720 77772 169726 77784
rect 176626 77772 176654 77880
rect 177390 77868 177396 77880
rect 177448 77868 177454 77920
rect 176838 77800 176844 77852
rect 176896 77840 176902 77852
rect 580350 77840 580356 77852
rect 176896 77812 580356 77840
rect 176896 77800 176902 77812
rect 580350 77800 580356 77812
rect 580408 77800 580414 77852
rect 169720 77744 176654 77772
rect 169720 77732 169726 77744
rect 177298 77732 177304 77784
rect 177356 77772 177362 77784
rect 191098 77772 191104 77784
rect 177356 77744 191104 77772
rect 177356 77732 177362 77744
rect 191098 77732 191104 77744
rect 191156 77732 191162 77784
rect 177206 77704 177212 77716
rect 169082 77676 177212 77704
rect 177206 77664 177212 77676
rect 177264 77664 177270 77716
rect 168282 77636 168288 77648
rect 159876 77608 162072 77636
rect 162136 77608 168288 77636
rect 159876 77596 159882 77608
rect 161106 77568 161112 77580
rect 153166 77540 161112 77568
rect 161106 77528 161112 77540
rect 161164 77528 161170 77580
rect 162044 77568 162072 77608
rect 168282 77596 168288 77608
rect 168340 77596 168346 77648
rect 169754 77596 169760 77648
rect 169812 77636 169818 77648
rect 177298 77636 177304 77648
rect 169812 77608 177304 77636
rect 169812 77596 169818 77608
rect 177298 77596 177304 77608
rect 177356 77596 177362 77648
rect 167730 77568 167736 77580
rect 162044 77540 167736 77568
rect 167730 77528 167736 77540
rect 167788 77528 167794 77580
rect 168006 77528 168012 77580
rect 168064 77568 168070 77580
rect 176286 77568 176292 77580
rect 168064 77540 176292 77568
rect 168064 77528 168070 77540
rect 176286 77528 176292 77540
rect 176344 77528 176350 77580
rect 158438 77460 158444 77512
rect 158496 77500 158502 77512
rect 165430 77500 165436 77512
rect 158496 77472 165436 77500
rect 158496 77460 158502 77472
rect 165430 77460 165436 77472
rect 165488 77460 165494 77512
rect 166350 77460 166356 77512
rect 166408 77500 166414 77512
rect 181438 77500 181444 77512
rect 166408 77472 181444 77500
rect 166408 77460 166414 77472
rect 181438 77460 181444 77472
rect 181496 77460 181502 77512
rect 130470 77392 130476 77444
rect 130528 77432 130534 77444
rect 137830 77432 137836 77444
rect 130528 77404 137836 77432
rect 130528 77392 130534 77404
rect 137830 77392 137836 77404
rect 137888 77392 137894 77444
rect 155218 77392 155224 77444
rect 155276 77432 155282 77444
rect 155770 77432 155776 77444
rect 155276 77404 155776 77432
rect 155276 77392 155282 77404
rect 155770 77392 155776 77404
rect 155828 77392 155834 77444
rect 158714 77392 158720 77444
rect 158772 77432 158778 77444
rect 159634 77432 159640 77444
rect 158772 77404 159640 77432
rect 158772 77392 158778 77404
rect 159634 77392 159640 77404
rect 159692 77392 159698 77444
rect 160278 77392 160284 77444
rect 160336 77432 160342 77444
rect 168006 77432 168012 77444
rect 160336 77404 168012 77432
rect 160336 77392 160342 77404
rect 168006 77392 168012 77404
rect 168064 77392 168070 77444
rect 177666 77392 177672 77444
rect 177724 77432 177730 77444
rect 177850 77432 177856 77444
rect 177724 77404 177856 77432
rect 177724 77392 177730 77404
rect 177850 77392 177856 77404
rect 177908 77392 177914 77444
rect 178126 77392 178132 77444
rect 178184 77432 178190 77444
rect 179414 77432 179420 77444
rect 178184 77404 179420 77432
rect 178184 77392 178190 77404
rect 179414 77392 179420 77404
rect 179472 77392 179478 77444
rect 130194 77324 130200 77376
rect 130252 77364 130258 77376
rect 137646 77364 137652 77376
rect 130252 77336 137652 77364
rect 130252 77324 130258 77336
rect 137646 77324 137652 77336
rect 137704 77324 137710 77376
rect 164234 77324 164240 77376
rect 164292 77364 164298 77376
rect 165154 77364 165160 77376
rect 164292 77336 165160 77364
rect 164292 77324 164298 77336
rect 165154 77324 165160 77336
rect 165212 77324 165218 77376
rect 165614 77324 165620 77376
rect 165672 77364 165678 77376
rect 175826 77364 175832 77376
rect 165672 77336 175832 77364
rect 165672 77324 165678 77336
rect 175826 77324 175832 77336
rect 175884 77324 175890 77376
rect 131758 77256 131764 77308
rect 131816 77296 131822 77308
rect 135806 77296 135812 77308
rect 131816 77268 135812 77296
rect 131816 77256 131822 77268
rect 135806 77256 135812 77268
rect 135864 77256 135870 77308
rect 145374 77256 145380 77308
rect 145432 77296 145438 77308
rect 147214 77296 147220 77308
rect 145432 77268 147220 77296
rect 145432 77256 145438 77268
rect 147214 77256 147220 77268
rect 147272 77256 147278 77308
rect 151906 77256 151912 77308
rect 151964 77296 151970 77308
rect 152918 77296 152924 77308
rect 151964 77268 152924 77296
rect 151964 77256 151970 77268
rect 152918 77256 152924 77268
rect 152976 77256 152982 77308
rect 153378 77256 153384 77308
rect 153436 77296 153442 77308
rect 154114 77296 154120 77308
rect 153436 77268 154120 77296
rect 153436 77256 153442 77268
rect 154114 77256 154120 77268
rect 154172 77256 154178 77308
rect 154574 77256 154580 77308
rect 154632 77296 154638 77308
rect 154942 77296 154948 77308
rect 154632 77268 154948 77296
rect 154632 77256 154638 77268
rect 154942 77256 154948 77268
rect 155000 77256 155006 77308
rect 158898 77256 158904 77308
rect 158956 77296 158962 77308
rect 159082 77296 159088 77308
rect 158956 77268 159088 77296
rect 158956 77256 158962 77268
rect 159082 77256 159088 77268
rect 159140 77256 159146 77308
rect 173066 77256 173072 77308
rect 173124 77296 173130 77308
rect 176378 77296 176384 77308
rect 173124 77268 176384 77296
rect 173124 77256 173130 77268
rect 176378 77256 176384 77268
rect 176436 77256 176442 77308
rect 176746 77256 176752 77308
rect 176804 77296 176810 77308
rect 177850 77296 177856 77308
rect 176804 77268 177856 77296
rect 176804 77256 176810 77268
rect 177850 77256 177856 77268
rect 177908 77256 177914 77308
rect 150434 77188 150440 77240
rect 150492 77228 150498 77240
rect 151078 77228 151084 77240
rect 150492 77200 151084 77228
rect 150492 77188 150498 77200
rect 151078 77188 151084 77200
rect 151136 77188 151142 77240
rect 153194 77188 153200 77240
rect 153252 77228 153258 77240
rect 153746 77228 153752 77240
rect 153252 77200 153752 77228
rect 153252 77188 153258 77200
rect 153746 77188 153752 77200
rect 153804 77188 153810 77240
rect 154758 77188 154764 77240
rect 154816 77228 154822 77240
rect 158622 77228 158628 77240
rect 154816 77200 158628 77228
rect 154816 77188 154822 77200
rect 158622 77188 158628 77200
rect 158680 77188 158686 77240
rect 160370 77188 160376 77240
rect 160428 77228 160434 77240
rect 160830 77228 160836 77240
rect 160428 77200 160836 77228
rect 160428 77188 160434 77200
rect 160830 77188 160836 77200
rect 160888 77188 160894 77240
rect 161106 77188 161112 77240
rect 161164 77228 161170 77240
rect 186314 77228 186320 77240
rect 161164 77200 186320 77228
rect 161164 77188 161170 77200
rect 186314 77188 186320 77200
rect 186372 77188 186378 77240
rect 145926 77120 145932 77172
rect 145984 77160 145990 77172
rect 171870 77160 171876 77172
rect 145984 77132 171876 77160
rect 145984 77120 145990 77132
rect 171870 77120 171876 77132
rect 171928 77120 171934 77172
rect 140590 77052 140596 77104
rect 140648 77092 140654 77104
rect 141050 77092 141056 77104
rect 140648 77064 141056 77092
rect 140648 77052 140654 77064
rect 141050 77052 141056 77064
rect 141108 77052 141114 77104
rect 240134 77092 240140 77104
rect 157306 77064 240140 77092
rect 132586 76984 132592 77036
rect 132644 77024 132650 77036
rect 132954 77024 132960 77036
rect 132644 76996 132960 77024
rect 132644 76984 132650 76996
rect 132954 76984 132960 76996
rect 133012 76984 133018 77036
rect 156690 76984 156696 77036
rect 156748 77024 156754 77036
rect 157306 77024 157334 77064
rect 240134 77052 240140 77064
rect 240192 77052 240198 77104
rect 156748 76996 157334 77024
rect 156748 76984 156754 76996
rect 157518 76984 157524 77036
rect 157576 77024 157582 77036
rect 158070 77024 158076 77036
rect 157576 76996 158076 77024
rect 157576 76984 157582 76996
rect 158070 76984 158076 76996
rect 158128 76984 158134 77036
rect 171134 76984 171140 77036
rect 171192 77024 171198 77036
rect 260834 77024 260840 77036
rect 171192 76996 260840 77024
rect 171192 76984 171198 76996
rect 260834 76984 260840 76996
rect 260892 76984 260898 77036
rect 151446 76916 151452 76968
rect 151504 76956 151510 76968
rect 267734 76956 267740 76968
rect 151504 76928 267740 76956
rect 151504 76916 151510 76928
rect 267734 76916 267740 76928
rect 267792 76916 267798 76968
rect 126974 76848 126980 76900
rect 127032 76888 127038 76900
rect 140498 76888 140504 76900
rect 127032 76860 140504 76888
rect 127032 76848 127038 76860
rect 140498 76848 140504 76860
rect 140556 76848 140562 76900
rect 142706 76848 142712 76900
rect 142764 76888 142770 76900
rect 143074 76888 143080 76900
rect 142764 76860 143080 76888
rect 142764 76848 142770 76860
rect 143074 76848 143080 76860
rect 143132 76848 143138 76900
rect 150526 76848 150532 76900
rect 150584 76888 150590 76900
rect 150710 76888 150716 76900
rect 150584 76860 150716 76888
rect 150584 76848 150590 76860
rect 150710 76848 150716 76860
rect 150768 76848 150774 76900
rect 157426 76848 157432 76900
rect 157484 76888 157490 76900
rect 158254 76888 158260 76900
rect 157484 76860 158260 76888
rect 157484 76848 157490 76860
rect 158254 76848 158260 76860
rect 158312 76848 158318 76900
rect 165614 76848 165620 76900
rect 165672 76888 165678 76900
rect 166166 76888 166172 76900
rect 165672 76860 166172 76888
rect 165672 76848 165678 76860
rect 166166 76848 166172 76860
rect 166224 76848 166230 76900
rect 171042 76848 171048 76900
rect 171100 76888 171106 76900
rect 327074 76888 327080 76900
rect 171100 76860 327080 76888
rect 171100 76848 171106 76860
rect 327074 76848 327080 76860
rect 327132 76848 327138 76900
rect 91094 76780 91100 76832
rect 91152 76820 91158 76832
rect 137738 76820 137744 76832
rect 91152 76792 137744 76820
rect 91152 76780 91158 76792
rect 137738 76780 137744 76792
rect 137796 76780 137802 76832
rect 142062 76780 142068 76832
rect 142120 76820 142126 76832
rect 142522 76820 142528 76832
rect 142120 76792 142528 76820
rect 142120 76780 142126 76792
rect 142522 76780 142528 76792
rect 142580 76780 142586 76832
rect 156874 76780 156880 76832
rect 156932 76820 156938 76832
rect 328454 76820 328460 76832
rect 156932 76792 328460 76820
rect 156932 76780 156938 76792
rect 328454 76780 328460 76792
rect 328512 76780 328518 76832
rect 104894 76712 104900 76764
rect 104952 76752 104958 76764
rect 138290 76752 138296 76764
rect 104952 76724 138296 76752
rect 104952 76712 104958 76724
rect 138290 76712 138296 76724
rect 138348 76712 138354 76764
rect 142430 76712 142436 76764
rect 142488 76752 142494 76764
rect 143074 76752 143080 76764
rect 142488 76724 143080 76752
rect 142488 76712 142494 76724
rect 143074 76712 143080 76724
rect 143132 76712 143138 76764
rect 147858 76712 147864 76764
rect 147916 76752 147922 76764
rect 148410 76752 148416 76764
rect 147916 76724 148416 76752
rect 147916 76712 147922 76724
rect 148410 76712 148416 76724
rect 148468 76712 148474 76764
rect 157426 76712 157432 76764
rect 157484 76752 157490 76764
rect 158162 76752 158168 76764
rect 157484 76724 158168 76752
rect 157484 76712 157490 76724
rect 158162 76712 158168 76724
rect 158220 76712 158226 76764
rect 160094 76712 160100 76764
rect 160152 76752 160158 76764
rect 160370 76752 160376 76764
rect 160152 76724 160376 76752
rect 160152 76712 160158 76724
rect 160370 76712 160376 76724
rect 160428 76712 160434 76764
rect 160738 76712 160744 76764
rect 160796 76712 160802 76764
rect 161290 76712 161296 76764
rect 161348 76752 161354 76764
rect 161348 76724 171364 76752
rect 161348 76712 161354 76724
rect 84194 76644 84200 76696
rect 84252 76684 84258 76696
rect 135254 76684 135260 76696
rect 84252 76656 135260 76684
rect 84252 76644 84258 76656
rect 135254 76644 135260 76656
rect 135312 76644 135318 76696
rect 159174 76644 159180 76696
rect 159232 76684 159238 76696
rect 159726 76684 159732 76696
rect 159232 76656 159732 76684
rect 159232 76644 159238 76656
rect 159726 76644 159732 76656
rect 159784 76644 159790 76696
rect 160756 76684 160784 76712
rect 160388 76656 160784 76684
rect 41414 76576 41420 76628
rect 41472 76616 41478 76628
rect 133506 76616 133512 76628
rect 41472 76588 133512 76616
rect 41472 76576 41478 76588
rect 133506 76576 133512 76588
rect 133564 76576 133570 76628
rect 154758 76576 154764 76628
rect 154816 76616 154822 76628
rect 155586 76616 155592 76628
rect 154816 76588 155592 76616
rect 154816 76576 154822 76588
rect 155586 76576 155592 76588
rect 155644 76576 155650 76628
rect 155954 76576 155960 76628
rect 156012 76616 156018 76628
rect 156414 76616 156420 76628
rect 156012 76588 156420 76616
rect 156012 76576 156018 76588
rect 156414 76576 156420 76588
rect 156472 76576 156478 76628
rect 158806 76576 158812 76628
rect 158864 76616 158870 76628
rect 159358 76616 159364 76628
rect 158864 76588 159364 76616
rect 158864 76576 158870 76588
rect 159358 76576 159364 76588
rect 159416 76576 159422 76628
rect 34514 76508 34520 76560
rect 34572 76548 34578 76560
rect 133046 76548 133052 76560
rect 34572 76520 133052 76548
rect 34572 76508 34578 76520
rect 133046 76508 133052 76520
rect 133104 76508 133110 76560
rect 158898 76508 158904 76560
rect 158956 76548 158962 76560
rect 159450 76548 159456 76560
rect 158956 76520 159456 76548
rect 158956 76508 158962 76520
rect 159450 76508 159456 76520
rect 159508 76508 159514 76560
rect 160388 76492 160416 76656
rect 165338 76644 165344 76696
rect 165396 76684 165402 76696
rect 165890 76684 165896 76696
rect 165396 76656 165896 76684
rect 165396 76644 165402 76656
rect 165890 76644 165896 76656
rect 165948 76644 165954 76696
rect 171336 76684 171364 76724
rect 172054 76712 172060 76764
rect 172112 76752 172118 76764
rect 368474 76752 368480 76764
rect 172112 76724 368480 76752
rect 172112 76712 172118 76724
rect 368474 76712 368480 76724
rect 368532 76712 368538 76764
rect 367094 76684 367100 76696
rect 171336 76656 367100 76684
rect 367094 76644 367100 76656
rect 367152 76644 367158 76696
rect 160738 76576 160744 76628
rect 160796 76616 160802 76628
rect 161014 76616 161020 76628
rect 160796 76588 161020 76616
rect 160796 76576 160802 76588
rect 161014 76576 161020 76588
rect 161072 76576 161078 76628
rect 161566 76576 161572 76628
rect 161624 76616 161630 76628
rect 161934 76616 161940 76628
rect 161624 76588 161940 76616
rect 161624 76576 161630 76588
rect 161934 76576 161940 76588
rect 161992 76576 161998 76628
rect 162118 76576 162124 76628
rect 162176 76616 162182 76628
rect 171134 76616 171140 76628
rect 162176 76588 171140 76616
rect 162176 76576 162182 76588
rect 171134 76576 171140 76588
rect 171192 76576 171198 76628
rect 485774 76616 485780 76628
rect 176626 76588 485780 76616
rect 160462 76508 160468 76560
rect 160520 76548 160526 76560
rect 160922 76548 160928 76560
rect 160520 76520 160928 76548
rect 160520 76508 160526 76520
rect 160922 76508 160928 76520
rect 160980 76508 160986 76560
rect 166166 76508 166172 76560
rect 166224 76548 166230 76560
rect 166534 76548 166540 76560
rect 166224 76520 166540 76548
rect 166224 76508 166230 76520
rect 166534 76508 166540 76520
rect 166592 76508 166598 76560
rect 168374 76508 168380 76560
rect 168432 76548 168438 76560
rect 176626 76548 176654 76588
rect 485774 76576 485780 76588
rect 485832 76576 485838 76628
rect 542354 76548 542360 76560
rect 168432 76520 176654 76548
rect 186286 76520 542360 76548
rect 168432 76508 168438 76520
rect 147950 76440 147956 76492
rect 148008 76480 148014 76492
rect 148134 76480 148140 76492
rect 148008 76452 148140 76480
rect 148008 76440 148014 76452
rect 148134 76440 148140 76452
rect 148192 76440 148198 76492
rect 149330 76440 149336 76492
rect 149388 76480 149394 76492
rect 149790 76480 149796 76492
rect 149388 76452 149796 76480
rect 149388 76440 149394 76452
rect 149790 76440 149796 76452
rect 149848 76440 149854 76492
rect 158990 76440 158996 76492
rect 159048 76480 159054 76492
rect 159542 76480 159548 76492
rect 159048 76452 159548 76480
rect 159048 76440 159054 76452
rect 159542 76440 159548 76452
rect 159600 76440 159606 76492
rect 160370 76440 160376 76492
rect 160428 76440 160434 76492
rect 160646 76440 160652 76492
rect 160704 76480 160710 76492
rect 161198 76480 161204 76492
rect 160704 76452 161204 76480
rect 160704 76440 160710 76452
rect 161198 76440 161204 76452
rect 161256 76440 161262 76492
rect 161934 76440 161940 76492
rect 161992 76480 161998 76492
rect 162302 76480 162308 76492
rect 161992 76452 162308 76480
rect 161992 76440 161998 76452
rect 162302 76440 162308 76452
rect 162360 76440 162366 76492
rect 171870 76440 171876 76492
rect 171928 76480 171934 76492
rect 178678 76480 178684 76492
rect 171928 76452 178684 76480
rect 171928 76440 171934 76452
rect 178678 76440 178684 76452
rect 178736 76440 178742 76492
rect 152274 76372 152280 76424
rect 152332 76412 152338 76424
rect 152550 76412 152556 76424
rect 152332 76384 152556 76412
rect 152332 76372 152338 76384
rect 152550 76372 152556 76384
rect 152608 76372 152614 76424
rect 162210 76372 162216 76424
rect 162268 76412 162274 76424
rect 172054 76412 172060 76424
rect 162268 76384 172060 76412
rect 162268 76372 162274 76384
rect 172054 76372 172060 76384
rect 172112 76372 172118 76424
rect 173158 76372 173164 76424
rect 173216 76412 173222 76424
rect 186286 76412 186314 76520
rect 542354 76508 542360 76520
rect 542412 76508 542418 76560
rect 173216 76384 186314 76412
rect 173216 76372 173222 76384
rect 147950 76304 147956 76356
rect 148008 76344 148014 76356
rect 148502 76344 148508 76356
rect 148008 76316 148508 76344
rect 148008 76304 148014 76316
rect 148502 76304 148508 76316
rect 148560 76304 148566 76356
rect 154574 76304 154580 76356
rect 154632 76344 154638 76356
rect 155494 76344 155500 76356
rect 154632 76316 155500 76344
rect 154632 76304 154638 76316
rect 155494 76304 155500 76316
rect 155552 76304 155558 76356
rect 168374 76304 168380 76356
rect 168432 76344 168438 76356
rect 168834 76344 168840 76356
rect 168432 76316 168840 76344
rect 168432 76304 168438 76316
rect 168834 76304 168840 76316
rect 168892 76304 168898 76356
rect 149146 76236 149152 76288
rect 149204 76276 149210 76288
rect 149698 76276 149704 76288
rect 149204 76248 149704 76276
rect 149204 76236 149210 76248
rect 149698 76236 149704 76248
rect 149756 76236 149762 76288
rect 144454 76168 144460 76220
rect 144512 76208 144518 76220
rect 145742 76208 145748 76220
rect 144512 76180 145748 76208
rect 144512 76168 144518 76180
rect 145742 76168 145748 76180
rect 145800 76168 145806 76220
rect 163314 76168 163320 76220
rect 163372 76208 163378 76220
rect 163498 76208 163504 76220
rect 163372 76180 163504 76208
rect 163372 76168 163378 76180
rect 163498 76168 163504 76180
rect 163556 76168 163562 76220
rect 139762 76100 139768 76152
rect 139820 76140 139826 76152
rect 139946 76140 139952 76152
rect 139820 76112 139952 76140
rect 139820 76100 139826 76112
rect 139946 76100 139952 76112
rect 140004 76100 140010 76152
rect 149146 76100 149152 76152
rect 149204 76140 149210 76152
rect 149422 76140 149428 76152
rect 149204 76112 149428 76140
rect 149204 76100 149210 76112
rect 149422 76100 149428 76112
rect 149480 76100 149486 76152
rect 168650 76100 168656 76152
rect 168708 76140 168714 76152
rect 169110 76140 169116 76152
rect 168708 76112 169116 76140
rect 168708 76100 168714 76112
rect 169110 76100 169116 76112
rect 169168 76100 169174 76152
rect 139946 75964 139952 76016
rect 140004 76004 140010 76016
rect 140222 76004 140228 76016
rect 140004 75976 140228 76004
rect 140004 75964 140010 75976
rect 140222 75964 140228 75976
rect 140280 75964 140286 76016
rect 143626 75964 143632 76016
rect 143684 76004 143690 76016
rect 144454 76004 144460 76016
rect 143684 75976 144460 76004
rect 143684 75964 143690 75976
rect 144454 75964 144460 75976
rect 144512 75964 144518 76016
rect 142522 75896 142528 75948
rect 142580 75936 142586 75948
rect 142798 75936 142804 75948
rect 142580 75908 142804 75936
rect 142580 75896 142586 75908
rect 142798 75896 142804 75908
rect 142856 75896 142862 75948
rect 150710 75896 150716 75948
rect 150768 75936 150774 75948
rect 151078 75936 151084 75948
rect 150768 75908 151084 75936
rect 150768 75896 150774 75908
rect 151078 75896 151084 75908
rect 151136 75896 151142 75948
rect 140222 75828 140228 75880
rect 140280 75868 140286 75880
rect 141234 75868 141240 75880
rect 140280 75840 141240 75868
rect 140280 75828 140286 75840
rect 141234 75828 141240 75840
rect 141292 75828 141298 75880
rect 150802 75828 150808 75880
rect 150860 75868 150866 75880
rect 151170 75868 151176 75880
rect 150860 75840 151176 75868
rect 150860 75828 150866 75840
rect 151170 75828 151176 75840
rect 151228 75828 151234 75880
rect 152182 75828 152188 75880
rect 152240 75868 152246 75880
rect 152642 75868 152648 75880
rect 152240 75840 152648 75868
rect 152240 75828 152246 75840
rect 152642 75828 152648 75840
rect 152700 75828 152706 75880
rect 151998 75760 152004 75812
rect 152056 75800 152062 75812
rect 152274 75800 152280 75812
rect 152056 75772 152280 75800
rect 152056 75760 152062 75772
rect 152274 75760 152280 75772
rect 152332 75760 152338 75812
rect 169570 75760 169576 75812
rect 169628 75800 169634 75812
rect 175090 75800 175096 75812
rect 169628 75772 175096 75800
rect 169628 75760 169634 75772
rect 175090 75760 175096 75772
rect 175148 75760 175154 75812
rect 131022 75692 131028 75744
rect 131080 75732 131086 75744
rect 137462 75732 137468 75744
rect 131080 75704 137468 75732
rect 131080 75692 131086 75704
rect 137462 75692 137468 75704
rect 137520 75692 137526 75744
rect 141234 75692 141240 75744
rect 141292 75732 141298 75744
rect 141602 75732 141608 75744
rect 141292 75704 141608 75732
rect 141292 75692 141298 75704
rect 141602 75692 141608 75704
rect 141660 75692 141666 75744
rect 170674 75692 170680 75744
rect 170732 75732 170738 75744
rect 174998 75732 175004 75744
rect 170732 75704 175004 75732
rect 170732 75692 170738 75704
rect 174998 75692 175004 75704
rect 175056 75692 175062 75744
rect 130102 75624 130108 75676
rect 130160 75664 130166 75676
rect 140774 75664 140780 75676
rect 130160 75636 140780 75664
rect 130160 75624 130166 75636
rect 140774 75624 140780 75636
rect 140832 75624 140838 75676
rect 148318 75624 148324 75676
rect 148376 75664 148382 75676
rect 176746 75664 176752 75676
rect 148376 75636 176752 75664
rect 148376 75624 148382 75636
rect 176746 75624 176752 75636
rect 176804 75624 176810 75676
rect 128354 75556 128360 75608
rect 128412 75596 128418 75608
rect 140682 75596 140688 75608
rect 128412 75568 140688 75596
rect 128412 75556 128418 75568
rect 140682 75556 140688 75568
rect 140740 75556 140746 75608
rect 145650 75556 145656 75608
rect 145708 75596 145714 75608
rect 191834 75596 191840 75608
rect 145708 75568 191840 75596
rect 145708 75556 145714 75568
rect 191834 75556 191840 75568
rect 191892 75556 191898 75608
rect 127066 75488 127072 75540
rect 127124 75528 127130 75540
rect 140406 75528 140412 75540
rect 127124 75500 140412 75528
rect 127124 75488 127130 75500
rect 140406 75488 140412 75500
rect 140464 75488 140470 75540
rect 147490 75488 147496 75540
rect 147548 75528 147554 75540
rect 201494 75528 201500 75540
rect 147548 75500 201500 75528
rect 147548 75488 147554 75500
rect 201494 75488 201500 75500
rect 201552 75488 201558 75540
rect 81434 75420 81440 75472
rect 81492 75460 81498 75472
rect 131022 75460 131028 75472
rect 81492 75432 131028 75460
rect 81492 75420 81498 75432
rect 131022 75420 131028 75432
rect 131080 75420 131086 75472
rect 135990 75460 135996 75472
rect 131224 75432 135996 75460
rect 69014 75352 69020 75404
rect 69072 75392 69078 75404
rect 131224 75392 131252 75432
rect 135990 75420 135996 75432
rect 136048 75420 136054 75472
rect 153194 75420 153200 75472
rect 153252 75460 153258 75472
rect 154022 75460 154028 75472
rect 153252 75432 154028 75460
rect 153252 75420 153258 75432
rect 154022 75420 154028 75432
rect 154080 75420 154086 75472
rect 170490 75420 170496 75472
rect 170548 75460 170554 75472
rect 170548 75432 174952 75460
rect 170548 75420 170554 75432
rect 134610 75392 134616 75404
rect 69072 75364 131252 75392
rect 131316 75364 134616 75392
rect 69072 75352 69078 75364
rect 51074 75284 51080 75336
rect 51132 75324 51138 75336
rect 131316 75324 131344 75364
rect 134610 75352 134616 75364
rect 134668 75352 134674 75404
rect 139670 75352 139676 75404
rect 139728 75392 139734 75404
rect 140038 75392 140044 75404
rect 139728 75364 140044 75392
rect 139728 75352 139734 75364
rect 140038 75352 140044 75364
rect 140096 75352 140102 75404
rect 142338 75352 142344 75404
rect 142396 75392 142402 75404
rect 142614 75392 142620 75404
rect 142396 75364 142620 75392
rect 142396 75352 142402 75364
rect 142614 75352 142620 75364
rect 142672 75352 142678 75404
rect 164418 75352 164424 75404
rect 164476 75392 164482 75404
rect 164878 75392 164884 75404
rect 164476 75364 164884 75392
rect 164476 75352 164482 75364
rect 164878 75352 164884 75364
rect 164936 75352 164942 75404
rect 171502 75352 171508 75404
rect 171560 75392 171566 75404
rect 171560 75364 174860 75392
rect 171560 75352 171566 75364
rect 51132 75296 131344 75324
rect 51132 75284 51138 75296
rect 131390 75284 131396 75336
rect 131448 75324 131454 75336
rect 132218 75324 132224 75336
rect 131448 75296 132224 75324
rect 131448 75284 131454 75296
rect 132218 75284 132224 75296
rect 132276 75284 132282 75336
rect 132678 75284 132684 75336
rect 132736 75324 132742 75336
rect 133782 75324 133788 75336
rect 132736 75296 133788 75324
rect 132736 75284 132742 75296
rect 133782 75284 133788 75296
rect 133840 75284 133846 75336
rect 138566 75284 138572 75336
rect 138624 75324 138630 75336
rect 139302 75324 139308 75336
rect 138624 75296 139308 75324
rect 138624 75284 138630 75296
rect 139302 75284 139308 75296
rect 139360 75284 139366 75336
rect 162946 75284 162952 75336
rect 163004 75324 163010 75336
rect 164142 75324 164148 75336
rect 163004 75296 164148 75324
rect 163004 75284 163010 75296
rect 164142 75284 164148 75296
rect 164200 75284 164206 75336
rect 167178 75284 167184 75336
rect 167236 75324 167242 75336
rect 167914 75324 167920 75336
rect 167236 75296 167920 75324
rect 167236 75284 167242 75296
rect 167914 75284 167920 75296
rect 167972 75284 167978 75336
rect 168742 75284 168748 75336
rect 168800 75324 168806 75336
rect 169478 75324 169484 75336
rect 168800 75296 169484 75324
rect 168800 75284 168806 75296
rect 169478 75284 169484 75296
rect 169536 75284 169542 75336
rect 46934 75216 46940 75268
rect 46992 75256 46998 75268
rect 131114 75256 131120 75268
rect 46992 75228 131120 75256
rect 46992 75216 46998 75228
rect 131114 75216 131120 75228
rect 131172 75216 131178 75268
rect 131574 75216 131580 75268
rect 131632 75256 131638 75268
rect 132402 75256 132408 75268
rect 131632 75228 132408 75256
rect 131632 75216 131638 75228
rect 132402 75216 132408 75228
rect 132460 75216 132466 75268
rect 133046 75216 133052 75268
rect 133104 75256 133110 75268
rect 133598 75256 133604 75268
rect 133104 75228 133604 75256
rect 133104 75216 133110 75228
rect 133598 75216 133604 75228
rect 133656 75216 133662 75268
rect 133874 75216 133880 75268
rect 133932 75256 133938 75268
rect 134150 75256 134156 75268
rect 133932 75228 134156 75256
rect 133932 75216 133938 75228
rect 134150 75216 134156 75228
rect 134208 75216 134214 75268
rect 134242 75216 134248 75268
rect 134300 75256 134306 75268
rect 134794 75256 134800 75268
rect 134300 75228 134800 75256
rect 134300 75216 134306 75228
rect 134794 75216 134800 75228
rect 134852 75216 134858 75268
rect 135990 75216 135996 75268
rect 136048 75256 136054 75268
rect 136450 75256 136456 75268
rect 136048 75228 136456 75256
rect 136048 75216 136054 75228
rect 136450 75216 136456 75228
rect 136508 75216 136514 75268
rect 138290 75216 138296 75268
rect 138348 75256 138354 75268
rect 139210 75256 139216 75268
rect 138348 75228 139216 75256
rect 138348 75216 138354 75228
rect 139210 75216 139216 75228
rect 139268 75216 139274 75268
rect 140038 75216 140044 75268
rect 140096 75256 140102 75268
rect 140866 75256 140872 75268
rect 140096 75228 140872 75256
rect 140096 75216 140102 75228
rect 140866 75216 140872 75228
rect 140924 75216 140930 75268
rect 141326 75216 141332 75268
rect 141384 75256 141390 75268
rect 141786 75256 141792 75268
rect 141384 75228 141792 75256
rect 141384 75216 141390 75228
rect 141786 75216 141792 75228
rect 141844 75216 141850 75268
rect 141878 75216 141884 75268
rect 141936 75256 141942 75268
rect 142338 75256 142344 75268
rect 141936 75228 142344 75256
rect 141936 75216 141942 75228
rect 142338 75216 142344 75228
rect 142396 75216 142402 75268
rect 145282 75216 145288 75268
rect 145340 75256 145346 75268
rect 146018 75256 146024 75268
rect 145340 75228 146024 75256
rect 145340 75216 145346 75228
rect 146018 75216 146024 75228
rect 146076 75216 146082 75268
rect 146754 75216 146760 75268
rect 146812 75256 146818 75268
rect 146938 75256 146944 75268
rect 146812 75228 146944 75256
rect 146812 75216 146818 75228
rect 146938 75216 146944 75228
rect 146996 75216 147002 75268
rect 164418 75216 164424 75268
rect 164476 75256 164482 75268
rect 165062 75256 165068 75268
rect 164476 75228 165068 75256
rect 164476 75216 164482 75228
rect 165062 75216 165068 75228
rect 165120 75216 165126 75268
rect 168834 75216 168840 75268
rect 168892 75256 168898 75268
rect 169202 75256 169208 75268
rect 168892 75228 169208 75256
rect 168892 75216 168898 75228
rect 169202 75216 169208 75228
rect 169260 75216 169266 75268
rect 170306 75216 170312 75268
rect 170364 75256 170370 75268
rect 170766 75256 170772 75268
rect 170364 75228 170772 75256
rect 170364 75216 170370 75228
rect 170766 75216 170772 75228
rect 170824 75216 170830 75268
rect 171502 75216 171508 75268
rect 171560 75256 171566 75268
rect 171962 75256 171968 75268
rect 171560 75228 171968 75256
rect 171560 75216 171566 75228
rect 171962 75216 171968 75228
rect 172020 75216 172026 75268
rect 172606 75216 172612 75268
rect 172664 75256 172670 75268
rect 173066 75256 173072 75268
rect 172664 75228 173072 75256
rect 172664 75216 172670 75228
rect 173066 75216 173072 75228
rect 173124 75216 173130 75268
rect 174354 75216 174360 75268
rect 174412 75256 174418 75268
rect 174722 75256 174728 75268
rect 174412 75228 174728 75256
rect 174412 75216 174418 75228
rect 174722 75216 174728 75228
rect 174780 75216 174786 75268
rect 174832 75256 174860 75364
rect 174924 75324 174952 75432
rect 175090 75420 175096 75472
rect 175148 75460 175154 75472
rect 499574 75460 499580 75472
rect 175148 75432 499580 75460
rect 175148 75420 175154 75432
rect 499574 75420 499580 75432
rect 499632 75420 499638 75472
rect 174998 75352 175004 75404
rect 175056 75392 175062 75404
rect 506474 75392 506480 75404
rect 175056 75364 506480 75392
rect 175056 75352 175062 75364
rect 506474 75352 506480 75364
rect 506532 75352 506538 75404
rect 514754 75324 514760 75336
rect 174924 75296 514760 75324
rect 514754 75284 514760 75296
rect 514812 75284 514818 75336
rect 521654 75256 521660 75268
rect 174832 75228 521660 75256
rect 521654 75216 521660 75228
rect 521712 75216 521718 75268
rect 1394 75148 1400 75200
rect 1452 75188 1458 75200
rect 130654 75188 130660 75200
rect 1452 75160 130660 75188
rect 1452 75148 1458 75160
rect 130654 75148 130660 75160
rect 130712 75148 130718 75200
rect 131482 75148 131488 75200
rect 131540 75188 131546 75200
rect 132310 75188 132316 75200
rect 131540 75160 132316 75188
rect 131540 75148 131546 75160
rect 132310 75148 132316 75160
rect 132368 75148 132374 75200
rect 132954 75148 132960 75200
rect 133012 75188 133018 75200
rect 133322 75188 133328 75200
rect 133012 75160 133328 75188
rect 133012 75148 133018 75160
rect 133322 75148 133328 75160
rect 133380 75148 133386 75200
rect 134334 75148 134340 75200
rect 134392 75188 134398 75200
rect 134978 75188 134984 75200
rect 134392 75160 134984 75188
rect 134392 75148 134398 75160
rect 134978 75148 134984 75160
rect 135036 75148 135042 75200
rect 135530 75148 135536 75200
rect 135588 75188 135594 75200
rect 136542 75188 136548 75200
rect 135588 75160 136548 75188
rect 135588 75148 135594 75160
rect 136542 75148 136548 75160
rect 136600 75148 136606 75200
rect 138382 75148 138388 75200
rect 138440 75188 138446 75200
rect 139026 75188 139032 75200
rect 138440 75160 139032 75188
rect 138440 75148 138446 75160
rect 139026 75148 139032 75160
rect 139084 75148 139090 75200
rect 140130 75148 140136 75200
rect 140188 75188 140194 75200
rect 140958 75188 140964 75200
rect 140188 75160 140964 75188
rect 140188 75148 140194 75160
rect 140958 75148 140964 75160
rect 141016 75148 141022 75200
rect 141050 75148 141056 75200
rect 141108 75188 141114 75200
rect 141970 75188 141976 75200
rect 141108 75160 141976 75188
rect 141108 75148 141114 75160
rect 141970 75148 141976 75160
rect 142028 75148 142034 75200
rect 146478 75148 146484 75200
rect 146536 75188 146542 75200
rect 147030 75188 147036 75200
rect 146536 75160 147036 75188
rect 146536 75148 146542 75160
rect 147030 75148 147036 75160
rect 147088 75148 147094 75200
rect 163038 75148 163044 75200
rect 163096 75188 163102 75200
rect 163866 75188 163872 75200
rect 163096 75160 163872 75188
rect 163096 75148 163102 75160
rect 163866 75148 163872 75160
rect 163924 75148 163930 75200
rect 167086 75148 167092 75200
rect 167144 75188 167150 75200
rect 167822 75188 167828 75200
rect 167144 75160 167828 75188
rect 167144 75148 167150 75160
rect 167822 75148 167828 75160
rect 167880 75148 167886 75200
rect 171134 75148 171140 75200
rect 171192 75188 171198 75200
rect 172238 75188 172244 75200
rect 171192 75160 172244 75188
rect 171192 75148 171198 75160
rect 172238 75148 172244 75160
rect 172296 75148 172302 75200
rect 173434 75148 173440 75200
rect 173492 75188 173498 75200
rect 549254 75188 549260 75200
rect 173492 75160 549260 75188
rect 173492 75148 173498 75160
rect 549254 75148 549260 75160
rect 549312 75148 549318 75200
rect 138014 75080 138020 75132
rect 138072 75120 138078 75132
rect 139118 75120 139124 75132
rect 138072 75092 139124 75120
rect 138072 75080 138078 75092
rect 139118 75080 139124 75092
rect 139176 75080 139182 75132
rect 145742 75080 145748 75132
rect 145800 75120 145806 75132
rect 146018 75120 146024 75132
rect 145800 75092 146024 75120
rect 145800 75080 145806 75092
rect 146018 75080 146024 75092
rect 146076 75080 146082 75132
rect 146754 75080 146760 75132
rect 146812 75120 146818 75132
rect 147122 75120 147128 75132
rect 146812 75092 147128 75120
rect 146812 75080 146818 75092
rect 147122 75080 147128 75092
rect 147180 75080 147186 75132
rect 149422 75080 149428 75132
rect 149480 75120 149486 75132
rect 149974 75120 149980 75132
rect 149480 75092 149980 75120
rect 149480 75080 149486 75092
rect 149974 75080 149980 75092
rect 150032 75080 150038 75132
rect 151998 75080 152004 75132
rect 152056 75120 152062 75132
rect 152734 75120 152740 75132
rect 152056 75092 152740 75120
rect 152056 75080 152062 75092
rect 152734 75080 152740 75092
rect 152792 75080 152798 75132
rect 163314 75080 163320 75132
rect 163372 75120 163378 75132
rect 163682 75120 163688 75132
rect 163372 75092 163688 75120
rect 163372 75080 163378 75092
rect 163682 75080 163688 75092
rect 163740 75080 163746 75132
rect 167362 75080 167368 75132
rect 167420 75120 167426 75132
rect 167638 75120 167644 75132
rect 167420 75092 167644 75120
rect 167420 75080 167426 75092
rect 167638 75080 167644 75092
rect 167696 75080 167702 75132
rect 172606 75080 172612 75132
rect 172664 75120 172670 75132
rect 173342 75120 173348 75132
rect 172664 75092 173348 75120
rect 172664 75080 172670 75092
rect 173342 75080 173348 75092
rect 173400 75080 173406 75132
rect 174354 75080 174360 75132
rect 174412 75120 174418 75132
rect 175182 75120 175188 75132
rect 174412 75092 175188 75120
rect 174412 75080 174418 75092
rect 175182 75080 175188 75092
rect 175240 75080 175246 75132
rect 149330 75012 149336 75064
rect 149388 75052 149394 75064
rect 150158 75052 150164 75064
rect 149388 75024 150164 75052
rect 149388 75012 149394 75024
rect 150158 75012 150164 75024
rect 150216 75012 150222 75064
rect 157886 75012 157892 75064
rect 157944 75052 157950 75064
rect 170674 75052 170680 75064
rect 157944 75024 170680 75052
rect 157944 75012 157950 75024
rect 170674 75012 170680 75024
rect 170732 75012 170738 75064
rect 120718 74196 120724 74248
rect 120776 74236 120782 74248
rect 135162 74236 135168 74248
rect 120776 74208 135168 74236
rect 120776 74196 120782 74208
rect 135162 74196 135168 74208
rect 135220 74196 135226 74248
rect 168098 74196 168104 74248
rect 168156 74236 168162 74248
rect 185578 74236 185584 74248
rect 168156 74208 185584 74236
rect 168156 74196 168162 74208
rect 185578 74196 185584 74208
rect 185636 74196 185642 74248
rect 114554 74128 114560 74180
rect 114612 74168 114618 74180
rect 139486 74168 139492 74180
rect 114612 74140 139492 74168
rect 114612 74128 114618 74140
rect 139486 74128 139492 74140
rect 139544 74128 139550 74180
rect 150250 74128 150256 74180
rect 150308 74168 150314 74180
rect 202138 74168 202144 74180
rect 150308 74140 202144 74168
rect 150308 74128 150314 74140
rect 202138 74128 202144 74140
rect 202196 74128 202202 74180
rect 82814 74060 82820 74112
rect 82872 74100 82878 74112
rect 136910 74100 136916 74112
rect 82872 74072 136916 74100
rect 82872 74060 82878 74072
rect 136910 74060 136916 74072
rect 136968 74060 136974 74112
rect 148594 74060 148600 74112
rect 148652 74100 148658 74112
rect 230474 74100 230480 74112
rect 148652 74072 230480 74100
rect 148652 74060 148658 74072
rect 230474 74060 230480 74072
rect 230532 74060 230538 74112
rect 64874 73992 64880 74044
rect 64932 74032 64938 74044
rect 136174 74032 136180 74044
rect 64932 74004 136180 74032
rect 64932 73992 64938 74004
rect 136174 73992 136180 74004
rect 136232 73992 136238 74044
rect 150986 73992 150992 74044
rect 151044 74032 151050 74044
rect 259454 74032 259460 74044
rect 151044 74004 259460 74032
rect 151044 73992 151050 74004
rect 259454 73992 259460 74004
rect 259512 73992 259518 74044
rect 28994 73924 29000 73976
rect 29052 73964 29058 73976
rect 132586 73964 132592 73976
rect 29052 73936 132592 73964
rect 29052 73924 29058 73936
rect 132586 73924 132592 73936
rect 132644 73924 132650 73976
rect 155310 73924 155316 73976
rect 155368 73964 155374 73976
rect 266354 73964 266360 73976
rect 155368 73936 266360 73964
rect 155368 73924 155374 73936
rect 266354 73924 266360 73936
rect 266412 73924 266418 73976
rect 16574 73856 16580 73908
rect 16632 73896 16638 73908
rect 131850 73896 131856 73908
rect 16632 73868 131856 73896
rect 16632 73856 16638 73868
rect 131850 73856 131856 73868
rect 131908 73856 131914 73908
rect 151538 73856 151544 73908
rect 151596 73896 151602 73908
rect 273254 73896 273260 73908
rect 151596 73868 273260 73896
rect 151596 73856 151602 73868
rect 273254 73856 273260 73868
rect 273312 73856 273318 73908
rect 2866 73788 2872 73840
rect 2924 73828 2930 73840
rect 130746 73828 130752 73840
rect 2924 73800 130752 73828
rect 2924 73788 2930 73800
rect 130746 73788 130752 73800
rect 130804 73788 130810 73840
rect 158254 73788 158260 73840
rect 158312 73828 158318 73840
rect 343634 73828 343640 73840
rect 158312 73800 343640 73828
rect 158312 73788 158318 73800
rect 343634 73788 343640 73800
rect 343692 73788 343698 73840
rect 158530 73720 158536 73772
rect 158588 73760 158594 73772
rect 159818 73760 159824 73772
rect 158588 73732 159824 73760
rect 158588 73720 158594 73732
rect 159818 73720 159824 73732
rect 159876 73720 159882 73772
rect 133874 73244 133880 73296
rect 133932 73284 133938 73296
rect 140590 73284 140596 73296
rect 133932 73256 140596 73284
rect 133932 73244 133938 73256
rect 140590 73244 140596 73256
rect 140648 73244 140654 73296
rect 176194 73244 176200 73296
rect 176252 73284 176258 73296
rect 177942 73284 177948 73296
rect 176252 73256 177948 73284
rect 176252 73244 176258 73256
rect 177942 73244 177948 73256
rect 178000 73244 178006 73296
rect 136910 73176 136916 73228
rect 136968 73216 136974 73228
rect 141418 73216 141424 73228
rect 136968 73188 141424 73216
rect 136968 73176 136974 73188
rect 141418 73176 141424 73188
rect 141476 73176 141482 73228
rect 176010 73108 176016 73160
rect 176068 73148 176074 73160
rect 580166 73148 580172 73160
rect 176068 73120 580172 73148
rect 176068 73108 176074 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 175826 73040 175832 73092
rect 175884 73080 175890 73092
rect 176194 73080 176200 73092
rect 175884 73052 176200 73080
rect 175884 73040 175890 73052
rect 176194 73040 176200 73052
rect 176252 73040 176258 73092
rect 175274 72836 175280 72888
rect 175332 72876 175338 72888
rect 176102 72876 176108 72888
rect 175332 72848 176108 72876
rect 175332 72836 175338 72848
rect 176102 72836 176108 72848
rect 176160 72836 176166 72888
rect 153930 72768 153936 72820
rect 153988 72808 153994 72820
rect 293954 72808 293960 72820
rect 153988 72780 293960 72808
rect 153988 72768 153994 72780
rect 293954 72768 293960 72780
rect 294012 72768 294018 72820
rect 154390 72700 154396 72752
rect 154448 72740 154454 72752
rect 300854 72740 300860 72752
rect 154448 72712 300860 72740
rect 154448 72700 154454 72712
rect 300854 72700 300860 72712
rect 300912 72700 300918 72752
rect 155770 72632 155776 72684
rect 155828 72672 155834 72684
rect 316126 72672 316132 72684
rect 155828 72644 316132 72672
rect 155828 72632 155834 72644
rect 316126 72632 316132 72644
rect 316184 72632 316190 72684
rect 107654 72564 107660 72616
rect 107712 72604 107718 72616
rect 138934 72604 138940 72616
rect 107712 72576 138940 72604
rect 107712 72564 107718 72576
rect 138934 72564 138940 72576
rect 138992 72564 138998 72616
rect 155678 72564 155684 72616
rect 155736 72604 155742 72616
rect 322934 72604 322940 72616
rect 155736 72576 322940 72604
rect 155736 72564 155742 72576
rect 322934 72564 322940 72576
rect 322992 72564 322998 72616
rect 57974 72496 57980 72548
rect 58032 72536 58038 72548
rect 135070 72536 135076 72548
rect 58032 72508 135076 72536
rect 58032 72496 58038 72508
rect 135070 72496 135076 72508
rect 135128 72496 135134 72548
rect 165430 72496 165436 72548
rect 165488 72536 165494 72548
rect 347774 72536 347780 72548
rect 165488 72508 347780 72536
rect 165488 72496 165494 72508
rect 347774 72496 347780 72508
rect 347832 72496 347838 72548
rect 14 72428 20 72480
rect 72 72468 78 72480
rect 130286 72468 130292 72480
rect 72 72440 130292 72468
rect 72 72428 78 72440
rect 130286 72428 130292 72440
rect 130344 72428 130350 72480
rect 159818 72428 159824 72480
rect 159876 72468 159882 72480
rect 354674 72468 354680 72480
rect 159876 72440 354680 72468
rect 159876 72428 159882 72440
rect 354674 72428 354680 72440
rect 354732 72428 354738 72480
rect 130378 72156 130384 72208
rect 130436 72196 130442 72208
rect 136266 72196 136272 72208
rect 130436 72168 136272 72196
rect 130436 72156 130442 72168
rect 136266 72156 136272 72168
rect 136324 72156 136330 72208
rect 135622 71748 135628 71800
rect 135680 71788 135686 71800
rect 139394 71788 139400 71800
rect 135680 71760 139400 71788
rect 135680 71748 135686 71760
rect 139394 71748 139400 71760
rect 139452 71748 139458 71800
rect 3418 71680 3424 71732
rect 3476 71720 3482 71732
rect 24210 71720 24216 71732
rect 3476 71692 24216 71720
rect 3476 71680 3482 71692
rect 24210 71680 24216 71692
rect 24268 71680 24274 71732
rect 158622 71136 158628 71188
rect 158680 71176 158686 71188
rect 309134 71176 309140 71188
rect 158680 71148 309140 71176
rect 158680 71136 158686 71148
rect 309134 71136 309140 71148
rect 309192 71136 309198 71188
rect 159634 71068 159640 71120
rect 159692 71108 159698 71120
rect 360194 71108 360200 71120
rect 159692 71080 360200 71108
rect 159692 71068 159698 71080
rect 360194 71068 360200 71080
rect 360252 71068 360258 71120
rect 53834 71000 53840 71052
rect 53892 71040 53898 71052
rect 134886 71040 134892 71052
rect 53892 71012 134892 71040
rect 53892 71000 53898 71012
rect 134886 71000 134892 71012
rect 134944 71000 134950 71052
rect 144362 71000 144368 71052
rect 144420 71040 144426 71052
rect 175274 71040 175280 71052
rect 144420 71012 175280 71040
rect 144420 71000 144426 71012
rect 175274 71000 175280 71012
rect 175332 71000 175338 71052
rect 176470 71000 176476 71052
rect 176528 71040 176534 71052
rect 487154 71040 487160 71052
rect 176528 71012 487160 71040
rect 176528 71000 176534 71012
rect 487154 71000 487160 71012
rect 487212 71000 487218 71052
rect 144178 69912 144184 69964
rect 144236 69952 144242 69964
rect 178034 69952 178040 69964
rect 144236 69924 178040 69952
rect 144236 69912 144242 69924
rect 178034 69912 178040 69924
rect 178092 69912 178098 69964
rect 163774 69844 163780 69896
rect 163832 69884 163838 69896
rect 415394 69884 415400 69896
rect 163832 69856 415400 69884
rect 163832 69844 163838 69856
rect 415394 69844 415400 69856
rect 415452 69844 415458 69896
rect 166350 69776 166356 69828
rect 166408 69816 166414 69828
rect 451274 69816 451280 69828
rect 166408 69788 451280 69816
rect 166408 69776 166414 69788
rect 451274 69776 451280 69788
rect 451332 69776 451338 69828
rect 143074 69708 143080 69760
rect 143132 69748 143138 69760
rect 151078 69748 151084 69760
rect 143132 69720 151084 69748
rect 143132 69708 143138 69720
rect 151078 69708 151084 69720
rect 151136 69708 151142 69760
rect 169018 69708 169024 69760
rect 169076 69748 169082 69760
rect 498194 69748 498200 69760
rect 169076 69720 498200 69748
rect 169076 69708 169082 69720
rect 498194 69708 498200 69720
rect 498252 69708 498258 69760
rect 5534 69640 5540 69692
rect 5592 69680 5598 69692
rect 130010 69680 130016 69692
rect 5592 69652 130016 69680
rect 5592 69640 5598 69652
rect 130010 69640 130016 69652
rect 130068 69640 130074 69692
rect 174722 69640 174728 69692
rect 174780 69680 174786 69692
rect 561674 69680 561680 69692
rect 174780 69652 561680 69680
rect 174780 69640 174786 69652
rect 561674 69640 561680 69652
rect 561732 69640 561738 69692
rect 142798 68960 142804 69012
rect 142856 69000 142862 69012
rect 145558 69000 145564 69012
rect 142856 68972 145564 69000
rect 142856 68960 142862 68972
rect 145558 68960 145564 68972
rect 145616 68960 145622 69012
rect 145834 68484 145840 68536
rect 145892 68524 145898 68536
rect 195974 68524 195980 68536
rect 145892 68496 195980 68524
rect 145892 68484 145898 68496
rect 195974 68484 195980 68496
rect 196032 68484 196038 68536
rect 164878 68416 164884 68468
rect 164936 68456 164942 68468
rect 433334 68456 433340 68468
rect 164936 68428 433340 68456
rect 164936 68416 164942 68428
rect 433334 68416 433340 68428
rect 433392 68416 433398 68468
rect 166258 68348 166264 68400
rect 166316 68388 166322 68400
rect 456794 68388 456800 68400
rect 166316 68360 456800 68388
rect 166316 68348 166322 68360
rect 456794 68348 456800 68360
rect 456852 68348 456858 68400
rect 170582 68280 170588 68332
rect 170640 68320 170646 68332
rect 514846 68320 514852 68332
rect 170640 68292 514852 68320
rect 170640 68280 170646 68292
rect 514846 68280 514852 68292
rect 514904 68280 514910 68332
rect 145374 67124 145380 67176
rect 145432 67164 145438 67176
rect 193214 67164 193220 67176
rect 145432 67136 193220 67164
rect 145432 67124 145438 67136
rect 193214 67124 193220 67136
rect 193272 67124 193278 67176
rect 159266 67056 159272 67108
rect 159324 67096 159330 67108
rect 365714 67096 365720 67108
rect 159324 67068 365720 67096
rect 159324 67056 159330 67068
rect 365714 67056 365720 67068
rect 365772 67056 365778 67108
rect 167546 66988 167552 67040
rect 167604 67028 167610 67040
rect 473354 67028 473360 67040
rect 167604 67000 473360 67028
rect 167604 66988 167610 67000
rect 473354 66988 473360 67000
rect 473412 66988 473418 67040
rect 170306 66920 170312 66972
rect 170364 66960 170370 66972
rect 511994 66960 512000 66972
rect 170364 66932 512000 66960
rect 170364 66920 170370 66932
rect 511994 66920 512000 66932
rect 512052 66920 512058 66972
rect 171778 66852 171784 66904
rect 171836 66892 171842 66904
rect 529934 66892 529940 66904
rect 171836 66864 529940 66892
rect 171836 66852 171842 66864
rect 529934 66852 529940 66864
rect 529992 66852 529998 66904
rect 153838 65900 153844 65952
rect 153896 65940 153902 65952
rect 295334 65940 295340 65952
rect 153896 65912 295340 65940
rect 153896 65900 153902 65912
rect 295334 65900 295340 65912
rect 295392 65900 295398 65952
rect 155218 65832 155224 65884
rect 155276 65872 155282 65884
rect 307754 65872 307760 65884
rect 155276 65844 307760 65872
rect 155276 65832 155282 65844
rect 307754 65832 307760 65844
rect 307812 65832 307818 65884
rect 3510 65764 3516 65816
rect 3568 65804 3574 65816
rect 190638 65804 190644 65816
rect 3568 65776 190644 65804
rect 3568 65764 3574 65776
rect 190638 65764 190644 65776
rect 190696 65764 190702 65816
rect 164786 65696 164792 65748
rect 164844 65736 164850 65748
rect 437474 65736 437480 65748
rect 164844 65708 437480 65736
rect 164844 65696 164850 65708
rect 437474 65696 437480 65708
rect 437532 65696 437538 65748
rect 170214 65628 170220 65680
rect 170272 65668 170278 65680
rect 510614 65668 510620 65680
rect 170272 65640 510620 65668
rect 170272 65628 170278 65640
rect 510614 65628 510620 65640
rect 510672 65628 510678 65680
rect 174538 65560 174544 65612
rect 174596 65600 174602 65612
rect 564434 65600 564440 65612
rect 174596 65572 564440 65600
rect 174596 65560 174602 65572
rect 564434 65560 564440 65572
rect 564492 65560 564498 65612
rect 174630 65492 174636 65544
rect 174688 65532 174694 65544
rect 568574 65532 568580 65544
rect 174688 65504 568580 65532
rect 174688 65492 174694 65504
rect 568574 65492 568580 65504
rect 568632 65492 568638 65544
rect 165246 64336 165252 64388
rect 165304 64376 165310 64388
rect 382274 64376 382280 64388
rect 165304 64348 382280 64376
rect 165304 64336 165310 64348
rect 382274 64336 382280 64348
rect 382332 64336 382338 64388
rect 163498 64268 163504 64320
rect 163556 64308 163562 64320
rect 419534 64308 419540 64320
rect 163556 64280 419540 64308
rect 163556 64268 163562 64280
rect 419534 64268 419540 64280
rect 419592 64268 419598 64320
rect 163590 64200 163596 64252
rect 163648 64240 163654 64252
rect 423674 64240 423680 64252
rect 163648 64212 423680 64240
rect 163648 64200 163654 64212
rect 423674 64200 423680 64212
rect 423732 64200 423738 64252
rect 173802 64132 173808 64184
rect 173860 64172 173866 64184
rect 552014 64172 552020 64184
rect 173860 64144 552020 64172
rect 173860 64132 173866 64144
rect 552014 64132 552020 64144
rect 552072 64132 552078 64184
rect 144086 63248 144092 63300
rect 144144 63288 144150 63300
rect 145650 63288 145656 63300
rect 144144 63260 145656 63288
rect 144144 63248 144150 63260
rect 145650 63248 145656 63260
rect 145708 63248 145714 63300
rect 166626 62840 166632 62892
rect 166684 62880 166690 62892
rect 361574 62880 361580 62892
rect 166684 62852 361580 62880
rect 166684 62840 166690 62852
rect 361574 62840 361580 62852
rect 361632 62840 361638 62892
rect 168926 62772 168932 62824
rect 168984 62812 168990 62824
rect 488534 62812 488540 62824
rect 168984 62784 488540 62812
rect 168984 62772 168990 62784
rect 488534 62772 488540 62784
rect 488592 62772 488598 62824
rect 148410 61548 148416 61600
rect 148468 61588 148474 61600
rect 223574 61588 223580 61600
rect 148468 61560 223580 61588
rect 148468 61548 148474 61560
rect 223574 61548 223580 61560
rect 223632 61548 223638 61600
rect 152550 61480 152556 61532
rect 152608 61520 152614 61532
rect 277394 61520 277400 61532
rect 152608 61492 277400 61520
rect 152608 61480 152614 61492
rect 277394 61480 277400 61492
rect 277452 61480 277458 61532
rect 160830 61412 160836 61464
rect 160888 61452 160894 61464
rect 380894 61452 380900 61464
rect 160888 61424 380900 61452
rect 160888 61412 160894 61424
rect 380894 61412 380900 61424
rect 380952 61412 380958 61464
rect 171686 61344 171692 61396
rect 171744 61384 171750 61396
rect 525794 61384 525800 61396
rect 171744 61356 525800 61384
rect 171744 61344 171750 61356
rect 525794 61344 525800 61356
rect 525852 61344 525858 61396
rect 192662 60664 192668 60716
rect 192720 60704 192726 60716
rect 580166 60704 580172 60716
rect 192720 60676 580172 60704
rect 192720 60664 192726 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 170122 60052 170128 60104
rect 170180 60092 170186 60104
rect 506566 60092 506572 60104
rect 170180 60064 506572 60092
rect 170180 60052 170186 60064
rect 506566 60052 506572 60064
rect 506624 60052 506630 60104
rect 176378 59984 176384 60036
rect 176436 60024 176442 60036
rect 539594 60024 539600 60036
rect 176436 59996 539600 60024
rect 176436 59984 176442 59996
rect 539594 59984 539600 59996
rect 539652 59984 539658 60036
rect 156598 58624 156604 58676
rect 156656 58664 156662 58676
rect 333974 58664 333980 58676
rect 156656 58636 333980 58664
rect 156656 58624 156662 58636
rect 333974 58624 333980 58636
rect 334032 58624 334038 58676
rect 42794 57196 42800 57248
rect 42852 57236 42858 57248
rect 129366 57236 129372 57248
rect 42852 57208 129372 57236
rect 42852 57196 42858 57208
rect 129366 57196 129372 57208
rect 129424 57196 129430 57248
rect 157794 55836 157800 55888
rect 157852 55876 157858 55888
rect 346394 55876 346400 55888
rect 157852 55848 346400 55876
rect 157852 55836 157858 55848
rect 346394 55836 346400 55848
rect 346452 55836 346458 55888
rect 142706 51688 142712 51740
rect 142764 51728 142770 51740
rect 153838 51728 153844 51740
rect 142764 51700 153844 51728
rect 142764 51688 142770 51700
rect 153838 51688 153844 51700
rect 153896 51688 153902 51740
rect 160738 51688 160744 51740
rect 160796 51728 160802 51740
rect 390554 51728 390560 51740
rect 160796 51700 390560 51728
rect 160796 51688 160802 51700
rect 390554 51688 390560 51700
rect 390612 51688 390618 51740
rect 124214 51076 124220 51128
rect 124272 51116 124278 51128
rect 127618 51116 127624 51128
rect 124272 51088 127624 51116
rect 124272 51076 124278 51088
rect 127618 51076 127624 51088
rect 127676 51076 127682 51128
rect 148318 48968 148324 49020
rect 148376 49008 148382 49020
rect 226334 49008 226340 49020
rect 148376 48980 226340 49008
rect 148376 48968 148382 48980
rect 226334 48968 226340 48980
rect 226392 48968 226398 49020
rect 118510 46860 118516 46912
rect 118568 46900 118574 46912
rect 580166 46900 580172 46912
rect 118568 46872 580172 46900
rect 118568 46860 118574 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 3418 45500 3424 45552
rect 3476 45540 3482 45552
rect 178218 45540 178224 45552
rect 3476 45512 178224 45540
rect 3476 45500 3482 45512
rect 178218 45500 178224 45512
rect 178276 45500 178282 45552
rect 141326 44888 141332 44940
rect 141384 44928 141390 44940
rect 142890 44928 142896 44940
rect 141384 44900 142896 44928
rect 141384 44888 141390 44900
rect 142890 44888 142896 44900
rect 142948 44888 142954 44940
rect 38654 44820 38660 44872
rect 38712 44860 38718 44872
rect 133046 44860 133052 44872
rect 38712 44832 133052 44860
rect 38712 44820 38718 44832
rect 133046 44820 133052 44832
rect 133104 44820 133110 44872
rect 177206 44820 177212 44872
rect 177264 44860 177270 44872
rect 432046 44860 432052 44872
rect 177264 44832 432052 44860
rect 177264 44820 177270 44832
rect 432046 44820 432052 44832
rect 432104 44820 432110 44872
rect 142614 44140 142620 44192
rect 142672 44180 142678 44192
rect 144270 44180 144276 44192
rect 142672 44152 144276 44180
rect 142672 44140 142678 44152
rect 144270 44140 144276 44152
rect 144328 44140 144334 44192
rect 19334 39312 19340 39364
rect 19392 39352 19398 39364
rect 129274 39352 129280 39364
rect 19392 39324 129280 39352
rect 19392 39312 19398 39324
rect 129274 39312 129280 39324
rect 129332 39312 129338 39364
rect 146938 35640 146944 35692
rect 146996 35680 147002 35692
rect 205634 35680 205640 35692
rect 146996 35652 205640 35680
rect 146996 35640 147002 35652
rect 205634 35640 205640 35652
rect 205692 35640 205698 35692
rect 146846 35572 146852 35624
rect 146904 35612 146910 35624
rect 209866 35612 209872 35624
rect 146904 35584 209872 35612
rect 146904 35572 146910 35584
rect 209866 35572 209872 35584
rect 209924 35572 209930 35624
rect 150894 35504 150900 35556
rect 150952 35544 150958 35556
rect 255314 35544 255320 35556
rect 150952 35516 255320 35544
rect 150952 35504 150958 35516
rect 255314 35504 255320 35516
rect 255372 35504 255378 35556
rect 155126 35436 155132 35488
rect 155184 35476 155190 35488
rect 311894 35476 311900 35488
rect 155184 35448 311900 35476
rect 155184 35436 155190 35448
rect 311894 35436 311900 35448
rect 311952 35436 311958 35488
rect 167914 35368 167920 35420
rect 167972 35408 167978 35420
rect 375374 35408 375380 35420
rect 167972 35380 375380 35408
rect 167972 35368 167978 35380
rect 375374 35368 375380 35380
rect 375432 35368 375438 35420
rect 176194 35300 176200 35352
rect 176252 35340 176258 35352
rect 397454 35340 397460 35352
rect 176252 35312 397460 35340
rect 176252 35300 176258 35312
rect 397454 35300 397460 35312
rect 397512 35300 397518 35352
rect 176286 35232 176292 35284
rect 176344 35272 176350 35284
rect 404354 35272 404360 35284
rect 176344 35244 404360 35272
rect 176344 35232 176350 35244
rect 404354 35232 404360 35244
rect 404412 35232 404418 35284
rect 163406 35164 163412 35216
rect 163464 35204 163470 35216
rect 422294 35204 422300 35216
rect 163464 35176 422300 35204
rect 163464 35164 163470 35176
rect 422294 35164 422300 35176
rect 422352 35164 422358 35216
rect 145190 34280 145196 34332
rect 145248 34320 145254 34332
rect 187694 34320 187700 34332
rect 145248 34292 187700 34320
rect 145248 34280 145254 34292
rect 187694 34280 187700 34292
rect 187752 34280 187758 34332
rect 145098 34212 145104 34264
rect 145156 34252 145162 34264
rect 194594 34252 194600 34264
rect 145156 34224 194600 34252
rect 145156 34212 145162 34224
rect 194594 34212 194600 34224
rect 194652 34212 194658 34264
rect 145282 34144 145288 34196
rect 145340 34184 145346 34196
rect 198734 34184 198740 34196
rect 145340 34156 198740 34184
rect 145340 34144 145346 34156
rect 198734 34144 198740 34156
rect 198792 34144 198798 34196
rect 148226 34076 148232 34128
rect 148284 34116 148290 34128
rect 226426 34116 226432 34128
rect 148284 34088 226432 34116
rect 148284 34076 148290 34088
rect 226426 34076 226432 34088
rect 226484 34076 226490 34128
rect 149790 34008 149796 34060
rect 149848 34048 149854 34060
rect 241514 34048 241520 34060
rect 149848 34020 241520 34048
rect 149848 34008 149854 34020
rect 241514 34008 241520 34020
rect 241572 34008 241578 34060
rect 152458 33940 152464 33992
rect 152516 33980 152522 33992
rect 280154 33980 280160 33992
rect 152516 33952 280160 33980
rect 152516 33940 152522 33952
rect 280154 33940 280160 33952
rect 280212 33940 280218 33992
rect 153746 33872 153752 33924
rect 153804 33912 153810 33924
rect 291194 33912 291200 33924
rect 153804 33884 291200 33912
rect 153804 33872 153810 33884
rect 291194 33872 291200 33884
rect 291252 33872 291258 33924
rect 157702 33804 157708 33856
rect 157760 33844 157766 33856
rect 350534 33844 350540 33856
rect 157760 33816 350540 33844
rect 157760 33804 157766 33816
rect 350534 33804 350540 33816
rect 350592 33804 350598 33856
rect 164694 33736 164700 33788
rect 164752 33776 164758 33788
rect 441614 33776 441620 33788
rect 164752 33748 441620 33776
rect 164752 33736 164758 33748
rect 441614 33736 441620 33748
rect 441672 33736 441678 33788
rect 3510 33056 3516 33108
rect 3568 33096 3574 33108
rect 23014 33096 23020 33108
rect 3568 33068 23020 33096
rect 3568 33056 3574 33068
rect 23014 33056 23020 33068
rect 23072 33056 23078 33108
rect 177942 33056 177948 33108
rect 178000 33096 178006 33108
rect 580166 33096 580172 33108
rect 178000 33068 580172 33096
rect 178000 33056 178006 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 146754 32852 146760 32904
rect 146812 32892 146818 32904
rect 212534 32892 212540 32904
rect 146812 32864 212540 32892
rect 146812 32852 146818 32864
rect 212534 32852 212540 32864
rect 212592 32852 212598 32904
rect 148134 32784 148140 32836
rect 148192 32824 148198 32836
rect 219434 32824 219440 32836
rect 148192 32796 219440 32824
rect 148192 32784 148198 32796
rect 219434 32784 219440 32796
rect 219492 32784 219498 32836
rect 149698 32716 149704 32768
rect 149756 32756 149762 32768
rect 237374 32756 237380 32768
rect 149756 32728 237380 32756
rect 149756 32716 149762 32728
rect 237374 32716 237380 32728
rect 237432 32716 237438 32768
rect 3418 32648 3424 32700
rect 3476 32688 3482 32700
rect 178126 32688 178132 32700
rect 3476 32660 178132 32688
rect 3476 32648 3482 32660
rect 178126 32648 178132 32660
rect 178184 32648 178190 32700
rect 162026 32580 162032 32632
rect 162084 32620 162090 32632
rect 400214 32620 400220 32632
rect 162084 32592 400220 32620
rect 162084 32580 162090 32592
rect 400214 32580 400220 32592
rect 400272 32580 400278 32632
rect 163314 32512 163320 32564
rect 163372 32552 163378 32564
rect 423766 32552 423772 32564
rect 163372 32524 423772 32552
rect 163372 32512 163378 32524
rect 423766 32512 423772 32524
rect 423824 32512 423830 32564
rect 164510 32444 164516 32496
rect 164568 32484 164574 32496
rect 434714 32484 434720 32496
rect 164568 32456 434720 32484
rect 164568 32444 164574 32456
rect 434714 32444 434720 32456
rect 434772 32444 434778 32496
rect 164602 32376 164608 32428
rect 164660 32416 164666 32428
rect 438854 32416 438860 32428
rect 164660 32388 438860 32416
rect 164660 32376 164666 32388
rect 438854 32376 438860 32388
rect 438912 32376 438918 32428
rect 145006 31356 145012 31408
rect 145064 31396 145070 31408
rect 185026 31396 185032 31408
rect 145064 31368 185032 31396
rect 145064 31356 145070 31368
rect 185026 31356 185032 31368
rect 185084 31356 185090 31408
rect 153654 31288 153660 31340
rect 153712 31328 153718 31340
rect 292666 31328 292672 31340
rect 153712 31300 292672 31328
rect 153712 31288 153718 31300
rect 292666 31288 292672 31300
rect 292724 31288 292730 31340
rect 153562 31220 153568 31272
rect 153620 31260 153626 31272
rect 299474 31260 299480 31272
rect 153620 31232 299480 31260
rect 153620 31220 153626 31232
rect 299474 31220 299480 31232
rect 299532 31220 299538 31272
rect 158346 31152 158352 31204
rect 158404 31192 158410 31204
rect 339494 31192 339500 31204
rect 158404 31164 339500 31192
rect 158404 31152 158410 31164
rect 339494 31152 339500 31164
rect 339552 31152 339558 31204
rect 159174 31084 159180 31136
rect 159232 31124 159238 31136
rect 374086 31124 374092 31136
rect 159232 31096 374092 31124
rect 159232 31084 159238 31096
rect 374086 31084 374092 31096
rect 374144 31084 374150 31136
rect 168834 31016 168840 31068
rect 168892 31056 168898 31068
rect 496814 31056 496820 31068
rect 168892 31028 496820 31056
rect 168892 31016 168898 31028
rect 496814 31016 496820 31028
rect 496872 31016 496878 31068
rect 149514 29928 149520 29980
rect 149572 29968 149578 29980
rect 242894 29968 242900 29980
rect 149572 29940 242900 29968
rect 149572 29928 149578 29940
rect 242894 29928 242900 29940
rect 242952 29928 242958 29980
rect 149606 29860 149612 29912
rect 149664 29900 149670 29912
rect 247034 29900 247040 29912
rect 149664 29872 247040 29900
rect 149664 29860 149670 29872
rect 247034 29860 247040 29872
rect 247092 29860 247098 29912
rect 150802 29792 150808 29844
rect 150860 29832 150866 29844
rect 264974 29832 264980 29844
rect 150860 29804 264980 29832
rect 150860 29792 150866 29804
rect 264974 29792 264980 29804
rect 265032 29792 265038 29844
rect 155034 29724 155040 29776
rect 155092 29764 155098 29776
rect 317414 29764 317420 29776
rect 155092 29736 317420 29764
rect 155092 29724 155098 29736
rect 317414 29724 317420 29736
rect 317472 29724 317478 29776
rect 163222 29656 163228 29708
rect 163280 29696 163286 29708
rect 416774 29696 416780 29708
rect 163280 29668 416780 29696
rect 163280 29656 163286 29668
rect 416774 29656 416780 29668
rect 416832 29656 416838 29708
rect 174446 29588 174452 29640
rect 174504 29628 174510 29640
rect 564526 29628 564532 29640
rect 174504 29600 564532 29628
rect 174504 29588 174510 29600
rect 564526 29588 564532 29600
rect 564584 29588 564590 29640
rect 146662 28704 146668 28756
rect 146720 28744 146726 28756
rect 208394 28744 208400 28756
rect 146720 28716 208400 28744
rect 146720 28704 146726 28716
rect 208394 28704 208400 28716
rect 208452 28704 208458 28756
rect 148042 28636 148048 28688
rect 148100 28676 148106 28688
rect 222194 28676 222200 28688
rect 148100 28648 222200 28676
rect 148100 28636 148106 28648
rect 222194 28636 222200 28648
rect 222252 28636 222258 28688
rect 147950 28568 147956 28620
rect 148008 28608 148014 28620
rect 229094 28608 229100 28620
rect 148008 28580 229100 28608
rect 148008 28568 148014 28580
rect 229094 28568 229100 28580
rect 229152 28568 229158 28620
rect 152366 28500 152372 28552
rect 152424 28540 152430 28552
rect 278774 28540 278780 28552
rect 152424 28512 278780 28540
rect 152424 28500 152430 28512
rect 278774 28500 278780 28512
rect 278832 28500 278838 28552
rect 154942 28432 154948 28484
rect 155000 28472 155006 28484
rect 310514 28472 310520 28484
rect 155000 28444 310520 28472
rect 155000 28432 155006 28444
rect 310514 28432 310520 28444
rect 310572 28432 310578 28484
rect 159082 28364 159088 28416
rect 159140 28404 159146 28416
rect 364334 28404 364340 28416
rect 159140 28376 364340 28404
rect 159140 28364 159146 28376
rect 364334 28364 364340 28376
rect 364392 28364 364398 28416
rect 158990 28296 158996 28348
rect 159048 28336 159054 28348
rect 372614 28336 372620 28348
rect 159048 28308 372620 28336
rect 159048 28296 159054 28308
rect 372614 28296 372620 28308
rect 372672 28296 372678 28348
rect 173066 28228 173072 28280
rect 173124 28268 173130 28280
rect 539686 28268 539692 28280
rect 173124 28240 539692 28268
rect 173124 28228 173130 28240
rect 539686 28228 539692 28240
rect 539744 28228 539750 28280
rect 147214 27276 147220 27328
rect 147272 27316 147278 27328
rect 190454 27316 190460 27328
rect 147272 27288 190460 27316
rect 147272 27276 147278 27288
rect 190454 27276 190460 27288
rect 190512 27276 190518 27328
rect 146110 27208 146116 27260
rect 146168 27248 146174 27260
rect 193306 27248 193312 27260
rect 146168 27220 193312 27248
rect 146168 27208 146174 27220
rect 193306 27208 193312 27220
rect 193364 27208 193370 27260
rect 146570 27140 146576 27192
rect 146628 27180 146634 27192
rect 204254 27180 204260 27192
rect 146628 27152 204260 27180
rect 146628 27140 146634 27152
rect 204254 27140 204260 27152
rect 204312 27140 204318 27192
rect 152274 27072 152280 27124
rect 152332 27112 152338 27124
rect 276014 27112 276020 27124
rect 152332 27084 276020 27112
rect 152332 27072 152338 27084
rect 276014 27072 276020 27084
rect 276072 27072 276078 27124
rect 168006 27004 168012 27056
rect 168064 27044 168070 27056
rect 379514 27044 379520 27056
rect 168064 27016 379520 27044
rect 168064 27004 168070 27016
rect 379514 27004 379520 27016
rect 379572 27004 379578 27056
rect 158898 26936 158904 26988
rect 158956 26976 158962 26988
rect 371234 26976 371240 26988
rect 158956 26948 371240 26976
rect 158956 26936 158962 26948
rect 371234 26936 371240 26948
rect 371292 26936 371298 26988
rect 175366 26868 175372 26920
rect 175424 26908 175430 26920
rect 574094 26908 574100 26920
rect 175424 26880 574100 26908
rect 175424 26868 175430 26880
rect 574094 26868 574100 26880
rect 574152 26868 574158 26920
rect 146478 25916 146484 25968
rect 146536 25956 146542 25968
rect 211154 25956 211160 25968
rect 146536 25928 211160 25956
rect 146536 25916 146542 25928
rect 211154 25916 211160 25928
rect 211212 25916 211218 25968
rect 152182 25848 152188 25900
rect 152240 25888 152246 25900
rect 282914 25888 282920 25900
rect 152240 25860 282920 25888
rect 152240 25848 152246 25860
rect 282914 25848 282920 25860
rect 282972 25848 282978 25900
rect 154850 25780 154856 25832
rect 154908 25820 154914 25832
rect 314654 25820 314660 25832
rect 154908 25792 314660 25820
rect 154908 25780 154914 25792
rect 314654 25780 314660 25792
rect 314712 25780 314718 25832
rect 172882 25712 172888 25764
rect 172940 25752 172946 25764
rect 349890 25752 349896 25764
rect 172940 25724 349896 25752
rect 172940 25712 172946 25724
rect 349890 25712 349896 25724
rect 349948 25712 349954 25764
rect 177758 25644 177764 25696
rect 177816 25684 177822 25696
rect 411254 25684 411260 25696
rect 177816 25656 411260 25684
rect 177816 25644 177822 25656
rect 411254 25644 411260 25656
rect 411312 25644 411318 25696
rect 167454 25576 167460 25628
rect 167512 25616 167518 25628
rect 473446 25616 473452 25628
rect 167512 25588 473452 25616
rect 167512 25576 167518 25588
rect 473446 25576 473452 25588
rect 473504 25576 473510 25628
rect 172974 25508 172980 25560
rect 173032 25548 173038 25560
rect 546494 25548 546500 25560
rect 173032 25520 546500 25548
rect 173032 25508 173038 25520
rect 546494 25508 546500 25520
rect 546552 25508 546558 25560
rect 153470 24352 153476 24404
rect 153528 24392 153534 24404
rect 296714 24392 296720 24404
rect 153528 24364 296720 24392
rect 153528 24352 153534 24364
rect 296714 24352 296720 24364
rect 296772 24352 296778 24404
rect 154758 24284 154764 24336
rect 154816 24324 154822 24336
rect 321554 24324 321560 24336
rect 154816 24296 321560 24324
rect 154816 24284 154822 24296
rect 321554 24284 321560 24296
rect 321612 24284 321618 24336
rect 177574 24216 177580 24268
rect 177632 24256 177638 24268
rect 418154 24256 418160 24268
rect 177632 24228 418160 24256
rect 177632 24216 177638 24228
rect 418154 24216 418160 24228
rect 418212 24216 418218 24268
rect 172790 24148 172796 24200
rect 172848 24188 172854 24200
rect 540974 24188 540980 24200
rect 172848 24160 540980 24188
rect 172848 24148 172854 24160
rect 540974 24148 540980 24160
rect 541032 24148 541038 24200
rect 174354 24080 174360 24132
rect 174412 24120 174418 24132
rect 567194 24120 567200 24132
rect 174412 24092 567200 24120
rect 174412 24080 174418 24092
rect 567194 24080 567200 24092
rect 567252 24080 567258 24132
rect 3234 22992 3240 23044
rect 3292 23032 3298 23044
rect 189534 23032 189540 23044
rect 3292 23004 189540 23032
rect 3292 22992 3298 23004
rect 189534 22992 189540 23004
rect 189592 22992 189598 23044
rect 170030 22924 170036 22976
rect 170088 22964 170094 22976
rect 513374 22964 513380 22976
rect 170088 22936 513380 22964
rect 170088 22924 170094 22936
rect 513374 22924 513380 22936
rect 513432 22924 513438 22976
rect 171594 22856 171600 22908
rect 171652 22896 171658 22908
rect 528554 22896 528560 22908
rect 171652 22868 528560 22896
rect 171652 22856 171658 22868
rect 528554 22856 528560 22868
rect 528612 22856 528618 22908
rect 88334 22788 88340 22840
rect 88392 22828 88398 22840
rect 137186 22828 137192 22840
rect 88392 22800 137192 22828
rect 88392 22788 88398 22800
rect 137186 22788 137192 22800
rect 137244 22788 137250 22840
rect 171502 22788 171508 22840
rect 171560 22828 171566 22840
rect 531314 22828 531320 22840
rect 171560 22800 531320 22828
rect 171560 22788 171566 22800
rect 531314 22788 531320 22800
rect 531372 22788 531378 22840
rect 118326 22720 118332 22772
rect 118384 22760 118390 22772
rect 580258 22760 580264 22772
rect 118384 22732 580264 22760
rect 118384 22720 118390 22732
rect 580258 22720 580264 22732
rect 580316 22720 580322 22772
rect 163130 21632 163136 21684
rect 163188 21672 163194 21684
rect 415486 21672 415492 21684
rect 163188 21644 415492 21672
rect 163188 21632 163194 21644
rect 415486 21632 415492 21644
rect 415544 21632 415550 21684
rect 167362 21564 167368 21616
rect 167420 21604 167426 21616
rect 476114 21604 476120 21616
rect 167420 21576 476120 21604
rect 167420 21564 167426 21576
rect 476114 21564 476120 21576
rect 476172 21564 476178 21616
rect 168650 21496 168656 21548
rect 168708 21536 168714 21548
rect 495434 21536 495440 21548
rect 168708 21508 495440 21536
rect 168708 21496 168714 21508
rect 495434 21496 495440 21508
rect 495492 21496 495498 21548
rect 168742 21428 168748 21480
rect 168800 21468 168806 21480
rect 498286 21468 498292 21480
rect 168800 21440 498292 21468
rect 168800 21428 168806 21440
rect 498286 21428 498292 21440
rect 498344 21428 498350 21480
rect 174262 21360 174268 21412
rect 174320 21400 174326 21412
rect 563054 21400 563060 21412
rect 174320 21372 563060 21400
rect 174320 21360 174326 21372
rect 563054 21360 563060 21372
rect 563112 21360 563118 21412
rect 347038 20612 347044 20664
rect 347096 20652 347102 20664
rect 579982 20652 579988 20664
rect 347096 20624 579988 20652
rect 347096 20612 347102 20624
rect 579982 20612 579988 20624
rect 580040 20612 580046 20664
rect 152090 20272 152096 20324
rect 152148 20312 152154 20324
rect 276106 20312 276112 20324
rect 152148 20284 276112 20312
rect 152148 20272 152154 20284
rect 276106 20272 276112 20284
rect 276164 20272 276170 20324
rect 151998 20204 152004 20256
rect 152056 20244 152062 20256
rect 284294 20244 284300 20256
rect 152056 20216 284300 20244
rect 152056 20204 152062 20216
rect 284294 20204 284300 20216
rect 284352 20204 284358 20256
rect 268378 20136 268384 20188
rect 268436 20176 268442 20188
rect 467834 20176 467840 20188
rect 268436 20148 467840 20176
rect 268436 20136 268442 20148
rect 467834 20136 467840 20148
rect 467892 20136 467898 20188
rect 167270 20068 167276 20120
rect 167328 20108 167334 20120
rect 228358 20108 228364 20120
rect 167328 20080 228364 20108
rect 167328 20068 167334 20080
rect 228358 20068 228364 20080
rect 228416 20068 228422 20120
rect 260098 20068 260104 20120
rect 260156 20108 260162 20120
rect 460934 20108 460940 20120
rect 260156 20080 460940 20108
rect 260156 20068 260162 20080
rect 460934 20068 460940 20080
rect 460992 20068 460998 20120
rect 166166 20000 166172 20052
rect 166224 20040 166230 20052
rect 462314 20040 462320 20052
rect 166224 20012 462320 20040
rect 166224 20000 166230 20012
rect 462314 20000 462320 20012
rect 462372 20000 462378 20052
rect 169938 19932 169944 19984
rect 169996 19972 170002 19984
rect 509234 19972 509240 19984
rect 169996 19944 509240 19972
rect 169996 19932 170002 19944
rect 509234 19932 509240 19944
rect 509292 19932 509298 19984
rect 161934 18980 161940 19032
rect 161992 19020 161998 19032
rect 407114 19020 407120 19032
rect 161992 18992 407120 19020
rect 161992 18980 161998 18992
rect 407114 18980 407120 18992
rect 407172 18980 407178 19032
rect 163038 18912 163044 18964
rect 163096 18952 163102 18964
rect 426434 18952 426440 18964
rect 163096 18924 426440 18952
rect 163096 18912 163102 18924
rect 426434 18912 426440 18924
rect 426492 18912 426498 18964
rect 117314 18844 117320 18896
rect 117372 18884 117378 18896
rect 129182 18884 129188 18896
rect 117372 18856 129188 18884
rect 117372 18844 117378 18856
rect 129182 18844 129188 18856
rect 129240 18844 129246 18896
rect 164418 18844 164424 18896
rect 164476 18884 164482 18896
rect 440234 18884 440240 18896
rect 164476 18856 440240 18884
rect 164476 18844 164482 18856
rect 440234 18844 440240 18856
rect 440292 18844 440298 18896
rect 120074 18776 120080 18828
rect 120132 18816 120138 18828
rect 139670 18816 139676 18828
rect 120132 18788 139676 18816
rect 120132 18776 120138 18788
rect 139670 18776 139676 18788
rect 139728 18776 139734 18828
rect 172698 18776 172704 18828
rect 172756 18816 172762 18828
rect 553394 18816 553400 18828
rect 172756 18788 553400 18816
rect 172756 18776 172762 18788
rect 553394 18776 553400 18788
rect 553452 18776 553458 18828
rect 111794 18708 111800 18760
rect 111852 18748 111858 18760
rect 138566 18748 138572 18760
rect 111852 18720 138572 18748
rect 111852 18708 111858 18720
rect 138566 18708 138572 18720
rect 138624 18708 138630 18760
rect 173986 18708 173992 18760
rect 174044 18748 174050 18760
rect 556246 18748 556252 18760
rect 174044 18720 556252 18748
rect 174044 18708 174050 18720
rect 556246 18708 556252 18720
rect 556304 18708 556310 18760
rect 35894 18640 35900 18692
rect 35952 18680 35958 18692
rect 126330 18680 126336 18692
rect 35952 18652 126336 18680
rect 35952 18640 35958 18652
rect 126330 18640 126336 18652
rect 126388 18640 126394 18692
rect 174078 18640 174084 18692
rect 174136 18680 174142 18692
rect 558914 18680 558920 18692
rect 174136 18652 558920 18680
rect 174136 18640 174142 18652
rect 558914 18640 558920 18652
rect 558972 18640 558978 18692
rect 15194 18572 15200 18624
rect 15252 18612 15258 18624
rect 131666 18612 131672 18624
rect 15252 18584 131672 18612
rect 15252 18572 15258 18584
rect 131666 18572 131672 18584
rect 131724 18572 131730 18624
rect 174170 18572 174176 18624
rect 174228 18612 174234 18624
rect 560294 18612 560300 18624
rect 174228 18584 560300 18612
rect 174228 18572 174234 18584
rect 560294 18572 560300 18584
rect 560352 18572 560358 18624
rect 154666 17416 154672 17468
rect 154724 17456 154730 17468
rect 318794 17456 318800 17468
rect 154724 17428 318800 17456
rect 154724 17416 154730 17428
rect 318794 17416 318800 17428
rect 318852 17416 318858 17468
rect 161842 17348 161848 17400
rect 161900 17388 161906 17400
rect 405734 17388 405740 17400
rect 161900 17360 405740 17388
rect 161900 17348 161906 17360
rect 405734 17348 405740 17360
rect 405792 17348 405798 17400
rect 168558 17280 168564 17332
rect 168616 17320 168622 17332
rect 492674 17320 492680 17332
rect 168616 17292 492680 17320
rect 168616 17280 168622 17292
rect 492674 17280 492680 17292
rect 492732 17280 492738 17332
rect 171410 17212 171416 17264
rect 171468 17252 171474 17264
rect 531406 17252 531412 17264
rect 171468 17224 531412 17252
rect 171468 17212 171474 17224
rect 531406 17212 531412 17224
rect 531464 17212 531470 17264
rect 160554 16124 160560 16176
rect 160612 16164 160618 16176
rect 384298 16164 384304 16176
rect 160612 16136 384304 16164
rect 160612 16124 160618 16136
rect 384298 16124 384304 16136
rect 384356 16124 384362 16176
rect 160646 16056 160652 16108
rect 160704 16096 160710 16108
rect 387794 16096 387800 16108
rect 160704 16068 387800 16096
rect 160704 16056 160710 16068
rect 387794 16056 387800 16068
rect 387852 16056 387858 16108
rect 167086 15988 167092 16040
rect 167144 16028 167150 16040
rect 478138 16028 478144 16040
rect 167144 16000 478144 16028
rect 167144 15988 167150 16000
rect 478138 15988 478144 16000
rect 478196 15988 478202 16040
rect 167178 15920 167184 15972
rect 167236 15960 167242 15972
rect 478874 15960 478880 15972
rect 167236 15932 478880 15960
rect 167236 15920 167242 15932
rect 478874 15920 478880 15932
rect 478932 15920 478938 15972
rect 142522 15852 142528 15904
rect 142580 15892 142586 15904
rect 156138 15892 156144 15904
rect 142580 15864 156144 15892
rect 142580 15852 142586 15864
rect 156138 15852 156144 15864
rect 156196 15852 156202 15904
rect 171318 15852 171324 15904
rect 171376 15892 171382 15904
rect 527818 15892 527824 15904
rect 171376 15864 527824 15892
rect 171376 15852 171382 15864
rect 527818 15852 527824 15864
rect 527876 15852 527882 15904
rect 162394 15036 162400 15088
rect 162452 15076 162458 15088
rect 256694 15076 256700 15088
rect 162452 15048 256700 15076
rect 162452 15036 162458 15048
rect 256694 15036 256700 15048
rect 256752 15036 256758 15088
rect 150710 14968 150716 15020
rect 150768 15008 150774 15020
rect 262490 15008 262496 15020
rect 150768 14980 262496 15008
rect 150768 14968 150774 14980
rect 262490 14968 262496 14980
rect 262548 14968 262554 15020
rect 158806 14900 158812 14952
rect 158864 14940 158870 14952
rect 370130 14940 370136 14952
rect 158864 14912 370136 14940
rect 158864 14900 158870 14912
rect 370130 14900 370136 14912
rect 370188 14900 370194 14952
rect 160462 14832 160468 14884
rect 160520 14872 160526 14884
rect 390646 14872 390652 14884
rect 160520 14844 390652 14872
rect 160520 14832 160526 14844
rect 390646 14832 390652 14844
rect 390704 14832 390710 14884
rect 161750 14764 161756 14816
rect 161808 14804 161814 14816
rect 398834 14804 398840 14816
rect 161808 14776 398840 14804
rect 161808 14764 161814 14776
rect 398834 14764 398840 14776
rect 398892 14764 398898 14816
rect 162854 14696 162860 14748
rect 162912 14736 162918 14748
rect 420914 14736 420920 14748
rect 162912 14708 420920 14736
rect 162912 14696 162918 14708
rect 420914 14696 420920 14708
rect 420972 14696 420978 14748
rect 162946 14628 162952 14680
rect 163004 14668 163010 14680
rect 428458 14668 428464 14680
rect 163004 14640 428464 14668
rect 163004 14628 163010 14640
rect 428458 14628 428464 14640
rect 428516 14628 428522 14680
rect 129550 14560 129556 14612
rect 129608 14600 129614 14612
rect 402514 14600 402520 14612
rect 129608 14572 402520 14600
rect 129608 14560 129614 14572
rect 402514 14560 402520 14572
rect 402572 14560 402578 14612
rect 181438 14492 181444 14544
rect 181496 14532 181502 14544
rect 454034 14532 454040 14544
rect 181496 14504 454040 14532
rect 181496 14492 181502 14504
rect 454034 14492 454040 14504
rect 454092 14492 454098 14544
rect 172606 14424 172612 14476
rect 172664 14464 172670 14476
rect 465718 14464 465724 14476
rect 172664 14436 465724 14464
rect 172664 14424 172670 14436
rect 465718 14424 465724 14436
rect 465776 14424 465782 14476
rect 149422 13472 149428 13524
rect 149480 13512 149486 13524
rect 248414 13512 248420 13524
rect 149480 13484 248420 13512
rect 149480 13472 149486 13484
rect 248414 13472 248420 13484
rect 248472 13472 248478 13524
rect 157610 13404 157616 13456
rect 157668 13444 157674 13456
rect 345290 13444 345296 13456
rect 157668 13416 345296 13444
rect 157668 13404 157674 13416
rect 345290 13404 345296 13416
rect 345348 13404 345354 13456
rect 157518 13336 157524 13388
rect 157576 13376 157582 13388
rect 352834 13376 352840 13388
rect 157576 13348 352840 13376
rect 157576 13336 157582 13348
rect 352834 13336 352840 13348
rect 352892 13336 352898 13388
rect 161566 13268 161572 13320
rect 161624 13308 161630 13320
rect 403618 13308 403624 13320
rect 161624 13280 403624 13308
rect 161624 13268 161630 13280
rect 403618 13268 403624 13280
rect 403676 13268 403682 13320
rect 161658 13200 161664 13252
rect 161716 13240 161722 13252
rect 407206 13240 407212 13252
rect 161716 13212 407212 13240
rect 161716 13200 161722 13212
rect 407206 13200 407212 13212
rect 407264 13200 407270 13252
rect 180242 13132 180248 13184
rect 180300 13172 180306 13184
rect 447410 13172 447416 13184
rect 180300 13144 447416 13172
rect 180300 13132 180306 13144
rect 447410 13132 447416 13144
rect 447468 13132 447474 13184
rect 168466 13064 168472 13116
rect 168524 13104 168530 13116
rect 490006 13104 490012 13116
rect 168524 13076 490012 13104
rect 168524 13064 168530 13076
rect 490006 13064 490012 13076
rect 490064 13064 490070 13116
rect 154574 12316 154580 12368
rect 154632 12356 154638 12368
rect 320450 12356 320456 12368
rect 154632 12328 320456 12356
rect 154632 12316 154638 12328
rect 320450 12316 320456 12328
rect 320508 12316 320514 12368
rect 156414 12248 156420 12300
rect 156472 12288 156478 12300
rect 326338 12288 326344 12300
rect 156472 12260 326344 12288
rect 156472 12248 156478 12260
rect 326338 12248 326344 12260
rect 326396 12248 326402 12300
rect 156506 12180 156512 12232
rect 156564 12220 156570 12232
rect 330386 12220 330392 12232
rect 156564 12192 330392 12220
rect 156564 12180 156570 12192
rect 330386 12180 330392 12192
rect 330444 12180 330450 12232
rect 156230 12112 156236 12164
rect 156288 12152 156294 12164
rect 331214 12152 331220 12164
rect 156288 12124 331220 12152
rect 156288 12112 156294 12124
rect 331214 12112 331220 12124
rect 331272 12112 331278 12164
rect 156322 12044 156328 12096
rect 156380 12084 156386 12096
rect 332594 12084 332600 12096
rect 156380 12056 332600 12084
rect 156380 12044 156386 12056
rect 332594 12044 332600 12056
rect 332652 12044 332658 12096
rect 156046 11976 156052 12028
rect 156104 12016 156110 12028
rect 337010 12016 337016 12028
rect 156104 11988 337016 12016
rect 156104 11976 156110 11988
rect 337010 11976 337016 11988
rect 337068 11976 337074 12028
rect 158714 11908 158720 11960
rect 158772 11948 158778 11960
rect 365806 11948 365812 11960
rect 158772 11920 365812 11948
rect 158772 11908 158778 11920
rect 365806 11908 365812 11920
rect 365864 11908 365870 11960
rect 160370 11840 160376 11892
rect 160428 11880 160434 11892
rect 386690 11880 386696 11892
rect 160428 11852 386696 11880
rect 160428 11840 160434 11852
rect 386690 11840 386696 11852
rect 386748 11840 386754 11892
rect 130746 11812 130752 11824
rect 122806 11784 130752 11812
rect 102134 11704 102140 11756
rect 102192 11744 102198 11756
rect 122806 11744 122834 11784
rect 130746 11772 130752 11784
rect 130804 11772 130810 11824
rect 161474 11772 161480 11824
rect 161532 11812 161538 11824
rect 398926 11812 398932 11824
rect 161532 11784 398932 11812
rect 161532 11772 161538 11784
rect 398926 11772 398932 11784
rect 398984 11772 398990 11824
rect 102192 11716 122834 11744
rect 102192 11704 102198 11716
rect 126974 11704 126980 11756
rect 127032 11744 127038 11756
rect 128170 11744 128176 11756
rect 127032 11716 128176 11744
rect 127032 11704 127038 11716
rect 128170 11704 128176 11716
rect 128228 11704 128234 11756
rect 168374 11704 168380 11756
rect 168432 11744 168438 11756
rect 492306 11744 492312 11756
rect 168432 11716 492312 11744
rect 168432 11704 168438 11716
rect 492306 11704 492312 11716
rect 492364 11704 492370 11756
rect 99834 10684 99840 10736
rect 99892 10724 99898 10736
rect 130654 10724 130660 10736
rect 99892 10696 130660 10724
rect 99892 10684 99898 10696
rect 130654 10684 130660 10696
rect 130712 10684 130718 10736
rect 153194 10684 153200 10736
rect 153252 10724 153258 10736
rect 298094 10724 298100 10736
rect 153252 10696 298100 10724
rect 153252 10684 153258 10696
rect 298094 10684 298100 10696
rect 298152 10684 298158 10736
rect 106458 10616 106464 10668
rect 106516 10656 106522 10668
rect 138474 10656 138480 10668
rect 106516 10628 138480 10656
rect 106516 10616 106522 10628
rect 138474 10616 138480 10628
rect 138532 10616 138538 10668
rect 153378 10616 153384 10668
rect 153436 10656 153442 10668
rect 299658 10656 299664 10668
rect 153436 10628 299664 10656
rect 153436 10616 153442 10628
rect 299658 10616 299664 10628
rect 299716 10616 299722 10668
rect 92474 10548 92480 10600
rect 92532 10588 92538 10600
rect 130562 10588 130568 10600
rect 92532 10560 130568 10588
rect 92532 10548 92538 10560
rect 130562 10548 130568 10560
rect 130620 10548 130626 10600
rect 153286 10548 153292 10600
rect 153344 10588 153350 10600
rect 303154 10588 303160 10600
rect 153344 10560 303160 10588
rect 153344 10548 153350 10560
rect 303154 10548 303160 10560
rect 303212 10548 303218 10600
rect 85666 10480 85672 10532
rect 85724 10520 85730 10532
rect 130470 10520 130476 10532
rect 85724 10492 130476 10520
rect 85724 10480 85730 10492
rect 130470 10480 130476 10492
rect 130528 10480 130534 10532
rect 157426 10480 157432 10532
rect 157484 10520 157490 10532
rect 353570 10520 353576 10532
rect 157484 10492 353576 10520
rect 157484 10480 157490 10492
rect 353570 10480 353576 10492
rect 353628 10480 353634 10532
rect 74994 10412 75000 10464
rect 75052 10452 75058 10464
rect 134518 10452 134524 10464
rect 75052 10424 134524 10452
rect 75052 10412 75058 10424
rect 134518 10412 134524 10424
rect 134576 10412 134582 10464
rect 157334 10412 157340 10464
rect 157392 10452 157398 10464
rect 349246 10452 349252 10464
rect 157392 10424 349252 10452
rect 157392 10412 157398 10424
rect 349246 10412 349252 10424
rect 349304 10412 349310 10464
rect 349798 10412 349804 10464
rect 349856 10452 349862 10464
rect 583386 10452 583392 10464
rect 349856 10424 583392 10452
rect 349856 10412 349862 10424
rect 583386 10412 583392 10424
rect 583444 10412 583450 10464
rect 67634 10344 67640 10396
rect 67692 10384 67698 10396
rect 131758 10384 131764 10396
rect 67692 10356 131764 10384
rect 67692 10344 67698 10356
rect 131758 10344 131764 10356
rect 131816 10344 131822 10396
rect 180150 10344 180156 10396
rect 180208 10384 180214 10396
rect 440326 10384 440332 10396
rect 180208 10356 440332 10384
rect 180208 10344 180214 10356
rect 440326 10344 440332 10356
rect 440384 10344 440390 10396
rect 71498 10276 71504 10328
rect 71556 10316 71562 10328
rect 135806 10316 135812 10328
rect 71556 10288 135812 10316
rect 71556 10276 71562 10288
rect 135806 10276 135812 10288
rect 135864 10276 135870 10328
rect 166074 10276 166080 10328
rect 166132 10316 166138 10328
rect 456886 10316 456892 10328
rect 166132 10288 456892 10316
rect 166132 10276 166138 10288
rect 456886 10276 456892 10288
rect 456944 10276 456950 10328
rect 151814 9596 151820 9648
rect 151872 9636 151878 9648
rect 281902 9636 281908 9648
rect 151872 9608 281908 9636
rect 151872 9596 151878 9608
rect 281902 9596 281908 9608
rect 281960 9596 281966 9648
rect 151906 9528 151912 9580
rect 151964 9568 151970 9580
rect 285398 9568 285404 9580
rect 151964 9540 285404 9568
rect 151964 9528 151970 9540
rect 285398 9528 285404 9540
rect 285456 9528 285462 9580
rect 155954 9460 155960 9512
rect 156012 9500 156018 9512
rect 332686 9500 332692 9512
rect 156012 9472 332692 9500
rect 156012 9460 156018 9472
rect 332686 9460 332692 9472
rect 332744 9460 332750 9512
rect 156966 9392 156972 9444
rect 157024 9432 157030 9444
rect 336274 9432 336280 9444
rect 157024 9404 336280 9432
rect 157024 9392 157030 9404
rect 336274 9392 336280 9404
rect 336332 9392 336338 9444
rect 160186 9324 160192 9376
rect 160244 9364 160250 9376
rect 382366 9364 382372 9376
rect 160244 9336 382372 9364
rect 160244 9324 160250 9336
rect 382366 9324 382372 9336
rect 382424 9324 382430 9376
rect 160278 9256 160284 9308
rect 160336 9296 160342 9308
rect 385954 9296 385960 9308
rect 160336 9268 385960 9296
rect 160336 9256 160342 9268
rect 385954 9256 385960 9268
rect 386012 9256 386018 9308
rect 160094 9188 160100 9240
rect 160152 9228 160158 9240
rect 389450 9228 389456 9240
rect 160152 9200 389456 9228
rect 160152 9188 160158 9200
rect 389450 9188 389456 9200
rect 389508 9188 389514 9240
rect 57238 9120 57244 9172
rect 57296 9160 57302 9172
rect 134334 9160 134340 9172
rect 57296 9132 134340 9160
rect 57296 9120 57302 9132
rect 134334 9120 134340 9132
rect 134392 9120 134398 9172
rect 164326 9120 164332 9172
rect 164384 9160 164390 9172
rect 436738 9160 436744 9172
rect 164384 9132 436744 9160
rect 164384 9120 164390 9132
rect 436738 9120 436744 9132
rect 436796 9120 436802 9172
rect 53742 9052 53748 9104
rect 53800 9092 53806 9104
rect 134242 9092 134248 9104
rect 53800 9064 134248 9092
rect 53800 9052 53806 9064
rect 134242 9052 134248 9064
rect 134300 9052 134306 9104
rect 165982 9052 165988 9104
rect 166040 9092 166046 9104
rect 453298 9092 453304 9104
rect 166040 9064 453304 9092
rect 166040 9052 166046 9064
rect 453298 9052 453304 9064
rect 453356 9052 453362 9104
rect 50154 8984 50160 9036
rect 50212 9024 50218 9036
rect 134150 9024 134156 9036
rect 50212 8996 134156 9024
rect 50212 8984 50218 8996
rect 134150 8984 134156 8996
rect 134208 8984 134214 9036
rect 165890 8984 165896 9036
rect 165948 9024 165954 9036
rect 459186 9024 459192 9036
rect 165948 8996 459192 9024
rect 165948 8984 165954 8996
rect 459186 8984 459192 8996
rect 459244 8984 459250 9036
rect 38378 8916 38384 8968
rect 38436 8956 38442 8968
rect 132954 8956 132960 8968
rect 38436 8928 132960 8956
rect 38436 8916 38442 8928
rect 132954 8916 132960 8928
rect 133012 8916 133018 8968
rect 171226 8916 171232 8968
rect 171284 8956 171290 8968
rect 525426 8956 525432 8968
rect 171284 8928 525432 8956
rect 171284 8916 171290 8928
rect 525426 8916 525432 8928
rect 525484 8916 525490 8968
rect 150618 8848 150624 8900
rect 150676 8888 150682 8900
rect 264146 8888 264152 8900
rect 150676 8860 264152 8888
rect 150676 8848 150682 8860
rect 264146 8848 264152 8860
rect 264204 8848 264210 8900
rect 150526 8780 150532 8832
rect 150584 8820 150590 8832
rect 258258 8820 258264 8832
rect 150584 8792 258264 8820
rect 150584 8780 150590 8792
rect 258258 8780 258264 8792
rect 258316 8780 258322 8832
rect 177482 8712 177488 8764
rect 177540 8752 177546 8764
rect 267734 8752 267740 8764
rect 177540 8724 267740 8752
rect 177540 8712 177546 8724
rect 267734 8712 267740 8724
rect 267792 8712 267798 8764
rect 123478 8032 123484 8084
rect 123536 8072 123542 8084
rect 139578 8072 139584 8084
rect 123536 8044 139584 8072
rect 123536 8032 123542 8044
rect 139578 8032 139584 8044
rect 139636 8032 139642 8084
rect 110506 7964 110512 8016
rect 110564 8004 110570 8016
rect 129090 8004 129096 8016
rect 110564 7976 129096 8004
rect 110564 7964 110570 7976
rect 129090 7964 129096 7976
rect 129148 7964 129154 8016
rect 111610 7896 111616 7948
rect 111668 7936 111674 7948
rect 138290 7936 138296 7948
rect 111668 7908 138296 7936
rect 111668 7896 111674 7908
rect 138290 7896 138296 7908
rect 138348 7896 138354 7948
rect 109310 7828 109316 7880
rect 109368 7868 109374 7880
rect 138382 7868 138388 7880
rect 109368 7840 138388 7868
rect 109368 7828 109374 7840
rect 138382 7828 138388 7840
rect 138440 7828 138446 7880
rect 337378 7828 337384 7880
rect 337436 7868 337442 7880
rect 580994 7868 581000 7880
rect 337436 7840 581000 7868
rect 337436 7828 337442 7840
rect 580994 7828 581000 7840
rect 581052 7828 581058 7880
rect 102226 7760 102232 7812
rect 102284 7800 102290 7812
rect 138198 7800 138204 7812
rect 102284 7772 138204 7800
rect 102284 7760 102290 7772
rect 138198 7760 138204 7772
rect 138256 7760 138262 7812
rect 176102 7760 176108 7812
rect 176160 7800 176166 7812
rect 426158 7800 426164 7812
rect 176160 7772 426164 7800
rect 176160 7760 176166 7772
rect 426158 7760 426164 7772
rect 426216 7760 426222 7812
rect 95142 7692 95148 7744
rect 95200 7732 95206 7744
rect 137094 7732 137100 7744
rect 95200 7704 137100 7732
rect 95200 7692 95206 7704
rect 137094 7692 137100 7704
rect 137152 7692 137158 7744
rect 165798 7692 165804 7744
rect 165856 7732 165862 7744
rect 455690 7732 455696 7744
rect 165856 7704 455696 7732
rect 165856 7692 165862 7704
rect 455690 7692 455696 7704
rect 455748 7692 455754 7744
rect 66714 7624 66720 7676
rect 66772 7664 66778 7676
rect 135714 7664 135720 7676
rect 66772 7636 135720 7664
rect 66772 7624 66778 7636
rect 135714 7624 135720 7636
rect 135772 7624 135778 7676
rect 169846 7624 169852 7676
rect 169904 7664 169910 7676
rect 469950 7664 469956 7676
rect 169904 7636 469956 7664
rect 169904 7624 169910 7636
rect 469950 7624 469956 7636
rect 470008 7624 470014 7676
rect 31294 7556 31300 7608
rect 31352 7596 31358 7608
rect 132862 7596 132868 7608
rect 31352 7568 132868 7596
rect 31352 7556 31358 7568
rect 132862 7556 132868 7568
rect 132920 7556 132926 7608
rect 166994 7556 167000 7608
rect 167052 7596 167058 7608
rect 471054 7596 471060 7608
rect 167052 7568 471060 7596
rect 167052 7556 167058 7568
rect 471054 7556 471060 7568
rect 471112 7556 471118 7608
rect 129642 6740 129648 6792
rect 129700 6780 129706 6792
rect 189718 6780 189724 6792
rect 129700 6752 189724 6780
rect 129700 6740 129706 6752
rect 189718 6740 189724 6752
rect 189776 6740 189782 6792
rect 92566 6672 92572 6724
rect 92624 6712 92630 6724
rect 132770 6712 132776 6724
rect 92624 6684 132776 6712
rect 92624 6672 92630 6684
rect 132770 6672 132776 6684
rect 132828 6672 132834 6724
rect 147858 6672 147864 6724
rect 147916 6712 147922 6724
rect 228726 6712 228732 6724
rect 147916 6684 228732 6712
rect 147916 6672 147922 6684
rect 228726 6672 228732 6684
rect 228784 6672 228790 6724
rect 87966 6604 87972 6656
rect 88024 6644 88030 6656
rect 137002 6644 137008 6656
rect 88024 6616 137008 6644
rect 88024 6604 88030 6616
rect 137002 6604 137008 6616
rect 137060 6604 137066 6656
rect 149238 6604 149244 6656
rect 149296 6644 149302 6656
rect 239306 6644 239312 6656
rect 149296 6616 239312 6644
rect 149296 6604 149302 6616
rect 239306 6604 239312 6616
rect 239364 6604 239370 6656
rect 77386 6536 77392 6588
rect 77444 6576 77450 6588
rect 135530 6576 135536 6588
rect 77444 6548 135536 6576
rect 77444 6536 77450 6548
rect 135530 6536 135536 6548
rect 135588 6536 135594 6588
rect 149146 6536 149152 6588
rect 149204 6576 149210 6588
rect 242986 6576 242992 6588
rect 149204 6548 242992 6576
rect 149204 6536 149210 6548
rect 242986 6536 242992 6548
rect 243044 6536 243050 6588
rect 73798 6468 73804 6520
rect 73856 6508 73862 6520
rect 135438 6508 135444 6520
rect 73856 6480 135444 6508
rect 73856 6468 73862 6480
rect 135438 6468 135444 6480
rect 135496 6468 135502 6520
rect 149054 6468 149060 6520
rect 149112 6508 149118 6520
rect 246390 6508 246396 6520
rect 149112 6480 246396 6508
rect 149112 6468 149118 6480
rect 246390 6468 246396 6480
rect 246448 6468 246454 6520
rect 56042 6400 56048 6452
rect 56100 6440 56106 6452
rect 134058 6440 134064 6452
rect 56100 6412 134064 6440
rect 56100 6400 56106 6412
rect 134058 6400 134064 6412
rect 134116 6400 134122 6452
rect 149330 6400 149336 6452
rect 149388 6440 149394 6452
rect 249978 6440 249984 6452
rect 149388 6412 249984 6440
rect 149388 6400 149394 6412
rect 249978 6400 249984 6412
rect 250036 6400 250042 6452
rect 52546 6332 52552 6384
rect 52604 6372 52610 6384
rect 134702 6372 134708 6384
rect 52604 6344 134708 6372
rect 52604 6332 52610 6344
rect 134702 6332 134708 6344
rect 134760 6332 134766 6384
rect 150434 6332 150440 6384
rect 150492 6372 150498 6384
rect 260650 6372 260656 6384
rect 150492 6344 260656 6372
rect 150492 6332 150498 6344
rect 260650 6332 260656 6344
rect 260708 6332 260714 6384
rect 40678 6264 40684 6316
rect 40736 6304 40742 6316
rect 132678 6304 132684 6316
rect 40736 6276 132684 6304
rect 40736 6264 40742 6276
rect 132678 6264 132684 6276
rect 132736 6264 132742 6316
rect 165706 6264 165712 6316
rect 165764 6304 165770 6316
rect 450906 6304 450912 6316
rect 165764 6276 450912 6304
rect 165764 6264 165770 6276
rect 450906 6264 450912 6276
rect 450964 6264 450970 6316
rect 24210 6196 24216 6248
rect 24268 6236 24274 6248
rect 131574 6236 131580 6248
rect 24268 6208 131580 6236
rect 24268 6196 24274 6208
rect 131574 6196 131580 6208
rect 131632 6196 131638 6248
rect 142430 6196 142436 6248
rect 142488 6236 142494 6248
rect 155402 6236 155408 6248
rect 142488 6208 155408 6236
rect 142488 6196 142494 6208
rect 155402 6196 155408 6208
rect 155460 6196 155466 6248
rect 165614 6196 165620 6248
rect 165672 6236 165678 6248
rect 460382 6236 460388 6248
rect 165672 6208 460388 6236
rect 165672 6196 165678 6208
rect 460382 6196 460388 6208
rect 460440 6196 460446 6248
rect 23014 6128 23020 6180
rect 23072 6168 23078 6180
rect 131482 6168 131488 6180
rect 23072 6140 131488 6168
rect 23072 6128 23078 6140
rect 131482 6128 131488 6140
rect 131540 6128 131546 6180
rect 143994 6128 144000 6180
rect 144052 6168 144058 6180
rect 170766 6168 170772 6180
rect 144052 6140 170772 6168
rect 144052 6128 144058 6140
rect 170766 6128 170772 6140
rect 170824 6128 170830 6180
rect 176562 6128 176568 6180
rect 176620 6168 176626 6180
rect 578602 6168 578608 6180
rect 176620 6140 578608 6168
rect 176620 6128 176626 6140
rect 578602 6128 578608 6140
rect 578660 6128 578666 6180
rect 126882 5380 126888 5432
rect 126940 5420 126946 5432
rect 133322 5420 133328 5432
rect 126940 5392 133328 5420
rect 126940 5380 126946 5392
rect 133322 5380 133328 5392
rect 133380 5380 133386 5432
rect 104526 5176 104532 5228
rect 104584 5216 104590 5228
rect 139026 5216 139032 5228
rect 104584 5188 139032 5216
rect 104584 5176 104590 5188
rect 139026 5176 139032 5188
rect 139084 5176 139090 5228
rect 143810 5176 143816 5228
rect 143868 5216 143874 5228
rect 173158 5216 173164 5228
rect 143868 5188 173164 5216
rect 143868 5176 143874 5188
rect 173158 5176 173164 5188
rect 173216 5176 173222 5228
rect 20622 5108 20628 5160
rect 20680 5148 20686 5160
rect 43438 5148 43444 5160
rect 20680 5120 43444 5148
rect 20680 5108 20686 5120
rect 43438 5108 43444 5120
rect 43496 5108 43502 5160
rect 70302 5108 70308 5160
rect 70360 5148 70366 5160
rect 136082 5148 136088 5160
rect 70360 5120 136088 5148
rect 70360 5108 70366 5120
rect 136082 5108 136088 5120
rect 136140 5108 136146 5160
rect 143718 5108 143724 5160
rect 143776 5148 143782 5160
rect 174262 5148 174268 5160
rect 143776 5120 174268 5148
rect 143776 5108 143782 5120
rect 174262 5108 174268 5120
rect 174320 5108 174326 5160
rect 431218 5108 431224 5160
rect 431276 5148 431282 5160
rect 475746 5148 475752 5160
rect 431276 5120 475752 5148
rect 431276 5108 431282 5120
rect 475746 5108 475752 5120
rect 475804 5108 475810 5160
rect 28902 5040 28908 5092
rect 28960 5080 28966 5092
rect 126238 5080 126244 5092
rect 28960 5052 126244 5080
rect 28960 5040 28966 5052
rect 126238 5040 126244 5052
rect 126296 5040 126302 5092
rect 164234 5040 164240 5092
rect 164292 5080 164298 5092
rect 443822 5080 443828 5092
rect 164292 5052 443828 5080
rect 164292 5040 164298 5052
rect 443822 5040 443828 5052
rect 443880 5040 443886 5092
rect 33594 4972 33600 5024
rect 33652 5012 33658 5024
rect 133138 5012 133144 5024
rect 33652 4984 133144 5012
rect 33652 4972 33658 4984
rect 133138 4972 133144 4984
rect 133196 4972 133202 5024
rect 142338 4972 142344 5024
rect 142396 5012 142402 5024
rect 151814 5012 151820 5024
rect 142396 4984 151820 5012
rect 142396 4972 142402 4984
rect 151814 4972 151820 4984
rect 151872 4972 151878 5024
rect 170858 4972 170864 5024
rect 170916 5012 170922 5024
rect 508866 5012 508872 5024
rect 170916 4984 508872 5012
rect 170916 4972 170922 4984
rect 508866 4972 508872 4984
rect 508924 4972 508930 5024
rect 21818 4904 21824 4956
rect 21876 4944 21882 4956
rect 131390 4944 131396 4956
rect 21876 4916 131396 4944
rect 21876 4904 21882 4916
rect 131390 4904 131396 4916
rect 131448 4904 131454 4956
rect 142246 4904 142252 4956
rect 142304 4944 142310 4956
rect 157794 4944 157800 4956
rect 142304 4916 157800 4944
rect 142304 4904 142310 4916
rect 157794 4904 157800 4916
rect 157852 4904 157858 4956
rect 171134 4904 171140 4956
rect 171192 4944 171198 4956
rect 533706 4944 533712 4956
rect 171192 4916 533712 4944
rect 171192 4904 171198 4916
rect 533706 4904 533712 4916
rect 533764 4904 533770 4956
rect 14734 4836 14740 4888
rect 14792 4876 14798 4888
rect 131298 4876 131304 4888
rect 14792 4848 131304 4876
rect 14792 4836 14798 4848
rect 131298 4836 131304 4848
rect 131356 4836 131362 4888
rect 143626 4836 143632 4888
rect 143684 4876 143690 4888
rect 167178 4876 167184 4888
rect 143684 4848 167184 4876
rect 143684 4836 143690 4848
rect 167178 4836 167184 4848
rect 167236 4836 167242 4888
rect 173618 4836 173624 4888
rect 173676 4876 173682 4888
rect 551462 4876 551468 4888
rect 173676 4848 551468 4876
rect 173676 4836 173682 4848
rect 551462 4836 551468 4848
rect 551520 4836 551526 4888
rect 13538 4768 13544 4820
rect 13596 4808 13602 4820
rect 131206 4808 131212 4820
rect 13596 4780 131212 4808
rect 13596 4768 13602 4780
rect 131206 4768 131212 4780
rect 131264 4768 131270 4820
rect 143902 4768 143908 4820
rect 143960 4808 143966 4820
rect 169570 4808 169576 4820
rect 143960 4780 169576 4808
rect 143960 4768 143966 4780
rect 169570 4768 169576 4780
rect 169628 4768 169634 4820
rect 174906 4768 174912 4820
rect 174964 4808 174970 4820
rect 566826 4808 566832 4820
rect 174964 4780 566832 4808
rect 174964 4768 174970 4780
rect 566826 4768 566832 4780
rect 566884 4768 566890 4820
rect 201420 4168 202828 4196
rect 18230 4088 18236 4140
rect 18288 4128 18294 4140
rect 131942 4128 131948 4140
rect 18288 4100 131948 4128
rect 18288 4088 18294 4100
rect 131942 4088 131948 4100
rect 132000 4088 132006 4140
rect 140958 4088 140964 4140
rect 141016 4128 141022 4140
rect 144730 4128 144736 4140
rect 141016 4100 144736 4128
rect 141016 4088 141022 4100
rect 144730 4088 144736 4100
rect 144788 4088 144794 4140
rect 146294 4088 146300 4140
rect 146352 4128 146358 4140
rect 201420 4128 201448 4168
rect 146352 4100 201448 4128
rect 146352 4088 146358 4100
rect 201494 4088 201500 4140
rect 201552 4128 201558 4140
rect 202690 4128 202696 4140
rect 201552 4100 202696 4128
rect 201552 4088 201558 4100
rect 202690 4088 202696 4100
rect 202748 4088 202754 4140
rect 202800 4128 202828 4168
rect 207382 4128 207388 4140
rect 202800 4100 207388 4128
rect 207382 4088 207388 4100
rect 207440 4088 207446 4140
rect 125870 4020 125876 4072
rect 125928 4060 125934 4072
rect 139946 4060 139952 4072
rect 125928 4032 139952 4060
rect 125928 4020 125934 4032
rect 139946 4020 139952 4032
rect 140004 4020 140010 4072
rect 146386 4020 146392 4072
rect 146444 4060 146450 4072
rect 210970 4060 210976 4072
rect 146444 4032 210976 4060
rect 146444 4020 146450 4032
rect 210970 4020 210976 4032
rect 211028 4020 211034 4072
rect 90358 3952 90364 4004
rect 90416 3992 90422 4004
rect 137370 3992 137376 4004
rect 90416 3964 137376 3992
rect 90416 3952 90422 3964
rect 137370 3952 137376 3964
rect 137428 3952 137434 4004
rect 147766 3952 147772 4004
rect 147824 3992 147830 4004
rect 221550 3992 221556 4004
rect 147824 3964 221556 3992
rect 147824 3952 147830 3964
rect 221550 3952 221556 3964
rect 221608 3952 221614 4004
rect 251174 3952 251180 4004
rect 251232 3992 251238 4004
rect 252370 3992 252376 4004
rect 251232 3964 252376 3992
rect 251232 3952 251238 3964
rect 252370 3952 252376 3964
rect 252428 3952 252434 4004
rect 86862 3884 86868 3936
rect 86920 3924 86926 3936
rect 137278 3924 137284 3936
rect 86920 3896 137284 3924
rect 86920 3884 86926 3896
rect 137278 3884 137284 3896
rect 137336 3884 137342 3936
rect 170674 3884 170680 3936
rect 170732 3924 170738 3936
rect 349154 3924 349160 3936
rect 170732 3896 349160 3924
rect 170732 3884 170738 3896
rect 349154 3884 349160 3896
rect 349212 3884 349218 3936
rect 349890 3884 349896 3936
rect 349948 3924 349954 3936
rect 545482 3924 545488 3936
rect 349948 3896 545488 3924
rect 349948 3884 349954 3896
rect 545482 3884 545488 3896
rect 545540 3884 545546 3936
rect 72602 3816 72608 3868
rect 72660 3856 72666 3868
rect 130378 3856 130384 3868
rect 72660 3828 130384 3856
rect 72660 3816 72666 3828
rect 130378 3816 130384 3828
rect 130436 3816 130442 3868
rect 141050 3816 141056 3868
rect 141108 3856 141114 3868
rect 147122 3856 147128 3868
rect 141108 3828 147128 3856
rect 141108 3816 141114 3828
rect 147122 3816 147128 3828
rect 147180 3816 147186 3868
rect 148594 3816 148600 3868
rect 148652 3856 148658 3868
rect 225138 3856 225144 3868
rect 148652 3828 225144 3856
rect 148652 3816 148658 3828
rect 225138 3816 225144 3828
rect 225196 3816 225202 3868
rect 228358 3816 228364 3868
rect 228416 3856 228422 3868
rect 469858 3856 469864 3868
rect 228416 3828 469864 3856
rect 228416 3816 228422 3828
rect 469858 3816 469864 3828
rect 469916 3816 469922 3868
rect 469950 3816 469956 3868
rect 470008 3856 470014 3868
rect 504174 3856 504180 3868
rect 470008 3828 504180 3856
rect 470008 3816 470014 3828
rect 504174 3816 504180 3828
rect 504232 3816 504238 3868
rect 76190 3748 76196 3800
rect 76248 3788 76254 3800
rect 135990 3788 135996 3800
rect 76248 3760 135996 3788
rect 76248 3748 76254 3760
rect 135990 3748 135996 3760
rect 136048 3748 136054 3800
rect 142154 3748 142160 3800
rect 142212 3788 142218 3800
rect 154206 3788 154212 3800
rect 142212 3760 154212 3788
rect 142212 3748 142218 3760
rect 154206 3748 154212 3760
rect 154264 3748 154270 3800
rect 159358 3748 159364 3800
rect 159416 3788 159422 3800
rect 180242 3788 180248 3800
rect 159416 3760 180248 3788
rect 159416 3748 159422 3760
rect 180242 3748 180248 3760
rect 180300 3748 180306 3800
rect 185578 3748 185584 3800
rect 185636 3788 185642 3800
rect 472250 3788 472256 3800
rect 185636 3760 472256 3788
rect 185636 3748 185642 3760
rect 472250 3748 472256 3760
rect 472308 3748 472314 3800
rect 32398 3680 32404 3732
rect 32456 3720 32462 3732
rect 92566 3720 92572 3732
rect 32456 3692 92572 3720
rect 32456 3680 32462 3692
rect 92566 3680 92572 3692
rect 92624 3680 92630 3732
rect 93946 3680 93952 3732
rect 94004 3720 94010 3732
rect 136818 3720 136824 3732
rect 94004 3692 136824 3720
rect 94004 3680 94010 3692
rect 136818 3680 136824 3692
rect 136876 3680 136882 3732
rect 141234 3680 141240 3732
rect 141292 3720 141298 3732
rect 142430 3720 142436 3732
rect 141292 3692 142436 3720
rect 141292 3680 141298 3692
rect 142430 3680 142436 3692
rect 142488 3680 142494 3732
rect 144454 3680 144460 3732
rect 144512 3720 144518 3732
rect 160094 3720 160100 3732
rect 144512 3692 160100 3720
rect 144512 3680 144518 3692
rect 160094 3680 160100 3692
rect 160152 3680 160158 3732
rect 176010 3680 176016 3732
rect 176068 3720 176074 3732
rect 465166 3720 465172 3732
rect 176068 3692 465172 3720
rect 176068 3680 176074 3692
rect 465166 3680 465172 3692
rect 465224 3680 465230 3732
rect 465718 3680 465724 3732
rect 465776 3720 465782 3732
rect 549070 3720 549076 3732
rect 465776 3692 549076 3720
rect 465776 3680 465782 3692
rect 549070 3680 549076 3692
rect 549128 3680 549134 3732
rect 59630 3612 59636 3664
rect 59688 3652 59694 3664
rect 120718 3652 120724 3664
rect 59688 3624 120724 3652
rect 59688 3612 59694 3624
rect 120718 3612 120724 3624
rect 120776 3612 120782 3664
rect 144178 3612 144184 3664
rect 144236 3652 144242 3664
rect 164878 3652 164884 3664
rect 144236 3624 164884 3652
rect 144236 3612 144242 3624
rect 164878 3612 164884 3624
rect 164936 3612 164942 3664
rect 177390 3612 177396 3664
rect 177448 3652 177454 3664
rect 494698 3652 494704 3664
rect 177448 3624 494704 3652
rect 177448 3612 177454 3624
rect 494698 3612 494704 3624
rect 494756 3612 494762 3664
rect 46658 3544 46664 3596
rect 46716 3584 46722 3596
rect 128998 3584 129004 3596
rect 46716 3556 129004 3584
rect 46716 3544 46722 3556
rect 128998 3544 129004 3556
rect 129056 3544 129062 3596
rect 136450 3544 136456 3596
rect 136508 3584 136514 3596
rect 140222 3584 140228 3596
rect 136508 3556 140228 3584
rect 136508 3544 136514 3556
rect 140222 3544 140228 3556
rect 140280 3544 140286 3596
rect 141602 3544 141608 3596
rect 141660 3584 141666 3596
rect 143534 3584 143540 3596
rect 141660 3556 143540 3584
rect 141660 3544 141666 3556
rect 143534 3544 143540 3556
rect 143592 3544 143598 3596
rect 146018 3544 146024 3596
rect 146076 3584 146082 3596
rect 146076 3556 149652 3584
rect 146076 3544 146082 3556
rect 2774 3476 2780 3528
rect 2832 3516 2838 3528
rect 3694 3516 3700 3528
rect 2832 3488 3700 3516
rect 2832 3476 2838 3488
rect 3694 3476 3700 3488
rect 3752 3476 3758 3528
rect 11146 3476 11152 3528
rect 11204 3516 11210 3528
rect 13078 3516 13084 3528
rect 11204 3488 13084 3516
rect 11204 3476 11210 3488
rect 13078 3476 13084 3488
rect 13136 3476 13142 3528
rect 37182 3476 37188 3528
rect 37240 3516 37246 3528
rect 126882 3516 126888 3528
rect 37240 3488 126888 3516
rect 37240 3476 37246 3488
rect 126882 3476 126888 3488
rect 126940 3476 126946 3528
rect 140038 3476 140044 3528
rect 140096 3516 140102 3528
rect 141142 3516 141148 3528
rect 140096 3488 141148 3516
rect 140096 3476 140102 3488
rect 141142 3476 141148 3488
rect 141200 3476 141206 3528
rect 144270 3476 144276 3528
rect 144328 3516 144334 3528
rect 149514 3516 149520 3528
rect 144328 3488 149520 3516
rect 144328 3476 144334 3488
rect 149514 3476 149520 3488
rect 149572 3476 149578 3528
rect 149624 3516 149652 3556
rect 151078 3544 151084 3596
rect 151136 3584 151142 3596
rect 153010 3584 153016 3596
rect 151136 3556 153016 3584
rect 151136 3544 151142 3556
rect 153010 3544 153016 3556
rect 153068 3544 153074 3596
rect 156414 3544 156420 3596
rect 156472 3584 156478 3596
rect 171962 3584 171968 3596
rect 156472 3556 171968 3584
rect 156472 3544 156478 3556
rect 171962 3544 171968 3556
rect 172020 3544 172026 3596
rect 177298 3544 177304 3596
rect 177356 3584 177362 3596
rect 505370 3584 505376 3596
rect 177356 3556 505376 3584
rect 177356 3544 177362 3556
rect 505370 3544 505376 3556
rect 505428 3544 505434 3596
rect 168374 3516 168380 3528
rect 149624 3488 168380 3516
rect 168374 3476 168380 3488
rect 168432 3476 168438 3528
rect 170398 3476 170404 3528
rect 170456 3516 170462 3528
rect 501782 3516 501788 3528
rect 170456 3488 501788 3516
rect 170456 3476 170462 3488
rect 501782 3476 501788 3488
rect 501840 3476 501846 3528
rect 506474 3476 506480 3528
rect 506532 3516 506538 3528
rect 507302 3516 507308 3528
rect 506532 3488 507308 3516
rect 506532 3476 506538 3488
rect 507302 3476 507308 3488
rect 507360 3476 507366 3528
rect 531314 3476 531320 3528
rect 531372 3516 531378 3528
rect 532142 3516 532148 3528
rect 531372 3488 532148 3516
rect 531372 3476 531378 3488
rect 532142 3476 532148 3488
rect 532200 3476 532206 3528
rect 539594 3476 539600 3528
rect 539652 3516 539658 3528
rect 540422 3516 540428 3528
rect 539652 3488 540428 3516
rect 539652 3476 539658 3488
rect 540422 3476 540428 3488
rect 540480 3476 540486 3528
rect 564434 3476 564440 3528
rect 564492 3516 564498 3528
rect 565262 3516 565268 3528
rect 564492 3488 565268 3516
rect 564492 3476 564498 3488
rect 565262 3476 565268 3488
rect 565320 3476 565326 3528
rect 5258 3408 5264 3460
rect 5316 3448 5322 3460
rect 10318 3448 10324 3460
rect 5316 3420 10324 3448
rect 5316 3408 5322 3420
rect 10318 3408 10324 3420
rect 10376 3408 10382 3460
rect 102134 3408 102140 3460
rect 102192 3448 102198 3460
rect 103330 3448 103336 3460
rect 102192 3420 103336 3448
rect 102192 3408 102198 3420
rect 103330 3408 103336 3420
rect 103388 3408 103394 3460
rect 131758 3408 131764 3460
rect 131816 3448 131822 3460
rect 139946 3448 139952 3460
rect 131816 3420 139952 3448
rect 131816 3408 131822 3420
rect 139946 3408 139952 3420
rect 140004 3408 140010 3460
rect 144546 3408 144552 3460
rect 144604 3448 144610 3460
rect 176654 3448 176660 3460
rect 144604 3420 176660 3448
rect 144604 3408 144610 3420
rect 176654 3408 176660 3420
rect 176712 3408 176718 3460
rect 177942 3408 177948 3460
rect 178000 3448 178006 3460
rect 523034 3448 523040 3460
rect 178000 3420 523040 3448
rect 178000 3408 178006 3420
rect 523034 3408 523040 3420
rect 523092 3408 523098 3460
rect 122282 3340 122288 3392
rect 122340 3380 122346 3392
rect 139762 3380 139768 3392
rect 122340 3352 139768 3380
rect 122340 3340 122346 3352
rect 139762 3340 139768 3352
rect 139820 3340 139826 3392
rect 145650 3340 145656 3392
rect 145708 3380 145714 3392
rect 145708 3352 146156 3380
rect 145708 3340 145714 3352
rect 142890 3272 142896 3324
rect 142948 3312 142954 3324
rect 145926 3312 145932 3324
rect 142948 3284 145932 3312
rect 142948 3272 142954 3284
rect 145926 3272 145932 3284
rect 145984 3272 145990 3324
rect 146128 3312 146156 3352
rect 151262 3340 151268 3392
rect 151320 3380 151326 3392
rect 203886 3380 203892 3392
rect 151320 3352 203892 3380
rect 151320 3340 151326 3352
rect 203886 3340 203892 3352
rect 203944 3340 203950 3392
rect 242894 3340 242900 3392
rect 242952 3380 242958 3392
rect 244090 3380 244096 3392
rect 242952 3352 244096 3380
rect 242952 3340 242958 3352
rect 244090 3340 244096 3352
rect 244148 3340 244154 3392
rect 299474 3340 299480 3392
rect 299532 3380 299538 3392
rect 300762 3380 300768 3392
rect 299532 3352 300768 3380
rect 299532 3340 299538 3352
rect 300762 3340 300768 3352
rect 300820 3340 300826 3392
rect 307754 3340 307760 3392
rect 307812 3380 307818 3392
rect 309042 3380 309048 3392
rect 307812 3352 309048 3380
rect 307812 3340 307818 3352
rect 309042 3340 309048 3352
rect 309100 3340 309106 3392
rect 316034 3340 316040 3392
rect 316092 3380 316098 3392
rect 317322 3380 317328 3392
rect 316092 3352 317328 3380
rect 316092 3340 316098 3352
rect 317322 3340 317328 3352
rect 317380 3340 317386 3392
rect 324314 3340 324320 3392
rect 324372 3380 324378 3392
rect 325602 3380 325608 3392
rect 324372 3352 325608 3380
rect 324372 3340 324378 3352
rect 325602 3340 325608 3352
rect 325660 3340 325666 3392
rect 332594 3340 332600 3392
rect 332652 3380 332658 3392
rect 333882 3380 333888 3392
rect 332652 3352 333888 3380
rect 332652 3340 332658 3352
rect 333882 3340 333888 3352
rect 333940 3340 333946 3392
rect 340874 3340 340880 3392
rect 340932 3380 340938 3392
rect 342162 3380 342168 3392
rect 340932 3352 342168 3380
rect 340932 3340 340938 3352
rect 342162 3340 342168 3352
rect 342220 3340 342226 3392
rect 349246 3340 349252 3392
rect 349304 3380 349310 3392
rect 350442 3380 350448 3392
rect 349304 3352 350448 3380
rect 349304 3340 349310 3352
rect 350442 3340 350448 3352
rect 350500 3340 350506 3392
rect 357434 3340 357440 3392
rect 357492 3380 357498 3392
rect 358722 3380 358728 3392
rect 357492 3352 358728 3380
rect 357492 3340 357498 3352
rect 358722 3340 358728 3352
rect 358780 3340 358786 3392
rect 374086 3340 374092 3392
rect 374144 3380 374150 3392
rect 375282 3380 375288 3392
rect 374144 3352 375288 3380
rect 374144 3340 374150 3352
rect 375282 3340 375288 3352
rect 375340 3340 375346 3392
rect 382274 3340 382280 3392
rect 382332 3380 382338 3392
rect 383562 3380 383568 3392
rect 382332 3352 383568 3380
rect 382332 3340 382338 3352
rect 383562 3340 383568 3352
rect 383620 3340 383626 3392
rect 390554 3340 390560 3392
rect 390612 3380 390618 3392
rect 391842 3380 391848 3392
rect 390612 3352 391848 3380
rect 390612 3340 390618 3352
rect 391842 3340 391848 3352
rect 391900 3340 391906 3392
rect 398926 3340 398932 3392
rect 398984 3380 398990 3392
rect 400122 3380 400128 3392
rect 398984 3352 400128 3380
rect 398984 3340 398990 3352
rect 400122 3340 400128 3352
rect 400180 3340 400186 3392
rect 407114 3340 407120 3392
rect 407172 3380 407178 3392
rect 408402 3380 408408 3392
rect 407172 3352 408408 3380
rect 407172 3340 407178 3352
rect 408402 3340 408408 3352
rect 408460 3340 408466 3392
rect 415394 3340 415400 3392
rect 415452 3380 415458 3392
rect 416682 3380 416688 3392
rect 415452 3352 416688 3380
rect 415452 3340 415458 3352
rect 416682 3340 416688 3352
rect 416740 3340 416746 3392
rect 423766 3340 423772 3392
rect 423824 3380 423830 3392
rect 424962 3380 424968 3392
rect 423824 3352 424968 3380
rect 423824 3340 423830 3352
rect 424962 3340 424968 3352
rect 425020 3340 425026 3392
rect 432046 3340 432052 3392
rect 432104 3380 432110 3392
rect 433242 3380 433248 3392
rect 432104 3352 433248 3380
rect 432104 3340 432110 3352
rect 433242 3340 433248 3352
rect 433300 3340 433306 3392
rect 456794 3340 456800 3392
rect 456852 3380 456858 3392
rect 458082 3380 458088 3392
rect 456852 3352 458088 3380
rect 456852 3340 456858 3352
rect 458082 3340 458088 3352
rect 458140 3340 458146 3392
rect 481634 3340 481640 3392
rect 481692 3380 481698 3392
rect 482462 3380 482468 3392
rect 481692 3352 482468 3380
rect 481692 3340 481698 3352
rect 482462 3340 482468 3352
rect 482520 3340 482526 3392
rect 489914 3340 489920 3392
rect 489972 3380 489978 3392
rect 490742 3380 490748 3392
rect 489972 3352 490748 3380
rect 489972 3340 489978 3352
rect 490742 3340 490748 3352
rect 490800 3340 490806 3392
rect 156414 3312 156420 3324
rect 146128 3284 156420 3312
rect 156414 3272 156420 3284
rect 156472 3272 156478 3324
rect 178678 3272 178684 3324
rect 178736 3312 178742 3324
rect 197906 3312 197912 3324
rect 178736 3284 197912 3312
rect 178736 3272 178742 3284
rect 197906 3272 197912 3284
rect 197964 3272 197970 3324
rect 202138 3272 202144 3324
rect 202196 3312 202202 3324
rect 245194 3312 245200 3324
rect 202196 3284 245200 3312
rect 202196 3272 202202 3284
rect 245194 3272 245200 3284
rect 245252 3272 245258 3324
rect 448514 3272 448520 3324
rect 448572 3312 448578 3324
rect 449802 3312 449808 3324
rect 448572 3284 449808 3312
rect 448572 3272 448578 3284
rect 449802 3272 449808 3284
rect 449860 3272 449866 3324
rect 142798 3204 142804 3256
rect 142856 3244 142862 3256
rect 148318 3244 148324 3256
rect 142856 3216 148324 3244
rect 142856 3204 142862 3216
rect 148318 3204 148324 3216
rect 148376 3204 148382 3256
rect 153838 3204 153844 3256
rect 153896 3244 153902 3256
rect 158898 3244 158904 3256
rect 153896 3216 158904 3244
rect 153896 3204 153902 3216
rect 158898 3204 158904 3216
rect 158956 3204 158962 3256
rect 180058 3204 180064 3256
rect 180116 3244 180122 3256
rect 219250 3244 219256 3256
rect 180116 3216 219256 3244
rect 180116 3204 180122 3216
rect 219250 3204 219256 3216
rect 219308 3204 219314 3256
rect 177666 3136 177672 3188
rect 177724 3176 177730 3188
rect 186130 3176 186136 3188
rect 177724 3148 186136 3176
rect 177724 3136 177730 3148
rect 186130 3136 186136 3148
rect 186188 3136 186194 3188
rect 132954 3068 132960 3120
rect 133012 3108 133018 3120
rect 140130 3108 140136 3120
rect 133012 3080 140136 3108
rect 133012 3068 133018 3080
rect 140130 3068 140136 3080
rect 140188 3068 140194 3120
rect 145558 2932 145564 2984
rect 145616 2972 145622 2984
rect 150618 2972 150624 2984
rect 145616 2944 150624 2972
rect 145616 2932 145622 2944
rect 150618 2932 150624 2944
rect 150676 2932 150682 2984
rect 365714 1232 365720 1284
rect 365772 1272 365778 1284
rect 367002 1272 367008 1284
rect 365772 1244 367008 1272
rect 365772 1232 365778 1244
rect 367002 1232 367008 1244
rect 367060 1232 367066 1284
rect 440234 552 440240 604
rect 440292 592 440298 604
rect 441522 592 441528 604
rect 440292 564 441528 592
rect 440292 552 440298 564
rect 441522 552 441528 564
rect 441580 552 441586 604
<< via1 >>
rect 201500 702992 201552 703044
rect 202788 702992 202840 703044
rect 331220 702992 331272 703044
rect 332508 702992 332560 703044
rect 207664 700612 207716 700664
rect 218980 700612 219032 700664
rect 206284 700544 206336 700596
rect 283840 700544 283892 700596
rect 203524 700476 203576 700528
rect 348792 700476 348844 700528
rect 154120 700408 154172 700460
rect 189080 700408 189132 700460
rect 200764 700408 200816 700460
rect 413652 700408 413704 700460
rect 72976 700340 73028 700392
rect 119344 700340 119396 700392
rect 137836 700340 137888 700392
rect 189356 700340 189408 700392
rect 199384 700340 199436 700392
rect 478512 700340 478564 700392
rect 24308 700272 24360 700324
rect 189172 700272 189224 700324
rect 198004 700272 198056 700324
rect 543464 700272 543516 700324
rect 105452 699660 105504 699712
rect 106924 699660 106976 699712
rect 266360 697552 266412 697604
rect 267648 697552 267700 697604
rect 2780 683612 2832 683664
rect 6184 683612 6236 683664
rect 196624 683136 196676 683188
rect 579620 683136 579672 683188
rect 3424 670760 3476 670812
rect 189264 670760 189316 670812
rect 120724 670692 120776 670744
rect 580172 670692 580224 670744
rect 191104 643084 191156 643136
rect 580172 643084 580224 643136
rect 2780 632068 2832 632120
rect 4804 632068 4856 632120
rect 193864 630640 193916 630692
rect 579988 630640 580040 630692
rect 3516 618264 3568 618316
rect 190460 618264 190512 618316
rect 118700 616836 118752 616888
rect 580172 616836 580224 616888
rect 192484 590656 192536 590708
rect 580172 590656 580224 590708
rect 3148 579776 3200 579828
rect 7564 579776 7616 579828
rect 193956 576852 194008 576904
rect 580172 576852 580224 576904
rect 3056 565836 3108 565888
rect 191840 565836 191892 565888
rect 120816 563048 120868 563100
rect 580172 563048 580224 563100
rect 3332 553392 3384 553444
rect 116584 553392 116636 553444
rect 192576 536800 192628 536852
rect 579896 536800 579948 536852
rect 2964 527144 3016 527196
rect 15844 527144 15896 527196
rect 194048 524424 194100 524476
rect 580172 524424 580224 524476
rect 120908 510620 120960 510672
rect 580172 510620 580224 510672
rect 3332 474716 3384 474768
rect 19984 474716 20036 474768
rect 121000 456764 121052 456816
rect 579620 456764 579672 456816
rect 2964 422288 3016 422340
rect 22744 422288 22796 422340
rect 192668 418140 192720 418192
rect 579712 418140 579764 418192
rect 3332 409844 3384 409896
rect 189448 409844 189500 409896
rect 118608 404336 118660 404388
rect 580172 404336 580224 404388
rect 192760 378156 192812 378208
rect 580172 378156 580224 378208
rect 3332 371220 3384 371272
rect 22836 371220 22888 371272
rect 366364 364352 366416 364404
rect 580172 364352 580224 364404
rect 3332 357416 3384 357468
rect 190552 357416 190604 357468
rect 118516 351908 118568 351960
rect 580172 351908 580224 351960
rect 3332 345040 3384 345092
rect 116676 345040 116728 345092
rect 2780 319064 2832 319116
rect 4896 319064 4948 319116
rect 362224 311856 362276 311908
rect 580172 311856 580224 311908
rect 2872 304988 2924 305040
rect 188344 304988 188396 305040
rect 280804 298120 280856 298172
rect 580172 298120 580224 298172
rect 3332 292544 3384 292596
rect 79324 292544 79376 292596
rect 118792 275272 118844 275324
rect 234620 275272 234672 275324
rect 192852 271872 192904 271924
rect 580172 271872 580224 271924
rect 3240 266364 3292 266416
rect 22928 266364 22980 266416
rect 531964 258068 532016 258120
rect 579620 258068 579672 258120
rect 2872 253920 2924 253972
rect 188436 253920 188488 253972
rect 360844 244264 360896 244316
rect 580172 244264 580224 244316
rect 3240 240116 3292 240168
rect 119436 240116 119488 240168
rect 118424 239368 118476 239420
rect 280804 239368 280856 239420
rect 532056 218016 532108 218068
rect 580172 218016 580224 218068
rect 3332 213936 3384 213988
rect 24124 213936 24176 213988
rect 280804 205640 280856 205692
rect 580172 205640 580224 205692
rect 118332 202104 118384 202156
rect 360844 202104 360896 202156
rect 3332 201492 3384 201544
rect 190736 201492 190788 201544
rect 196716 191836 196768 191888
rect 580172 191836 580224 191888
rect 358084 178032 358136 178084
rect 580172 178032 580224 178084
rect 122104 165588 122156 165640
rect 579620 165588 579672 165640
rect 3332 162868 3384 162920
rect 29644 162868 29696 162920
rect 196900 151784 196952 151836
rect 579988 151784 580040 151836
rect 118884 149676 118936 149728
rect 299480 149676 299532 149728
rect 3332 149064 3384 149116
rect 189724 149064 189776 149116
rect 3976 148316 4028 148368
rect 189632 148316 189684 148368
rect 3700 144168 3752 144220
rect 190920 144168 190972 144220
rect 88340 142876 88392 142928
rect 190828 142876 190880 142928
rect 118240 142808 118292 142860
rect 280804 142808 280856 142860
rect 118056 141448 118108 141500
rect 169760 141448 169812 141500
rect 119160 141380 119212 141432
rect 429200 141380 429252 141432
rect 119252 140156 119304 140208
rect 364340 140156 364392 140208
rect 119068 140088 119120 140140
rect 494060 140088 494112 140140
rect 118976 140020 119028 140072
rect 558920 140020 558972 140072
rect 118148 139408 118200 139460
rect 122104 139408 122156 139460
rect 188344 139340 188396 139392
rect 191932 139340 191984 139392
rect 188436 139272 188488 139324
rect 192024 139272 192076 139324
rect 3700 137980 3752 138032
rect 190644 137980 190696 138032
rect 2780 136688 2832 136740
rect 4988 136688 5040 136740
rect 23020 136620 23072 136672
rect 117320 136620 117372 136672
rect 24216 135260 24268 135312
rect 117320 135260 117372 135312
rect 190644 134444 190696 134496
rect 191012 134444 191064 134496
rect 21364 133900 21416 133952
rect 117320 133900 117372 133952
rect 29644 133832 29696 133884
rect 117412 133832 117464 133884
rect 24124 132404 24176 132456
rect 117320 132404 117372 132456
rect 22928 131044 22980 131096
rect 117320 131044 117372 131096
rect 4896 129684 4948 129736
rect 117320 129684 117372 129736
rect 22836 128256 22888 128308
rect 117320 128256 117372 128308
rect 22744 126896 22796 126948
rect 117320 126896 117372 126948
rect 19984 124108 20036 124160
rect 117320 124108 117372 124160
rect 15844 122748 15896 122800
rect 117320 122748 117372 122800
rect 7564 121388 7616 121440
rect 117320 121388 117372 121440
rect 4804 120028 4856 120080
rect 117320 120028 117372 120080
rect 6184 118600 6236 118652
rect 117320 118600 117372 118652
rect 189264 118600 189316 118652
rect 189448 118600 189500 118652
rect 40040 117240 40092 117292
rect 117320 117240 117372 117292
rect 189172 117240 189224 117292
rect 189448 117240 189500 117292
rect 106924 115880 106976 115932
rect 117320 115880 117372 115932
rect 189080 114452 189132 114504
rect 189448 114452 189500 114504
rect 193128 113092 193180 113144
rect 207664 113092 207716 113144
rect 189724 111800 189776 111852
rect 580080 111800 580132 111852
rect 3332 111732 3384 111784
rect 21364 111732 21416 111784
rect 193128 111732 193180 111784
rect 206284 111732 206336 111784
rect 193036 110372 193088 110424
rect 203524 110372 203576 110424
rect 193036 108944 193088 108996
rect 200764 108944 200816 108996
rect 193128 106156 193180 106208
rect 199384 106156 199436 106208
rect 193128 104660 193180 104712
rect 198004 104660 198056 104712
rect 193128 103164 193180 103216
rect 196624 103164 196676 103216
rect 192208 101736 192260 101788
rect 193864 101736 193916 101788
rect 192208 100376 192260 100428
rect 193956 100376 194008 100428
rect 192208 98812 192260 98864
rect 194048 98812 194100 98864
rect 193128 97928 193180 97980
rect 580448 97928 580500 97980
rect 193128 95140 193180 95192
rect 366364 95140 366416 95192
rect 193128 93780 193180 93832
rect 362224 93780 362276 93832
rect 193128 92420 193180 92472
rect 531964 92420 532016 92472
rect 193128 89632 193180 89684
rect 532056 89632 532108 89684
rect 193128 88272 193180 88324
rect 358084 88272 358136 88324
rect 193128 86912 193180 86964
rect 580724 86912 580776 86964
rect 193128 85484 193180 85536
rect 580908 85484 580960 85536
rect 192852 81404 192904 81456
rect 347044 81404 347096 81456
rect 118608 80928 118660 80980
rect 579988 80928 580040 80980
rect 4988 80792 5040 80844
rect 3700 80656 3752 80708
rect 179788 80656 179840 80708
rect 179512 80588 179564 80640
rect 127808 80384 127860 80436
rect 129372 80248 129424 80300
rect 129280 80112 129332 80164
rect 116584 79772 116636 79824
rect 130476 79976 130528 80028
rect 130706 79908 130758 79960
rect 130798 79908 130850 79960
rect 130660 79772 130712 79824
rect 130752 79772 130804 79824
rect 131350 79908 131402 79960
rect 131810 79908 131862 79960
rect 132086 79908 132138 79960
rect 132178 79908 132230 79960
rect 132270 79908 132322 79960
rect 132362 79908 132414 79960
rect 132638 79908 132690 79960
rect 133374 79908 133426 79960
rect 130568 79704 130620 79756
rect 131442 79840 131494 79892
rect 131764 79704 131816 79756
rect 132132 79704 132184 79756
rect 132224 79704 132276 79756
rect 131304 79636 131356 79688
rect 132316 79636 132368 79688
rect 132500 79636 132552 79688
rect 133006 79840 133058 79892
rect 132776 79636 132828 79688
rect 133236 79636 133288 79688
rect 133834 79908 133886 79960
rect 133926 79908 133978 79960
rect 135122 79908 135174 79960
rect 135214 79908 135266 79960
rect 135398 79908 135450 79960
rect 135582 79908 135634 79960
rect 136226 79908 136278 79960
rect 136502 79908 136554 79960
rect 133558 79840 133610 79892
rect 134478 79840 134530 79892
rect 134938 79840 134990 79892
rect 133972 79772 134024 79824
rect 133512 79636 133564 79688
rect 134570 79772 134622 79824
rect 134662 79772 134714 79824
rect 116676 79500 116728 79552
rect 127808 79500 127860 79552
rect 79324 79432 79376 79484
rect 131672 79432 131724 79484
rect 4068 79364 4120 79416
rect 3884 79296 3936 79348
rect 134064 79364 134116 79416
rect 134524 79500 134576 79552
rect 134708 79432 134760 79484
rect 134616 79364 134668 79416
rect 135076 79636 135128 79688
rect 135352 79636 135404 79688
rect 135168 79568 135220 79620
rect 135766 79840 135818 79892
rect 135858 79840 135910 79892
rect 135950 79840 136002 79892
rect 136042 79840 136094 79892
rect 135720 79704 135772 79756
rect 135812 79704 135864 79756
rect 135628 79568 135680 79620
rect 136318 79772 136370 79824
rect 136456 79772 136508 79824
rect 136088 79568 136140 79620
rect 135996 79500 136048 79552
rect 135536 79432 135588 79484
rect 136272 79432 136324 79484
rect 136870 79908 136922 79960
rect 137054 79908 137106 79960
rect 137238 79908 137290 79960
rect 137514 79908 137566 79960
rect 137974 79908 138026 79960
rect 138066 79908 138118 79960
rect 138158 79908 138210 79960
rect 138434 79908 138486 79960
rect 138526 79908 138578 79960
rect 137192 79636 137244 79688
rect 136640 79500 136692 79552
rect 137008 79500 137060 79552
rect 137422 79840 137474 79892
rect 138434 79772 138486 79824
rect 137928 79636 137980 79688
rect 138112 79636 138164 79688
rect 138020 79568 138072 79620
rect 137376 79500 137428 79552
rect 137652 79432 137704 79484
rect 138204 79432 138256 79484
rect 138480 79568 138532 79620
rect 138894 79908 138946 79960
rect 138986 79908 139038 79960
rect 139262 79908 139314 79960
rect 139354 79908 139406 79960
rect 138710 79840 138762 79892
rect 139538 79840 139590 79892
rect 139630 79772 139682 79824
rect 138940 79636 138992 79688
rect 139216 79636 139268 79688
rect 139308 79636 139360 79688
rect 139492 79636 139544 79688
rect 138664 79500 138716 79552
rect 139492 79500 139544 79552
rect 139998 79908 140050 79960
rect 140090 79908 140142 79960
rect 140182 79908 140234 79960
rect 141838 79908 141890 79960
rect 142390 79908 142442 79960
rect 142850 79908 142902 79960
rect 143218 79908 143270 79960
rect 144322 79908 144374 79960
rect 139952 79636 140004 79688
rect 136916 79364 136968 79416
rect 137468 79364 137520 79416
rect 138848 79364 138900 79416
rect 139124 79364 139176 79416
rect 139768 79364 139820 79416
rect 139952 79364 140004 79416
rect 140458 79840 140510 79892
rect 140734 79840 140786 79892
rect 140918 79840 140970 79892
rect 141010 79840 141062 79892
rect 141470 79840 141522 79892
rect 141654 79840 141706 79892
rect 140366 79772 140418 79824
rect 140228 79704 140280 79756
rect 140412 79636 140464 79688
rect 140780 79568 140832 79620
rect 141102 79772 141154 79824
rect 141286 79772 141338 79824
rect 141378 79704 141430 79756
rect 141056 79568 141108 79620
rect 140964 79500 141016 79552
rect 140596 79432 140648 79484
rect 141148 79364 141200 79416
rect 141792 79704 141844 79756
rect 141884 79704 141936 79756
rect 142252 79636 142304 79688
rect 142942 79840 142994 79892
rect 143862 79840 143914 79892
rect 144230 79840 144282 79892
rect 143080 79636 143132 79688
rect 143172 79636 143224 79688
rect 144000 79636 144052 79688
rect 144276 79636 144328 79688
rect 144690 79908 144742 79960
rect 144874 79908 144926 79960
rect 144644 79636 144696 79688
rect 145794 79908 145846 79960
rect 145978 79908 146030 79960
rect 145334 79840 145386 79892
rect 145518 79772 145570 79824
rect 145656 79636 145708 79688
rect 145748 79636 145800 79688
rect 145932 79636 145984 79688
rect 141608 79568 141660 79620
rect 144552 79568 144604 79620
rect 144828 79568 144880 79620
rect 145012 79568 145064 79620
rect 145104 79568 145156 79620
rect 145472 79568 145524 79620
rect 146162 79840 146214 79892
rect 146714 79908 146766 79960
rect 147358 79908 147410 79960
rect 148278 79908 148330 79960
rect 148370 79908 148422 79960
rect 148462 79908 148514 79960
rect 148554 79908 148606 79960
rect 148922 79908 148974 79960
rect 149198 79908 149250 79960
rect 150854 79908 150906 79960
rect 151038 79908 151090 79960
rect 146530 79840 146582 79892
rect 146806 79840 146858 79892
rect 146990 79840 147042 79892
rect 147312 79772 147364 79824
rect 147542 79772 147594 79824
rect 147726 79772 147778 79824
rect 148094 79772 148146 79824
rect 148232 79772 148284 79824
rect 146300 79636 146352 79688
rect 146576 79636 146628 79688
rect 146668 79636 146720 79688
rect 146392 79568 146444 79620
rect 146944 79568 146996 79620
rect 147864 79500 147916 79552
rect 147956 79500 148008 79552
rect 148416 79704 148468 79756
rect 148508 79704 148560 79756
rect 148738 79840 148790 79892
rect 148600 79636 148652 79688
rect 149382 79840 149434 79892
rect 149474 79840 149526 79892
rect 149566 79840 149618 79892
rect 149244 79704 149296 79756
rect 149336 79704 149388 79756
rect 148876 79636 148928 79688
rect 150302 79772 150354 79824
rect 150486 79772 150538 79824
rect 150670 79772 150722 79824
rect 149520 79636 149572 79688
rect 150164 79636 150216 79688
rect 148692 79568 148744 79620
rect 149428 79568 149480 79620
rect 151866 79908 151918 79960
rect 152418 79908 152470 79960
rect 152878 79908 152930 79960
rect 152970 79908 153022 79960
rect 151084 79772 151136 79824
rect 150992 79704 151044 79756
rect 150716 79636 150768 79688
rect 150624 79568 150676 79620
rect 151544 79568 151596 79620
rect 152326 79840 152378 79892
rect 152418 79772 152470 79824
rect 153016 79772 153068 79824
rect 152372 79636 152424 79688
rect 148784 79500 148836 79552
rect 153430 79908 153482 79960
rect 153614 79908 153666 79960
rect 153292 79500 153344 79552
rect 153890 79908 153942 79960
rect 153982 79908 154034 79960
rect 154074 79908 154126 79960
rect 153798 79840 153850 79892
rect 153844 79704 153896 79756
rect 153752 79636 153804 79688
rect 153568 79568 153620 79620
rect 153660 79500 153712 79552
rect 154350 79908 154402 79960
rect 154166 79772 154218 79824
rect 154258 79772 154310 79824
rect 154212 79636 154264 79688
rect 154810 79908 154862 79960
rect 155270 79908 155322 79960
rect 156098 79908 156150 79960
rect 156374 79908 156426 79960
rect 154718 79840 154770 79892
rect 155454 79772 155506 79824
rect 154764 79636 154816 79688
rect 155316 79636 155368 79688
rect 154580 79568 154632 79620
rect 154396 79500 154448 79552
rect 154488 79500 154540 79552
rect 154672 79500 154724 79552
rect 156466 79840 156518 79892
rect 156374 79772 156426 79824
rect 156052 79568 156104 79620
rect 156144 79568 156196 79620
rect 156834 79908 156886 79960
rect 156926 79908 156978 79960
rect 157662 79908 157714 79960
rect 156742 79840 156794 79892
rect 156788 79704 156840 79756
rect 156236 79500 156288 79552
rect 156696 79500 156748 79552
rect 157294 79840 157346 79892
rect 157156 79568 157208 79620
rect 180248 80520 180300 80572
rect 158030 79908 158082 79960
rect 157800 79568 157852 79620
rect 158214 79840 158266 79892
rect 158076 79568 158128 79620
rect 158490 79908 158542 79960
rect 158766 79908 158818 79960
rect 158858 79908 158910 79960
rect 158398 79840 158450 79892
rect 158352 79704 158404 79756
rect 159134 79840 159186 79892
rect 159502 79840 159554 79892
rect 159686 79908 159738 79960
rect 160790 79908 160842 79960
rect 161066 79908 161118 79960
rect 160146 79840 160198 79892
rect 160422 79840 160474 79892
rect 160698 79840 160750 79892
rect 158812 79704 158864 79756
rect 158536 79568 158588 79620
rect 158628 79568 158680 79620
rect 159548 79636 159600 79688
rect 159272 79568 159324 79620
rect 160284 79568 160336 79620
rect 160882 79840 160934 79892
rect 160744 79704 160796 79756
rect 160836 79704 160888 79756
rect 161342 79908 161394 79960
rect 161434 79908 161486 79960
rect 161480 79704 161532 79756
rect 162538 79908 162590 79960
rect 162630 79908 162682 79960
rect 161710 79840 161762 79892
rect 161894 79840 161946 79892
rect 162354 79840 162406 79892
rect 161572 79636 161624 79688
rect 158444 79500 158496 79552
rect 160376 79500 160428 79552
rect 160652 79500 160704 79552
rect 161020 79568 161072 79620
rect 161112 79568 161164 79620
rect 161296 79568 161348 79620
rect 161204 79500 161256 79552
rect 161480 79500 161532 79552
rect 162584 79772 162636 79824
rect 162814 79908 162866 79960
rect 162998 79908 163050 79960
rect 163090 79840 163142 79892
rect 163182 79840 163234 79892
rect 163366 79840 163418 79892
rect 163044 79636 163096 79688
rect 163228 79636 163280 79688
rect 162308 79568 162360 79620
rect 162492 79568 162544 79620
rect 162676 79568 162728 79620
rect 162860 79568 162912 79620
rect 163642 79772 163694 79824
rect 163918 79908 163970 79960
rect 163780 79636 163832 79688
rect 163688 79568 163740 79620
rect 164102 79840 164154 79892
rect 164056 79636 164108 79688
rect 164148 79568 164200 79620
rect 162124 79500 162176 79552
rect 164332 79500 164384 79552
rect 164654 79908 164706 79960
rect 165206 79908 165258 79960
rect 165666 79908 165718 79960
rect 165758 79908 165810 79960
rect 164562 79840 164614 79892
rect 164746 79840 164798 79892
rect 164608 79568 164660 79620
rect 165298 79840 165350 79892
rect 165390 79772 165442 79824
rect 165252 79704 165304 79756
rect 165850 79840 165902 79892
rect 166034 79840 166086 79892
rect 166310 79840 166362 79892
rect 166402 79840 166454 79892
rect 166218 79772 166270 79824
rect 165896 79704 165948 79756
rect 165988 79704 166040 79756
rect 165804 79636 165856 79688
rect 166172 79636 166224 79688
rect 165436 79568 165488 79620
rect 165528 79568 165580 79620
rect 165712 79568 165764 79620
rect 164792 79500 164844 79552
rect 164976 79500 165028 79552
rect 165344 79500 165396 79552
rect 166172 79500 166224 79552
rect 147680 79364 147732 79416
rect 153476 79432 153528 79484
rect 179696 80384 179748 80436
rect 179972 80180 180024 80232
rect 292580 80248 292632 80300
rect 316040 80180 316092 80232
rect 166862 79908 166914 79960
rect 166770 79840 166822 79892
rect 166816 79704 166868 79756
rect 166816 79568 166868 79620
rect 167414 79908 167466 79960
rect 167506 79908 167558 79960
rect 167138 79840 167190 79892
rect 167368 79772 167420 79824
rect 167460 79636 167512 79688
rect 167276 79568 167328 79620
rect 166632 79500 166684 79552
rect 167874 79840 167926 79892
rect 167966 79772 168018 79824
rect 168334 79908 168386 79960
rect 168150 79840 168202 79892
rect 168196 79704 168248 79756
rect 169162 79908 169214 79960
rect 169346 79908 169398 79960
rect 169438 79908 169490 79960
rect 170358 79908 170410 79960
rect 168426 79840 168478 79892
rect 168610 79840 168662 79892
rect 167920 79568 167972 79620
rect 168288 79636 168340 79688
rect 168104 79568 168156 79620
rect 168518 79772 168570 79824
rect 168702 79772 168754 79824
rect 168564 79568 168616 79620
rect 169254 79840 169306 79892
rect 169208 79704 169260 79756
rect 169300 79704 169352 79756
rect 169622 79840 169674 79892
rect 169898 79840 169950 79892
rect 169990 79840 170042 79892
rect 169484 79704 169536 79756
rect 168932 79636 168984 79688
rect 169116 79636 169168 79688
rect 168380 79500 168432 79552
rect 169392 79500 169444 79552
rect 169760 79568 169812 79620
rect 170082 79772 170134 79824
rect 170128 79636 170180 79688
rect 169944 79500 169996 79552
rect 170128 79500 170180 79552
rect 170634 79908 170686 79960
rect 170818 79908 170870 79960
rect 171002 79908 171054 79960
rect 170588 79772 170640 79824
rect 170496 79704 170548 79756
rect 170588 79568 170640 79620
rect 170496 79500 170548 79552
rect 170680 79500 170732 79552
rect 171048 79772 171100 79824
rect 170956 79636 171008 79688
rect 171370 79908 171422 79960
rect 172566 79908 172618 79960
rect 173026 79908 173078 79960
rect 173210 79908 173262 79960
rect 171830 79840 171882 79892
rect 172014 79772 172066 79824
rect 172198 79772 172250 79824
rect 172290 79772 172342 79824
rect 171784 79704 171836 79756
rect 171968 79568 172020 79620
rect 172842 79840 172894 79892
rect 172428 79568 172480 79620
rect 172152 79500 172204 79552
rect 172244 79500 172296 79552
rect 172888 79636 172940 79688
rect 173486 79840 173538 79892
rect 173854 79840 173906 79892
rect 174222 79840 174274 79892
rect 174314 79840 174366 79892
rect 173164 79636 173216 79688
rect 174498 79772 174550 79824
rect 173854 79636 173906 79688
rect 174176 79636 174228 79688
rect 174360 79636 174412 79688
rect 174452 79636 174504 79688
rect 179604 80112 179656 80164
rect 180156 80112 180208 80164
rect 180248 80112 180300 80164
rect 374000 80112 374052 80164
rect 179880 80044 179932 80096
rect 547972 80044 548024 80096
rect 179696 79976 179748 80028
rect 174774 79908 174826 79960
rect 175142 79908 175194 79960
rect 175418 79908 175470 79960
rect 175602 79908 175654 79960
rect 175970 79908 176022 79960
rect 174912 79636 174964 79688
rect 175004 79636 175056 79688
rect 175326 79840 175378 79892
rect 175878 79840 175930 79892
rect 175464 79704 175516 79756
rect 175556 79704 175608 79756
rect 176062 79840 176114 79892
rect 176246 79840 176298 79892
rect 176154 79772 176206 79824
rect 176062 79636 176114 79688
rect 175188 79568 175240 79620
rect 175372 79568 175424 79620
rect 175924 79568 175976 79620
rect 173164 79500 173216 79552
rect 176614 79908 176666 79960
rect 176706 79908 176758 79960
rect 177074 79908 177126 79960
rect 177166 79908 177218 79960
rect 177534 79908 177586 79960
rect 177626 79908 177678 79960
rect 176430 79840 176482 79892
rect 176752 79772 176804 79824
rect 176568 79704 176620 79756
rect 176660 79636 176712 79688
rect 177258 79840 177310 79892
rect 177580 79772 177632 79824
rect 177902 79908 177954 79960
rect 178086 79908 178138 79960
rect 178730 79908 178782 79960
rect 179190 79908 179242 79960
rect 179512 79908 179564 79960
rect 178178 79840 178230 79892
rect 178546 79840 178598 79892
rect 178086 79772 178138 79824
rect 177856 79704 177908 79756
rect 177304 79636 177356 79688
rect 177672 79636 177724 79688
rect 177764 79636 177816 79688
rect 177120 79568 177172 79620
rect 177212 79568 177264 79620
rect 177948 79568 178000 79620
rect 178040 79568 178092 79620
rect 178408 79636 178460 79688
rect 178500 79568 178552 79620
rect 178914 79840 178966 79892
rect 179696 79840 179748 79892
rect 179006 79772 179058 79824
rect 362960 79772 363012 79824
rect 179144 79704 179196 79756
rect 179788 79704 179840 79756
rect 179972 79636 180024 79688
rect 523132 79636 523184 79688
rect 179144 79568 179196 79620
rect 189724 79500 189776 79552
rect 134248 79228 134300 79280
rect 149612 79296 149664 79348
rect 164332 79364 164384 79416
rect 167736 79432 167788 79484
rect 165620 79364 165672 79416
rect 168288 79364 168340 79416
rect 171416 79364 171468 79416
rect 171600 79432 171652 79484
rect 171876 79432 171928 79484
rect 172060 79432 172112 79484
rect 178224 79432 178276 79484
rect 178868 79364 178920 79416
rect 138296 79160 138348 79212
rect 138756 79160 138808 79212
rect 139124 79160 139176 79212
rect 141332 79160 141384 79212
rect 153476 79228 153528 79280
rect 157800 79228 157852 79280
rect 162768 79228 162820 79280
rect 159180 79160 159232 79212
rect 161296 79160 161348 79212
rect 162032 79160 162084 79212
rect 162400 79160 162452 79212
rect 165620 79228 165672 79280
rect 167736 79228 167788 79280
rect 168564 79228 168616 79280
rect 171876 79228 171928 79280
rect 175280 79296 175332 79348
rect 176200 79296 176252 79348
rect 176292 79296 176344 79348
rect 178132 79296 178184 79348
rect 179788 79296 179840 79348
rect 527180 79296 527232 79348
rect 178684 79228 178736 79280
rect 180156 79228 180208 79280
rect 192760 79228 192812 79280
rect 166908 79160 166960 79212
rect 170956 79160 171008 79212
rect 171416 79160 171468 79212
rect 175648 79160 175700 79212
rect 176200 79160 176252 79212
rect 178316 79160 178368 79212
rect 180064 79160 180116 79212
rect 192944 79160 192996 79212
rect 130476 79024 130528 79076
rect 134248 79024 134300 79076
rect 135260 79024 135312 79076
rect 137100 79024 137152 79076
rect 139860 79024 139912 79076
rect 140136 79024 140188 79076
rect 144920 79024 144972 79076
rect 147680 79024 147732 79076
rect 3792 78956 3844 79008
rect 133880 78956 133932 79008
rect 138664 78956 138716 79008
rect 131672 78888 131724 78940
rect 144920 78888 144972 78940
rect 147220 78956 147272 79008
rect 150532 79092 150584 79144
rect 164332 79092 164384 79144
rect 168288 79092 168340 79144
rect 169392 79092 169444 79144
rect 156236 78956 156288 79008
rect 159916 78956 159968 79008
rect 162124 78956 162176 79008
rect 162216 78956 162268 79008
rect 162400 78956 162452 79008
rect 162768 78956 162820 79008
rect 168564 78956 168616 79008
rect 169668 79024 169720 79076
rect 172060 79024 172112 79076
rect 172612 79092 172664 79144
rect 176752 79092 176804 79144
rect 180708 79092 180760 79144
rect 201500 79092 201552 79144
rect 274640 79024 274692 79076
rect 171140 78956 171192 79008
rect 171508 78956 171560 79008
rect 173256 78956 173308 79008
rect 178592 78956 178644 79008
rect 3516 78820 3568 78872
rect 147220 78820 147272 78872
rect 157708 78820 157760 78872
rect 157984 78820 158036 78872
rect 158260 78820 158312 78872
rect 171048 78888 171100 78940
rect 172612 78888 172664 78940
rect 313280 78888 313332 78940
rect 133880 78752 133932 78804
rect 138664 78752 138716 78804
rect 150532 78752 150584 78804
rect 165620 78752 165672 78804
rect 169668 78752 169720 78804
rect 171876 78820 171928 78872
rect 178500 78820 178552 78872
rect 178408 78752 178460 78804
rect 178592 78752 178644 78804
rect 179236 78752 179288 78804
rect 126244 78684 126296 78736
rect 132684 78684 132736 78736
rect 157064 78684 157116 78736
rect 157984 78684 158036 78736
rect 168288 78684 168340 78736
rect 126336 78616 126388 78668
rect 133236 78616 133288 78668
rect 133328 78616 133380 78668
rect 133880 78616 133932 78668
rect 137100 78616 137152 78668
rect 138020 78616 138072 78668
rect 151912 78616 151964 78668
rect 169392 78616 169444 78668
rect 177856 78684 177908 78736
rect 174636 78616 174688 78668
rect 174820 78616 174872 78668
rect 174912 78616 174964 78668
rect 175188 78616 175240 78668
rect 176200 78616 176252 78668
rect 176568 78616 176620 78668
rect 127624 78548 127676 78600
rect 140320 78548 140372 78600
rect 149704 78548 149756 78600
rect 156696 78548 156748 78600
rect 168104 78548 168156 78600
rect 176476 78548 176528 78600
rect 177120 78548 177172 78600
rect 192484 78548 192536 78600
rect 143724 78480 143776 78532
rect 144184 78480 144236 78532
rect 153384 78480 153436 78532
rect 166816 78480 166868 78532
rect 170956 78480 171008 78532
rect 171508 78480 171560 78532
rect 177028 78480 177080 78532
rect 192576 78480 192628 78532
rect 129096 78412 129148 78464
rect 138848 78412 138900 78464
rect 162584 78412 162636 78464
rect 177672 78412 177724 78464
rect 177948 78412 178000 78464
rect 189356 78412 189408 78464
rect 130016 78344 130068 78396
rect 131120 78344 131172 78396
rect 134064 78344 134116 78396
rect 134616 78344 134668 78396
rect 170036 78344 170088 78396
rect 170404 78344 170456 78396
rect 171324 78344 171376 78396
rect 171600 78344 171652 78396
rect 175740 78344 175792 78396
rect 187608 78344 187660 78396
rect 96620 78208 96672 78260
rect 129648 78276 129700 78328
rect 145748 78276 145800 78328
rect 155776 78276 155828 78328
rect 177488 78276 177540 78328
rect 138112 78208 138164 78260
rect 143908 78208 143960 78260
rect 144092 78208 144144 78260
rect 155316 78208 155368 78260
rect 166908 78208 166960 78260
rect 167092 78208 167144 78260
rect 186136 78208 186188 78260
rect 186412 78208 186464 78260
rect 268384 78208 268436 78260
rect 78680 78140 78732 78192
rect 136732 78140 136784 78192
rect 161756 78140 161808 78192
rect 162032 78140 162084 78192
rect 164332 78140 164384 78192
rect 164608 78140 164660 78192
rect 164884 78140 164936 78192
rect 180156 78140 180208 78192
rect 187608 78140 187660 78192
rect 337384 78140 337436 78192
rect 10324 78072 10376 78124
rect 130936 78072 130988 78124
rect 131120 78072 131172 78124
rect 133972 78072 134024 78124
rect 43444 78004 43496 78056
rect 132132 78004 132184 78056
rect 137008 78004 137060 78056
rect 137376 78004 137428 78056
rect 2780 77936 2832 77988
rect 130844 77936 130896 77988
rect 130936 77936 130988 77988
rect 138572 77936 138624 77988
rect 131212 77732 131264 77784
rect 131580 77732 131632 77784
rect 139400 77732 139452 77784
rect 140596 77732 140648 77784
rect 144276 78072 144328 78124
rect 151360 78072 151412 78124
rect 155316 78072 155368 78124
rect 158812 78072 158864 78124
rect 166908 78072 166960 78124
rect 169024 78072 169076 78124
rect 169668 78072 169720 78124
rect 170220 78072 170272 78124
rect 170680 78072 170732 78124
rect 175924 78072 175976 78124
rect 349804 78072 349856 78124
rect 161204 78004 161256 78056
rect 164884 78004 164936 78056
rect 167552 78004 167604 78056
rect 431224 78004 431276 78056
rect 146484 77936 146536 77988
rect 151360 77936 151412 77988
rect 154948 77936 155000 77988
rect 161664 77868 161716 77920
rect 162400 77868 162452 77920
rect 164608 77936 164660 77988
rect 164976 77936 165028 77988
rect 168748 77936 168800 77988
rect 489920 77936 489972 77988
rect 172612 77868 172664 77920
rect 151636 77800 151688 77852
rect 162124 77800 162176 77852
rect 165804 77800 165856 77852
rect 166448 77800 166500 77852
rect 167368 77800 167420 77852
rect 167552 77800 167604 77852
rect 169944 77800 169996 77852
rect 170128 77800 170180 77852
rect 170588 77800 170640 77852
rect 170864 77800 170916 77852
rect 171048 77800 171100 77852
rect 171692 77800 171744 77852
rect 144368 77732 144420 77784
rect 150808 77732 150860 77784
rect 162400 77732 162452 77784
rect 164240 77732 164292 77784
rect 130568 77664 130620 77716
rect 138388 77664 138440 77716
rect 147864 77664 147916 77716
rect 129188 77596 129240 77648
rect 139676 77596 139728 77648
rect 145288 77596 145340 77648
rect 134524 77528 134576 77580
rect 136364 77528 136416 77580
rect 159824 77596 159876 77648
rect 165804 77664 165856 77716
rect 165988 77664 166040 77716
rect 169668 77732 169720 77784
rect 177396 77868 177448 77920
rect 176844 77800 176896 77852
rect 580356 77800 580408 77852
rect 177304 77732 177356 77784
rect 191104 77732 191156 77784
rect 177212 77664 177264 77716
rect 161112 77528 161164 77580
rect 168288 77596 168340 77648
rect 169760 77596 169812 77648
rect 177304 77596 177356 77648
rect 167736 77528 167788 77580
rect 168012 77528 168064 77580
rect 176292 77528 176344 77580
rect 158444 77460 158496 77512
rect 165436 77460 165488 77512
rect 166356 77460 166408 77512
rect 181444 77460 181496 77512
rect 130476 77392 130528 77444
rect 137836 77392 137888 77444
rect 155224 77392 155276 77444
rect 155776 77392 155828 77444
rect 158720 77392 158772 77444
rect 159640 77392 159692 77444
rect 160284 77392 160336 77444
rect 168012 77392 168064 77444
rect 177672 77392 177724 77444
rect 177856 77392 177908 77444
rect 178132 77392 178184 77444
rect 179420 77392 179472 77444
rect 130200 77324 130252 77376
rect 137652 77324 137704 77376
rect 164240 77324 164292 77376
rect 165160 77324 165212 77376
rect 165620 77324 165672 77376
rect 175832 77324 175884 77376
rect 131764 77256 131816 77308
rect 135812 77256 135864 77308
rect 145380 77256 145432 77308
rect 147220 77256 147272 77308
rect 151912 77256 151964 77308
rect 152924 77256 152976 77308
rect 153384 77256 153436 77308
rect 154120 77256 154172 77308
rect 154580 77256 154632 77308
rect 154948 77256 155000 77308
rect 158904 77256 158956 77308
rect 159088 77256 159140 77308
rect 173072 77256 173124 77308
rect 176384 77256 176436 77308
rect 176752 77256 176804 77308
rect 177856 77256 177908 77308
rect 150440 77188 150492 77240
rect 151084 77188 151136 77240
rect 153200 77188 153252 77240
rect 153752 77188 153804 77240
rect 154764 77188 154816 77240
rect 158628 77188 158680 77240
rect 160376 77188 160428 77240
rect 160836 77188 160888 77240
rect 161112 77188 161164 77240
rect 186320 77188 186372 77240
rect 145932 77120 145984 77172
rect 171876 77120 171928 77172
rect 140596 77052 140648 77104
rect 141056 77052 141108 77104
rect 132592 76984 132644 77036
rect 132960 76984 133012 77036
rect 156696 76984 156748 77036
rect 240140 77052 240192 77104
rect 157524 76984 157576 77036
rect 158076 76984 158128 77036
rect 171140 76984 171192 77036
rect 260840 76984 260892 77036
rect 151452 76916 151504 76968
rect 267740 76916 267792 76968
rect 126980 76848 127032 76900
rect 140504 76848 140556 76900
rect 142712 76848 142764 76900
rect 143080 76848 143132 76900
rect 150532 76848 150584 76900
rect 150716 76848 150768 76900
rect 157432 76848 157484 76900
rect 158260 76848 158312 76900
rect 165620 76848 165672 76900
rect 166172 76848 166224 76900
rect 171048 76848 171100 76900
rect 327080 76848 327132 76900
rect 91100 76780 91152 76832
rect 137744 76780 137796 76832
rect 142068 76780 142120 76832
rect 142528 76780 142580 76832
rect 156880 76780 156932 76832
rect 328460 76780 328512 76832
rect 104900 76712 104952 76764
rect 138296 76712 138348 76764
rect 142436 76712 142488 76764
rect 143080 76712 143132 76764
rect 147864 76712 147916 76764
rect 148416 76712 148468 76764
rect 157432 76712 157484 76764
rect 158168 76712 158220 76764
rect 160100 76712 160152 76764
rect 160376 76712 160428 76764
rect 160744 76712 160796 76764
rect 161296 76712 161348 76764
rect 84200 76644 84252 76696
rect 135260 76644 135312 76696
rect 159180 76644 159232 76696
rect 159732 76644 159784 76696
rect 41420 76576 41472 76628
rect 133512 76576 133564 76628
rect 154764 76576 154816 76628
rect 155592 76576 155644 76628
rect 155960 76576 156012 76628
rect 156420 76576 156472 76628
rect 158812 76576 158864 76628
rect 159364 76576 159416 76628
rect 34520 76508 34572 76560
rect 133052 76508 133104 76560
rect 158904 76508 158956 76560
rect 159456 76508 159508 76560
rect 165344 76644 165396 76696
rect 165896 76644 165948 76696
rect 172060 76712 172112 76764
rect 368480 76712 368532 76764
rect 367100 76644 367152 76696
rect 160744 76576 160796 76628
rect 161020 76576 161072 76628
rect 161572 76576 161624 76628
rect 161940 76576 161992 76628
rect 162124 76576 162176 76628
rect 171140 76576 171192 76628
rect 160468 76508 160520 76560
rect 160928 76508 160980 76560
rect 166172 76508 166224 76560
rect 166540 76508 166592 76560
rect 168380 76508 168432 76560
rect 485780 76576 485832 76628
rect 147956 76440 148008 76492
rect 148140 76440 148192 76492
rect 149336 76440 149388 76492
rect 149796 76440 149848 76492
rect 158996 76440 159048 76492
rect 159548 76440 159600 76492
rect 160376 76440 160428 76492
rect 160652 76440 160704 76492
rect 161204 76440 161256 76492
rect 161940 76440 161992 76492
rect 162308 76440 162360 76492
rect 171876 76440 171928 76492
rect 178684 76440 178736 76492
rect 152280 76372 152332 76424
rect 152556 76372 152608 76424
rect 162216 76372 162268 76424
rect 172060 76372 172112 76424
rect 173164 76372 173216 76424
rect 542360 76508 542412 76560
rect 147956 76304 148008 76356
rect 148508 76304 148560 76356
rect 154580 76304 154632 76356
rect 155500 76304 155552 76356
rect 168380 76304 168432 76356
rect 168840 76304 168892 76356
rect 149152 76236 149204 76288
rect 149704 76236 149756 76288
rect 144460 76168 144512 76220
rect 145748 76168 145800 76220
rect 163320 76168 163372 76220
rect 163504 76168 163556 76220
rect 139768 76100 139820 76152
rect 139952 76100 140004 76152
rect 149152 76100 149204 76152
rect 149428 76100 149480 76152
rect 168656 76100 168708 76152
rect 169116 76100 169168 76152
rect 139952 75964 140004 76016
rect 140228 75964 140280 76016
rect 143632 75964 143684 76016
rect 144460 75964 144512 76016
rect 142528 75896 142580 75948
rect 142804 75896 142856 75948
rect 150716 75896 150768 75948
rect 151084 75896 151136 75948
rect 140228 75828 140280 75880
rect 141240 75828 141292 75880
rect 150808 75828 150860 75880
rect 151176 75828 151228 75880
rect 152188 75828 152240 75880
rect 152648 75828 152700 75880
rect 152004 75760 152056 75812
rect 152280 75760 152332 75812
rect 169576 75760 169628 75812
rect 175096 75760 175148 75812
rect 131028 75692 131080 75744
rect 137468 75692 137520 75744
rect 141240 75692 141292 75744
rect 141608 75692 141660 75744
rect 170680 75692 170732 75744
rect 175004 75692 175056 75744
rect 130108 75624 130160 75676
rect 140780 75624 140832 75676
rect 148324 75624 148376 75676
rect 176752 75624 176804 75676
rect 128360 75556 128412 75608
rect 140688 75556 140740 75608
rect 145656 75556 145708 75608
rect 191840 75556 191892 75608
rect 127072 75488 127124 75540
rect 140412 75488 140464 75540
rect 147496 75488 147548 75540
rect 201500 75488 201552 75540
rect 81440 75420 81492 75472
rect 131028 75420 131080 75472
rect 69020 75352 69072 75404
rect 135996 75420 136048 75472
rect 153200 75420 153252 75472
rect 154028 75420 154080 75472
rect 170496 75420 170548 75472
rect 51080 75284 51132 75336
rect 134616 75352 134668 75404
rect 139676 75352 139728 75404
rect 140044 75352 140096 75404
rect 142344 75352 142396 75404
rect 142620 75352 142672 75404
rect 164424 75352 164476 75404
rect 164884 75352 164936 75404
rect 171508 75352 171560 75404
rect 131396 75284 131448 75336
rect 132224 75284 132276 75336
rect 132684 75284 132736 75336
rect 133788 75284 133840 75336
rect 138572 75284 138624 75336
rect 139308 75284 139360 75336
rect 162952 75284 163004 75336
rect 164148 75284 164200 75336
rect 167184 75284 167236 75336
rect 167920 75284 167972 75336
rect 168748 75284 168800 75336
rect 169484 75284 169536 75336
rect 46940 75216 46992 75268
rect 131120 75216 131172 75268
rect 131580 75216 131632 75268
rect 132408 75216 132460 75268
rect 133052 75216 133104 75268
rect 133604 75216 133656 75268
rect 133880 75216 133932 75268
rect 134156 75216 134208 75268
rect 134248 75216 134300 75268
rect 134800 75216 134852 75268
rect 135996 75216 136048 75268
rect 136456 75216 136508 75268
rect 138296 75216 138348 75268
rect 139216 75216 139268 75268
rect 140044 75216 140096 75268
rect 140872 75216 140924 75268
rect 141332 75216 141384 75268
rect 141792 75216 141844 75268
rect 141884 75216 141936 75268
rect 142344 75216 142396 75268
rect 145288 75216 145340 75268
rect 146024 75216 146076 75268
rect 146760 75216 146812 75268
rect 146944 75216 146996 75268
rect 164424 75216 164476 75268
rect 165068 75216 165120 75268
rect 168840 75216 168892 75268
rect 169208 75216 169260 75268
rect 170312 75216 170364 75268
rect 170772 75216 170824 75268
rect 171508 75216 171560 75268
rect 171968 75216 172020 75268
rect 172612 75216 172664 75268
rect 173072 75216 173124 75268
rect 174360 75216 174412 75268
rect 174728 75216 174780 75268
rect 175096 75420 175148 75472
rect 499580 75420 499632 75472
rect 175004 75352 175056 75404
rect 506480 75352 506532 75404
rect 514760 75284 514812 75336
rect 521660 75216 521712 75268
rect 1400 75148 1452 75200
rect 130660 75148 130712 75200
rect 131488 75148 131540 75200
rect 132316 75148 132368 75200
rect 132960 75148 133012 75200
rect 133328 75148 133380 75200
rect 134340 75148 134392 75200
rect 134984 75148 135036 75200
rect 135536 75148 135588 75200
rect 136548 75148 136600 75200
rect 138388 75148 138440 75200
rect 139032 75148 139084 75200
rect 140136 75148 140188 75200
rect 140964 75148 141016 75200
rect 141056 75148 141108 75200
rect 141976 75148 142028 75200
rect 146484 75148 146536 75200
rect 147036 75148 147088 75200
rect 163044 75148 163096 75200
rect 163872 75148 163924 75200
rect 167092 75148 167144 75200
rect 167828 75148 167880 75200
rect 171140 75148 171192 75200
rect 172244 75148 172296 75200
rect 173440 75148 173492 75200
rect 549260 75148 549312 75200
rect 138020 75080 138072 75132
rect 139124 75080 139176 75132
rect 145748 75080 145800 75132
rect 146024 75080 146076 75132
rect 146760 75080 146812 75132
rect 147128 75080 147180 75132
rect 149428 75080 149480 75132
rect 149980 75080 150032 75132
rect 152004 75080 152056 75132
rect 152740 75080 152792 75132
rect 163320 75080 163372 75132
rect 163688 75080 163740 75132
rect 167368 75080 167420 75132
rect 167644 75080 167696 75132
rect 172612 75080 172664 75132
rect 173348 75080 173400 75132
rect 174360 75080 174412 75132
rect 175188 75080 175240 75132
rect 149336 75012 149388 75064
rect 150164 75012 150216 75064
rect 157892 75012 157944 75064
rect 170680 75012 170732 75064
rect 120724 74196 120776 74248
rect 135168 74196 135220 74248
rect 168104 74196 168156 74248
rect 185584 74196 185636 74248
rect 114560 74128 114612 74180
rect 139492 74128 139544 74180
rect 150256 74128 150308 74180
rect 202144 74128 202196 74180
rect 82820 74060 82872 74112
rect 136916 74060 136968 74112
rect 148600 74060 148652 74112
rect 230480 74060 230532 74112
rect 64880 73992 64932 74044
rect 136180 73992 136232 74044
rect 150992 73992 151044 74044
rect 259460 73992 259512 74044
rect 29000 73924 29052 73976
rect 132592 73924 132644 73976
rect 155316 73924 155368 73976
rect 266360 73924 266412 73976
rect 16580 73856 16632 73908
rect 131856 73856 131908 73908
rect 151544 73856 151596 73908
rect 273260 73856 273312 73908
rect 2872 73788 2924 73840
rect 130752 73788 130804 73840
rect 158260 73788 158312 73840
rect 343640 73788 343692 73840
rect 158536 73720 158588 73772
rect 159824 73720 159876 73772
rect 133880 73244 133932 73296
rect 140596 73244 140648 73296
rect 176200 73244 176252 73296
rect 177948 73244 178000 73296
rect 136916 73176 136968 73228
rect 141424 73176 141476 73228
rect 176016 73108 176068 73160
rect 580172 73108 580224 73160
rect 175832 73040 175884 73092
rect 176200 73040 176252 73092
rect 175280 72836 175332 72888
rect 176108 72836 176160 72888
rect 153936 72768 153988 72820
rect 293960 72768 294012 72820
rect 154396 72700 154448 72752
rect 300860 72700 300912 72752
rect 155776 72632 155828 72684
rect 316132 72632 316184 72684
rect 107660 72564 107712 72616
rect 138940 72564 138992 72616
rect 155684 72564 155736 72616
rect 322940 72564 322992 72616
rect 57980 72496 58032 72548
rect 135076 72496 135128 72548
rect 165436 72496 165488 72548
rect 347780 72496 347832 72548
rect 20 72428 72 72480
rect 130292 72428 130344 72480
rect 159824 72428 159876 72480
rect 354680 72428 354732 72480
rect 130384 72156 130436 72208
rect 136272 72156 136324 72208
rect 135628 71748 135680 71800
rect 139400 71748 139452 71800
rect 3424 71680 3476 71732
rect 24216 71680 24268 71732
rect 158628 71136 158680 71188
rect 309140 71136 309192 71188
rect 159640 71068 159692 71120
rect 360200 71068 360252 71120
rect 53840 71000 53892 71052
rect 134892 71000 134944 71052
rect 144368 71000 144420 71052
rect 175280 71000 175332 71052
rect 176476 71000 176528 71052
rect 487160 71000 487212 71052
rect 144184 69912 144236 69964
rect 178040 69912 178092 69964
rect 163780 69844 163832 69896
rect 415400 69844 415452 69896
rect 166356 69776 166408 69828
rect 451280 69776 451332 69828
rect 143080 69708 143132 69760
rect 151084 69708 151136 69760
rect 169024 69708 169076 69760
rect 498200 69708 498252 69760
rect 5540 69640 5592 69692
rect 130016 69640 130068 69692
rect 174728 69640 174780 69692
rect 561680 69640 561732 69692
rect 142804 68960 142856 69012
rect 145564 68960 145616 69012
rect 145840 68484 145892 68536
rect 195980 68484 196032 68536
rect 164884 68416 164936 68468
rect 433340 68416 433392 68468
rect 166264 68348 166316 68400
rect 456800 68348 456852 68400
rect 170588 68280 170640 68332
rect 514852 68280 514904 68332
rect 145380 67124 145432 67176
rect 193220 67124 193272 67176
rect 159272 67056 159324 67108
rect 365720 67056 365772 67108
rect 167552 66988 167604 67040
rect 473360 66988 473412 67040
rect 170312 66920 170364 66972
rect 512000 66920 512052 66972
rect 171784 66852 171836 66904
rect 529940 66852 529992 66904
rect 153844 65900 153896 65952
rect 295340 65900 295392 65952
rect 155224 65832 155276 65884
rect 307760 65832 307812 65884
rect 3516 65764 3568 65816
rect 190644 65764 190696 65816
rect 164792 65696 164844 65748
rect 437480 65696 437532 65748
rect 170220 65628 170272 65680
rect 510620 65628 510672 65680
rect 174544 65560 174596 65612
rect 564440 65560 564492 65612
rect 174636 65492 174688 65544
rect 568580 65492 568632 65544
rect 165252 64336 165304 64388
rect 382280 64336 382332 64388
rect 163504 64268 163556 64320
rect 419540 64268 419592 64320
rect 163596 64200 163648 64252
rect 423680 64200 423732 64252
rect 173808 64132 173860 64184
rect 552020 64132 552072 64184
rect 144092 63248 144144 63300
rect 145656 63248 145708 63300
rect 166632 62840 166684 62892
rect 361580 62840 361632 62892
rect 168932 62772 168984 62824
rect 488540 62772 488592 62824
rect 148416 61548 148468 61600
rect 223580 61548 223632 61600
rect 152556 61480 152608 61532
rect 277400 61480 277452 61532
rect 160836 61412 160888 61464
rect 380900 61412 380952 61464
rect 171692 61344 171744 61396
rect 525800 61344 525852 61396
rect 192668 60664 192720 60716
rect 580172 60664 580224 60716
rect 170128 60052 170180 60104
rect 506572 60052 506624 60104
rect 176384 59984 176436 60036
rect 539600 59984 539652 60036
rect 156604 58624 156656 58676
rect 333980 58624 334032 58676
rect 42800 57196 42852 57248
rect 129372 57196 129424 57248
rect 157800 55836 157852 55888
rect 346400 55836 346452 55888
rect 142712 51688 142764 51740
rect 153844 51688 153896 51740
rect 160744 51688 160796 51740
rect 390560 51688 390612 51740
rect 124220 51076 124272 51128
rect 127624 51076 127676 51128
rect 148324 48968 148376 49020
rect 226340 48968 226392 49020
rect 118516 46860 118568 46912
rect 580172 46860 580224 46912
rect 3424 45500 3476 45552
rect 178224 45500 178276 45552
rect 141332 44888 141384 44940
rect 142896 44888 142948 44940
rect 38660 44820 38712 44872
rect 133052 44820 133104 44872
rect 177212 44820 177264 44872
rect 432052 44820 432104 44872
rect 142620 44140 142672 44192
rect 144276 44140 144328 44192
rect 19340 39312 19392 39364
rect 129280 39312 129332 39364
rect 146944 35640 146996 35692
rect 205640 35640 205692 35692
rect 146852 35572 146904 35624
rect 209872 35572 209924 35624
rect 150900 35504 150952 35556
rect 255320 35504 255372 35556
rect 155132 35436 155184 35488
rect 311900 35436 311952 35488
rect 167920 35368 167972 35420
rect 375380 35368 375432 35420
rect 176200 35300 176252 35352
rect 397460 35300 397512 35352
rect 176292 35232 176344 35284
rect 404360 35232 404412 35284
rect 163412 35164 163464 35216
rect 422300 35164 422352 35216
rect 145196 34280 145248 34332
rect 187700 34280 187752 34332
rect 145104 34212 145156 34264
rect 194600 34212 194652 34264
rect 145288 34144 145340 34196
rect 198740 34144 198792 34196
rect 148232 34076 148284 34128
rect 226432 34076 226484 34128
rect 149796 34008 149848 34060
rect 241520 34008 241572 34060
rect 152464 33940 152516 33992
rect 280160 33940 280212 33992
rect 153752 33872 153804 33924
rect 291200 33872 291252 33924
rect 157708 33804 157760 33856
rect 350540 33804 350592 33856
rect 164700 33736 164752 33788
rect 441620 33736 441672 33788
rect 3516 33056 3568 33108
rect 23020 33056 23072 33108
rect 177948 33056 178000 33108
rect 580172 33056 580224 33108
rect 146760 32852 146812 32904
rect 212540 32852 212592 32904
rect 148140 32784 148192 32836
rect 219440 32784 219492 32836
rect 149704 32716 149756 32768
rect 237380 32716 237432 32768
rect 3424 32648 3476 32700
rect 178132 32648 178184 32700
rect 162032 32580 162084 32632
rect 400220 32580 400272 32632
rect 163320 32512 163372 32564
rect 423772 32512 423824 32564
rect 164516 32444 164568 32496
rect 434720 32444 434772 32496
rect 164608 32376 164660 32428
rect 438860 32376 438912 32428
rect 145012 31356 145064 31408
rect 185032 31356 185084 31408
rect 153660 31288 153712 31340
rect 292672 31288 292724 31340
rect 153568 31220 153620 31272
rect 299480 31220 299532 31272
rect 158352 31152 158404 31204
rect 339500 31152 339552 31204
rect 159180 31084 159232 31136
rect 374092 31084 374144 31136
rect 168840 31016 168892 31068
rect 496820 31016 496872 31068
rect 149520 29928 149572 29980
rect 242900 29928 242952 29980
rect 149612 29860 149664 29912
rect 247040 29860 247092 29912
rect 150808 29792 150860 29844
rect 264980 29792 265032 29844
rect 155040 29724 155092 29776
rect 317420 29724 317472 29776
rect 163228 29656 163280 29708
rect 416780 29656 416832 29708
rect 174452 29588 174504 29640
rect 564532 29588 564584 29640
rect 146668 28704 146720 28756
rect 208400 28704 208452 28756
rect 148048 28636 148100 28688
rect 222200 28636 222252 28688
rect 147956 28568 148008 28620
rect 229100 28568 229152 28620
rect 152372 28500 152424 28552
rect 278780 28500 278832 28552
rect 154948 28432 155000 28484
rect 310520 28432 310572 28484
rect 159088 28364 159140 28416
rect 364340 28364 364392 28416
rect 158996 28296 159048 28348
rect 372620 28296 372672 28348
rect 173072 28228 173124 28280
rect 539692 28228 539744 28280
rect 147220 27276 147272 27328
rect 190460 27276 190512 27328
rect 146116 27208 146168 27260
rect 193312 27208 193364 27260
rect 146576 27140 146628 27192
rect 204260 27140 204312 27192
rect 152280 27072 152332 27124
rect 276020 27072 276072 27124
rect 168012 27004 168064 27056
rect 379520 27004 379572 27056
rect 158904 26936 158956 26988
rect 371240 26936 371292 26988
rect 175372 26868 175424 26920
rect 574100 26868 574152 26920
rect 146484 25916 146536 25968
rect 211160 25916 211212 25968
rect 152188 25848 152240 25900
rect 282920 25848 282972 25900
rect 154856 25780 154908 25832
rect 314660 25780 314712 25832
rect 172888 25712 172940 25764
rect 349896 25712 349948 25764
rect 177764 25644 177816 25696
rect 411260 25644 411312 25696
rect 167460 25576 167512 25628
rect 473452 25576 473504 25628
rect 172980 25508 173032 25560
rect 546500 25508 546552 25560
rect 153476 24352 153528 24404
rect 296720 24352 296772 24404
rect 154764 24284 154816 24336
rect 321560 24284 321612 24336
rect 177580 24216 177632 24268
rect 418160 24216 418212 24268
rect 172796 24148 172848 24200
rect 540980 24148 541032 24200
rect 174360 24080 174412 24132
rect 567200 24080 567252 24132
rect 3240 22992 3292 23044
rect 189540 22992 189592 23044
rect 170036 22924 170088 22976
rect 513380 22924 513432 22976
rect 171600 22856 171652 22908
rect 528560 22856 528612 22908
rect 88340 22788 88392 22840
rect 137192 22788 137244 22840
rect 171508 22788 171560 22840
rect 531320 22788 531372 22840
rect 118332 22720 118384 22772
rect 580264 22720 580316 22772
rect 163136 21632 163188 21684
rect 415492 21632 415544 21684
rect 167368 21564 167420 21616
rect 476120 21564 476172 21616
rect 168656 21496 168708 21548
rect 495440 21496 495492 21548
rect 168748 21428 168800 21480
rect 498292 21428 498344 21480
rect 174268 21360 174320 21412
rect 563060 21360 563112 21412
rect 347044 20612 347096 20664
rect 579988 20612 580040 20664
rect 152096 20272 152148 20324
rect 276112 20272 276164 20324
rect 152004 20204 152056 20256
rect 284300 20204 284352 20256
rect 268384 20136 268436 20188
rect 467840 20136 467892 20188
rect 167276 20068 167328 20120
rect 228364 20068 228416 20120
rect 260104 20068 260156 20120
rect 460940 20068 460992 20120
rect 166172 20000 166224 20052
rect 462320 20000 462372 20052
rect 169944 19932 169996 19984
rect 509240 19932 509292 19984
rect 161940 18980 161992 19032
rect 407120 18980 407172 19032
rect 163044 18912 163096 18964
rect 426440 18912 426492 18964
rect 117320 18844 117372 18896
rect 129188 18844 129240 18896
rect 164424 18844 164476 18896
rect 440240 18844 440292 18896
rect 120080 18776 120132 18828
rect 139676 18776 139728 18828
rect 172704 18776 172756 18828
rect 553400 18776 553452 18828
rect 111800 18708 111852 18760
rect 138572 18708 138624 18760
rect 173992 18708 174044 18760
rect 556252 18708 556304 18760
rect 35900 18640 35952 18692
rect 126336 18640 126388 18692
rect 174084 18640 174136 18692
rect 558920 18640 558972 18692
rect 15200 18572 15252 18624
rect 131672 18572 131724 18624
rect 174176 18572 174228 18624
rect 560300 18572 560352 18624
rect 154672 17416 154724 17468
rect 318800 17416 318852 17468
rect 161848 17348 161900 17400
rect 405740 17348 405792 17400
rect 168564 17280 168616 17332
rect 492680 17280 492732 17332
rect 171416 17212 171468 17264
rect 531412 17212 531464 17264
rect 160560 16124 160612 16176
rect 384304 16124 384356 16176
rect 160652 16056 160704 16108
rect 387800 16056 387852 16108
rect 167092 15988 167144 16040
rect 478144 15988 478196 16040
rect 167184 15920 167236 15972
rect 478880 15920 478932 15972
rect 142528 15852 142580 15904
rect 156144 15852 156196 15904
rect 171324 15852 171376 15904
rect 527824 15852 527876 15904
rect 162400 15036 162452 15088
rect 256700 15036 256752 15088
rect 150716 14968 150768 15020
rect 262496 14968 262548 15020
rect 158812 14900 158864 14952
rect 370136 14900 370188 14952
rect 160468 14832 160520 14884
rect 390652 14832 390704 14884
rect 161756 14764 161808 14816
rect 398840 14764 398892 14816
rect 162860 14696 162912 14748
rect 420920 14696 420972 14748
rect 162952 14628 163004 14680
rect 428464 14628 428516 14680
rect 129556 14560 129608 14612
rect 402520 14560 402572 14612
rect 181444 14492 181496 14544
rect 454040 14492 454092 14544
rect 172612 14424 172664 14476
rect 465724 14424 465776 14476
rect 149428 13472 149480 13524
rect 248420 13472 248472 13524
rect 157616 13404 157668 13456
rect 345296 13404 345348 13456
rect 157524 13336 157576 13388
rect 352840 13336 352892 13388
rect 161572 13268 161624 13320
rect 403624 13268 403676 13320
rect 161664 13200 161716 13252
rect 407212 13200 407264 13252
rect 180248 13132 180300 13184
rect 447416 13132 447468 13184
rect 168472 13064 168524 13116
rect 490012 13064 490064 13116
rect 154580 12316 154632 12368
rect 320456 12316 320508 12368
rect 156420 12248 156472 12300
rect 326344 12248 326396 12300
rect 156512 12180 156564 12232
rect 330392 12180 330444 12232
rect 156236 12112 156288 12164
rect 331220 12112 331272 12164
rect 156328 12044 156380 12096
rect 332600 12044 332652 12096
rect 156052 11976 156104 12028
rect 337016 11976 337068 12028
rect 158720 11908 158772 11960
rect 365812 11908 365864 11960
rect 160376 11840 160428 11892
rect 386696 11840 386748 11892
rect 102140 11704 102192 11756
rect 130752 11772 130804 11824
rect 161480 11772 161532 11824
rect 398932 11772 398984 11824
rect 126980 11704 127032 11756
rect 128176 11704 128228 11756
rect 168380 11704 168432 11756
rect 492312 11704 492364 11756
rect 99840 10684 99892 10736
rect 130660 10684 130712 10736
rect 153200 10684 153252 10736
rect 298100 10684 298152 10736
rect 106464 10616 106516 10668
rect 138480 10616 138532 10668
rect 153384 10616 153436 10668
rect 299664 10616 299716 10668
rect 92480 10548 92532 10600
rect 130568 10548 130620 10600
rect 153292 10548 153344 10600
rect 303160 10548 303212 10600
rect 85672 10480 85724 10532
rect 130476 10480 130528 10532
rect 157432 10480 157484 10532
rect 353576 10480 353628 10532
rect 75000 10412 75052 10464
rect 134524 10412 134576 10464
rect 157340 10412 157392 10464
rect 349252 10412 349304 10464
rect 349804 10412 349856 10464
rect 583392 10412 583444 10464
rect 67640 10344 67692 10396
rect 131764 10344 131816 10396
rect 180156 10344 180208 10396
rect 440332 10344 440384 10396
rect 71504 10276 71556 10328
rect 135812 10276 135864 10328
rect 166080 10276 166132 10328
rect 456892 10276 456944 10328
rect 151820 9596 151872 9648
rect 281908 9596 281960 9648
rect 151912 9528 151964 9580
rect 285404 9528 285456 9580
rect 155960 9460 156012 9512
rect 332692 9460 332744 9512
rect 156972 9392 157024 9444
rect 336280 9392 336332 9444
rect 160192 9324 160244 9376
rect 382372 9324 382424 9376
rect 160284 9256 160336 9308
rect 385960 9256 386012 9308
rect 160100 9188 160152 9240
rect 389456 9188 389508 9240
rect 57244 9120 57296 9172
rect 134340 9120 134392 9172
rect 164332 9120 164384 9172
rect 436744 9120 436796 9172
rect 53748 9052 53800 9104
rect 134248 9052 134300 9104
rect 165988 9052 166040 9104
rect 453304 9052 453356 9104
rect 50160 8984 50212 9036
rect 134156 8984 134208 9036
rect 165896 8984 165948 9036
rect 459192 8984 459244 9036
rect 38384 8916 38436 8968
rect 132960 8916 133012 8968
rect 171232 8916 171284 8968
rect 525432 8916 525484 8968
rect 150624 8848 150676 8900
rect 264152 8848 264204 8900
rect 150532 8780 150584 8832
rect 258264 8780 258316 8832
rect 177488 8712 177540 8764
rect 267740 8712 267792 8764
rect 123484 8032 123536 8084
rect 139584 8032 139636 8084
rect 110512 7964 110564 8016
rect 129096 7964 129148 8016
rect 111616 7896 111668 7948
rect 138296 7896 138348 7948
rect 109316 7828 109368 7880
rect 138388 7828 138440 7880
rect 337384 7828 337436 7880
rect 581000 7828 581052 7880
rect 102232 7760 102284 7812
rect 138204 7760 138256 7812
rect 176108 7760 176160 7812
rect 426164 7760 426216 7812
rect 95148 7692 95200 7744
rect 137100 7692 137152 7744
rect 165804 7692 165856 7744
rect 455696 7692 455748 7744
rect 66720 7624 66772 7676
rect 135720 7624 135772 7676
rect 169852 7624 169904 7676
rect 469956 7624 470008 7676
rect 31300 7556 31352 7608
rect 132868 7556 132920 7608
rect 167000 7556 167052 7608
rect 471060 7556 471112 7608
rect 129648 6740 129700 6792
rect 189724 6740 189776 6792
rect 92572 6672 92624 6724
rect 132776 6672 132828 6724
rect 147864 6672 147916 6724
rect 228732 6672 228784 6724
rect 87972 6604 88024 6656
rect 137008 6604 137060 6656
rect 149244 6604 149296 6656
rect 239312 6604 239364 6656
rect 77392 6536 77444 6588
rect 135536 6536 135588 6588
rect 149152 6536 149204 6588
rect 242992 6536 243044 6588
rect 73804 6468 73856 6520
rect 135444 6468 135496 6520
rect 149060 6468 149112 6520
rect 246396 6468 246448 6520
rect 56048 6400 56100 6452
rect 134064 6400 134116 6452
rect 149336 6400 149388 6452
rect 249984 6400 250036 6452
rect 52552 6332 52604 6384
rect 134708 6332 134760 6384
rect 150440 6332 150492 6384
rect 260656 6332 260708 6384
rect 40684 6264 40736 6316
rect 132684 6264 132736 6316
rect 165712 6264 165764 6316
rect 450912 6264 450964 6316
rect 24216 6196 24268 6248
rect 131580 6196 131632 6248
rect 142436 6196 142488 6248
rect 155408 6196 155460 6248
rect 165620 6196 165672 6248
rect 460388 6196 460440 6248
rect 23020 6128 23072 6180
rect 131488 6128 131540 6180
rect 144000 6128 144052 6180
rect 170772 6128 170824 6180
rect 176568 6128 176620 6180
rect 578608 6128 578660 6180
rect 126888 5380 126940 5432
rect 133328 5380 133380 5432
rect 104532 5176 104584 5228
rect 139032 5176 139084 5228
rect 143816 5176 143868 5228
rect 173164 5176 173216 5228
rect 20628 5108 20680 5160
rect 43444 5108 43496 5160
rect 70308 5108 70360 5160
rect 136088 5108 136140 5160
rect 143724 5108 143776 5160
rect 174268 5108 174320 5160
rect 431224 5108 431276 5160
rect 475752 5108 475804 5160
rect 28908 5040 28960 5092
rect 126244 5040 126296 5092
rect 164240 5040 164292 5092
rect 443828 5040 443880 5092
rect 33600 4972 33652 5024
rect 133144 4972 133196 5024
rect 142344 4972 142396 5024
rect 151820 4972 151872 5024
rect 170864 4972 170916 5024
rect 508872 4972 508924 5024
rect 21824 4904 21876 4956
rect 131396 4904 131448 4956
rect 142252 4904 142304 4956
rect 157800 4904 157852 4956
rect 171140 4904 171192 4956
rect 533712 4904 533764 4956
rect 14740 4836 14792 4888
rect 131304 4836 131356 4888
rect 143632 4836 143684 4888
rect 167184 4836 167236 4888
rect 173624 4836 173676 4888
rect 551468 4836 551520 4888
rect 13544 4768 13596 4820
rect 131212 4768 131264 4820
rect 143908 4768 143960 4820
rect 169576 4768 169628 4820
rect 174912 4768 174964 4820
rect 566832 4768 566884 4820
rect 18236 4088 18288 4140
rect 131948 4088 132000 4140
rect 140964 4088 141016 4140
rect 144736 4088 144788 4140
rect 146300 4088 146352 4140
rect 201500 4088 201552 4140
rect 202696 4088 202748 4140
rect 207388 4088 207440 4140
rect 125876 4020 125928 4072
rect 139952 4020 140004 4072
rect 146392 4020 146444 4072
rect 210976 4020 211028 4072
rect 90364 3952 90416 4004
rect 137376 3952 137428 4004
rect 147772 3952 147824 4004
rect 221556 3952 221608 4004
rect 251180 3952 251232 4004
rect 252376 3952 252428 4004
rect 86868 3884 86920 3936
rect 137284 3884 137336 3936
rect 170680 3884 170732 3936
rect 349160 3884 349212 3936
rect 349896 3884 349948 3936
rect 545488 3884 545540 3936
rect 72608 3816 72660 3868
rect 130384 3816 130436 3868
rect 141056 3816 141108 3868
rect 147128 3816 147180 3868
rect 148600 3816 148652 3868
rect 225144 3816 225196 3868
rect 228364 3816 228416 3868
rect 469864 3816 469916 3868
rect 469956 3816 470008 3868
rect 504180 3816 504232 3868
rect 76196 3748 76248 3800
rect 135996 3748 136048 3800
rect 142160 3748 142212 3800
rect 154212 3748 154264 3800
rect 159364 3748 159416 3800
rect 180248 3748 180300 3800
rect 185584 3748 185636 3800
rect 472256 3748 472308 3800
rect 32404 3680 32456 3732
rect 92572 3680 92624 3732
rect 93952 3680 94004 3732
rect 136824 3680 136876 3732
rect 141240 3680 141292 3732
rect 142436 3680 142488 3732
rect 144460 3680 144512 3732
rect 160100 3680 160152 3732
rect 176016 3680 176068 3732
rect 465172 3680 465224 3732
rect 465724 3680 465776 3732
rect 549076 3680 549128 3732
rect 59636 3612 59688 3664
rect 120724 3612 120776 3664
rect 144184 3612 144236 3664
rect 164884 3612 164936 3664
rect 177396 3612 177448 3664
rect 494704 3612 494756 3664
rect 46664 3544 46716 3596
rect 129004 3544 129056 3596
rect 136456 3544 136508 3596
rect 140228 3544 140280 3596
rect 141608 3544 141660 3596
rect 143540 3544 143592 3596
rect 146024 3544 146076 3596
rect 2780 3476 2832 3528
rect 3700 3476 3752 3528
rect 11152 3476 11204 3528
rect 13084 3476 13136 3528
rect 37188 3476 37240 3528
rect 126888 3476 126940 3528
rect 140044 3476 140096 3528
rect 141148 3476 141200 3528
rect 144276 3476 144328 3528
rect 149520 3476 149572 3528
rect 151084 3544 151136 3596
rect 153016 3544 153068 3596
rect 156420 3544 156472 3596
rect 171968 3544 172020 3596
rect 177304 3544 177356 3596
rect 505376 3544 505428 3596
rect 168380 3476 168432 3528
rect 170404 3476 170456 3528
rect 501788 3476 501840 3528
rect 506480 3476 506532 3528
rect 507308 3476 507360 3528
rect 531320 3476 531372 3528
rect 532148 3476 532200 3528
rect 539600 3476 539652 3528
rect 540428 3476 540480 3528
rect 564440 3476 564492 3528
rect 565268 3476 565320 3528
rect 5264 3408 5316 3460
rect 10324 3408 10376 3460
rect 102140 3408 102192 3460
rect 103336 3408 103388 3460
rect 131764 3408 131816 3460
rect 139952 3408 140004 3460
rect 144552 3408 144604 3460
rect 176660 3408 176712 3460
rect 177948 3408 178000 3460
rect 523040 3408 523092 3460
rect 122288 3340 122340 3392
rect 139768 3340 139820 3392
rect 145656 3340 145708 3392
rect 142896 3272 142948 3324
rect 145932 3272 145984 3324
rect 151268 3340 151320 3392
rect 203892 3340 203944 3392
rect 242900 3340 242952 3392
rect 244096 3340 244148 3392
rect 299480 3340 299532 3392
rect 300768 3340 300820 3392
rect 307760 3340 307812 3392
rect 309048 3340 309100 3392
rect 316040 3340 316092 3392
rect 317328 3340 317380 3392
rect 324320 3340 324372 3392
rect 325608 3340 325660 3392
rect 332600 3340 332652 3392
rect 333888 3340 333940 3392
rect 340880 3340 340932 3392
rect 342168 3340 342220 3392
rect 349252 3340 349304 3392
rect 350448 3340 350500 3392
rect 357440 3340 357492 3392
rect 358728 3340 358780 3392
rect 374092 3340 374144 3392
rect 375288 3340 375340 3392
rect 382280 3340 382332 3392
rect 383568 3340 383620 3392
rect 390560 3340 390612 3392
rect 391848 3340 391900 3392
rect 398932 3340 398984 3392
rect 400128 3340 400180 3392
rect 407120 3340 407172 3392
rect 408408 3340 408460 3392
rect 415400 3340 415452 3392
rect 416688 3340 416740 3392
rect 423772 3340 423824 3392
rect 424968 3340 425020 3392
rect 432052 3340 432104 3392
rect 433248 3340 433300 3392
rect 456800 3340 456852 3392
rect 458088 3340 458140 3392
rect 481640 3340 481692 3392
rect 482468 3340 482520 3392
rect 489920 3340 489972 3392
rect 490748 3340 490800 3392
rect 156420 3272 156472 3324
rect 178684 3272 178736 3324
rect 197912 3272 197964 3324
rect 202144 3272 202196 3324
rect 245200 3272 245252 3324
rect 448520 3272 448572 3324
rect 449808 3272 449860 3324
rect 142804 3204 142856 3256
rect 148324 3204 148376 3256
rect 153844 3204 153896 3256
rect 158904 3204 158956 3256
rect 180064 3204 180116 3256
rect 219256 3204 219308 3256
rect 177672 3136 177724 3188
rect 186136 3136 186188 3188
rect 132960 3068 133012 3120
rect 140136 3068 140188 3120
rect 145564 2932 145616 2984
rect 150624 2932 150676 2984
rect 365720 1232 365772 1284
rect 367008 1232 367060 1284
rect 440240 552 440292 604
rect 441528 552 441580 604
<< metal2 >>
rect 6932 703582 7972 703610
rect 2778 684312 2834 684321
rect 2778 684247 2834 684256
rect 2792 683670 2820 684247
rect 2780 683664 2832 683670
rect 2780 683606 2832 683612
rect 6184 683664 6236 683670
rect 6184 683606 6236 683612
rect 3422 671256 3478 671265
rect 3422 671191 3478 671200
rect 3436 670818 3464 671191
rect 3424 670812 3476 670818
rect 3424 670754 3476 670760
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 2780 632120 2832 632126
rect 2778 632088 2780 632097
rect 2832 632088 2834 632097
rect 2778 632023 2834 632032
rect 3146 580000 3202 580009
rect 3146 579935 3202 579944
rect 3160 579834 3188 579935
rect 3148 579828 3200 579834
rect 3148 579770 3200 579776
rect 3054 566944 3110 566953
rect 3054 566879 3110 566888
rect 3068 565894 3096 566879
rect 3056 565888 3108 565894
rect 3056 565830 3108 565836
rect 3330 553888 3386 553897
rect 3330 553823 3386 553832
rect 3344 553450 3372 553823
rect 3332 553444 3384 553450
rect 3332 553386 3384 553392
rect 2962 527912 3018 527921
rect 2962 527847 3018 527856
rect 2976 527202 3004 527847
rect 2964 527196 3016 527202
rect 2964 527138 3016 527144
rect 3330 475688 3386 475697
rect 3330 475623 3386 475632
rect 3344 474774 3372 475623
rect 3332 474768 3384 474774
rect 3332 474710 3384 474716
rect 2962 423600 3018 423609
rect 2962 423535 3018 423544
rect 2976 422346 3004 423535
rect 2964 422340 3016 422346
rect 2964 422282 3016 422288
rect 3330 410544 3386 410553
rect 3330 410479 3386 410488
rect 3344 409902 3372 410479
rect 3332 409896 3384 409902
rect 3332 409838 3384 409844
rect 3330 371376 3386 371385
rect 3330 371311 3386 371320
rect 3344 371278 3372 371311
rect 3332 371272 3384 371278
rect 3332 371214 3384 371220
rect 3330 358456 3386 358465
rect 3330 358391 3386 358400
rect 3344 357474 3372 358391
rect 3332 357468 3384 357474
rect 3332 357410 3384 357416
rect 3330 345400 3386 345409
rect 3330 345335 3386 345344
rect 3344 345098 3372 345335
rect 3332 345092 3384 345098
rect 3332 345034 3384 345040
rect 2778 319288 2834 319297
rect 2778 319223 2834 319232
rect 2792 319122 2820 319223
rect 2780 319116 2832 319122
rect 2780 319058 2832 319064
rect 2870 306232 2926 306241
rect 2870 306167 2926 306176
rect 2884 305046 2912 306167
rect 2872 305040 2924 305046
rect 2872 304982 2924 304988
rect 3330 293176 3386 293185
rect 3330 293111 3386 293120
rect 3344 292602 3372 293111
rect 3332 292596 3384 292602
rect 3332 292538 3384 292544
rect 3238 267200 3294 267209
rect 3238 267135 3294 267144
rect 3252 266422 3280 267135
rect 3240 266416 3292 266422
rect 3240 266358 3292 266364
rect 2870 254144 2926 254153
rect 2870 254079 2926 254088
rect 2884 253978 2912 254079
rect 2872 253972 2924 253978
rect 2872 253914 2924 253920
rect 3238 241088 3294 241097
rect 3238 241023 3294 241032
rect 3252 240174 3280 241023
rect 3240 240168 3292 240174
rect 3240 240110 3292 240116
rect 3330 214976 3386 214985
rect 3330 214911 3386 214920
rect 3344 213994 3372 214911
rect 3332 213988 3384 213994
rect 3332 213930 3384 213936
rect 3330 201920 3386 201929
rect 3330 201855 3386 201864
rect 3344 201550 3372 201855
rect 3332 201544 3384 201550
rect 3332 201486 3384 201492
rect 3332 162920 3384 162926
rect 3330 162888 3332 162897
rect 3384 162888 3386 162897
rect 3330 162823 3386 162832
rect 3330 149832 3386 149841
rect 3330 149767 3386 149776
rect 3344 149122 3372 149767
rect 3332 149116 3384 149122
rect 3332 149058 3384 149064
rect 2778 136776 2834 136785
rect 2778 136711 2780 136720
rect 2832 136711 2834 136720
rect 2780 136682 2832 136688
rect 3332 111784 3384 111790
rect 3332 111726 3384 111732
rect 3344 110673 3372 111726
rect 3330 110664 3386 110673
rect 3330 110599 3386 110608
rect 3436 79121 3464 658135
rect 4804 632120 4856 632126
rect 4804 632062 4856 632068
rect 3514 619168 3570 619177
rect 3514 619103 3570 619112
rect 3528 618322 3556 619103
rect 3516 618316 3568 618322
rect 3516 618258 3568 618264
rect 3606 606112 3662 606121
rect 3606 606047 3662 606056
rect 3514 501800 3570 501809
rect 3514 501735 3570 501744
rect 3422 79112 3478 79121
rect 3422 79047 3478 79056
rect 3528 78878 3556 501735
rect 3620 79257 3648 606047
rect 3698 514856 3754 514865
rect 3698 514791 3754 514800
rect 3712 144226 3740 514791
rect 3974 462632 4030 462641
rect 3974 462567 4030 462576
rect 3790 449576 3846 449585
rect 3790 449511 3846 449520
rect 3700 144220 3752 144226
rect 3700 144162 3752 144168
rect 3700 138032 3752 138038
rect 3700 137974 3752 137980
rect 3712 97617 3740 137974
rect 3698 97608 3754 97617
rect 3698 97543 3754 97552
rect 3698 84688 3754 84697
rect 3698 84623 3754 84632
rect 3712 80714 3740 84623
rect 3700 80708 3752 80714
rect 3700 80650 3752 80656
rect 3606 79248 3662 79257
rect 3606 79183 3662 79192
rect 3804 79014 3832 449511
rect 3882 397488 3938 397497
rect 3882 397423 3938 397432
rect 3896 79354 3924 397423
rect 3988 148374 4016 462567
rect 4066 188864 4122 188873
rect 4066 188799 4122 188808
rect 3976 148368 4028 148374
rect 3976 148310 4028 148316
rect 4080 79422 4108 188799
rect 4816 120086 4844 632062
rect 4896 319116 4948 319122
rect 4896 319058 4948 319064
rect 4908 129742 4936 319058
rect 4988 136740 5040 136746
rect 4988 136682 5040 136688
rect 4896 129736 4948 129742
rect 4896 129678 4948 129684
rect 4804 120080 4856 120086
rect 4804 120022 4856 120028
rect 5000 80850 5028 136682
rect 6196 118658 6224 683606
rect 6184 118652 6236 118658
rect 6184 118594 6236 118600
rect 4988 80844 5040 80850
rect 4988 80786 5040 80792
rect 4068 79416 4120 79422
rect 6932 79393 6960 703582
rect 7944 703474 7972 703582
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 8128 703474 8156 703520
rect 7944 703446 8156 703474
rect 24320 700330 24348 703520
rect 24308 700324 24360 700330
rect 24308 700266 24360 700272
rect 7564 579828 7616 579834
rect 7564 579770 7616 579776
rect 7576 121446 7604 579770
rect 15844 527196 15896 527202
rect 15844 527138 15896 527144
rect 15856 122806 15884 527138
rect 19984 474768 20036 474774
rect 19984 474710 20036 474716
rect 19996 124166 20024 474710
rect 22744 422340 22796 422346
rect 22744 422282 22796 422288
rect 21364 133952 21416 133958
rect 21364 133894 21416 133900
rect 19984 124160 20036 124166
rect 19984 124102 20036 124108
rect 15844 122800 15896 122806
rect 15844 122742 15896 122748
rect 7564 121440 7616 121446
rect 7564 121382 7616 121388
rect 21376 111790 21404 133894
rect 22756 126954 22784 422282
rect 22836 371272 22888 371278
rect 22836 371214 22888 371220
rect 22848 128314 22876 371214
rect 22928 266416 22980 266422
rect 22928 266358 22980 266364
rect 22940 131102 22968 266358
rect 24124 213988 24176 213994
rect 24124 213930 24176 213936
rect 23020 136672 23072 136678
rect 23020 136614 23072 136620
rect 22928 131096 22980 131102
rect 22928 131038 22980 131044
rect 22836 128308 22888 128314
rect 22836 128250 22888 128256
rect 22744 126948 22796 126954
rect 22744 126890 22796 126896
rect 21364 111784 21416 111790
rect 21364 111726 21416 111732
rect 4068 79358 4120 79364
rect 6918 79384 6974 79393
rect 3884 79348 3936 79354
rect 6918 79319 6974 79328
rect 3884 79290 3936 79296
rect 3792 79008 3844 79014
rect 3792 78950 3844 78956
rect 3516 78872 3568 78878
rect 3516 78814 3568 78820
rect 10324 78124 10376 78130
rect 10324 78066 10376 78072
rect 2780 77988 2832 77994
rect 2780 77930 2832 77936
rect 1400 75200 1452 75206
rect 1400 75142 1452 75148
rect 20 72480 72 72486
rect 20 72422 72 72428
rect 32 16574 60 72422
rect 32 16546 152 16574
rect 124 354 152 16546
rect 542 354 654 480
rect 124 326 654 354
rect 1412 354 1440 75142
rect 2792 3534 2820 77930
rect 6918 75168 6974 75177
rect 6918 75103 6974 75112
rect 2872 73840 2924 73846
rect 2872 73782 2924 73788
rect 2780 3528 2832 3534
rect 2780 3470 2832 3476
rect 2884 480 2912 73782
rect 3424 71732 3476 71738
rect 3424 71674 3476 71680
rect 3436 71641 3464 71674
rect 3422 71632 3478 71641
rect 3422 71567 3478 71576
rect 5540 69692 5592 69698
rect 5540 69634 5592 69640
rect 3516 65816 3568 65822
rect 3516 65758 3568 65764
rect 3528 58585 3556 65758
rect 3514 58576 3570 58585
rect 3514 58511 3570 58520
rect 3424 45552 3476 45558
rect 3422 45520 3424 45529
rect 3476 45520 3478 45529
rect 3422 45455 3478 45464
rect 3516 33108 3568 33114
rect 3516 33050 3568 33056
rect 3424 32700 3476 32706
rect 3424 32642 3476 32648
rect 3240 23044 3292 23050
rect 3240 22986 3292 22992
rect 3252 19417 3280 22986
rect 3238 19408 3294 19417
rect 3238 19343 3294 19352
rect 3436 6497 3464 32642
rect 3528 32473 3556 33050
rect 3514 32464 3570 32473
rect 3514 32399 3570 32408
rect 5552 16574 5580 69634
rect 6932 16574 6960 75103
rect 5552 16546 6040 16574
rect 6932 16546 7696 16574
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 3700 3528 3752 3534
rect 3700 3470 3752 3476
rect 1646 354 1758 480
rect 1412 326 1758 354
rect 542 -960 654 326
rect 1646 -960 1758 326
rect 2842 -960 2954 480
rect 3712 354 3740 3470
rect 5264 3460 5316 3466
rect 5264 3402 5316 3408
rect 5276 480 5304 3402
rect 4038 354 4150 480
rect 3712 326 4150 354
rect 4038 -960 4150 326
rect 5234 -960 5346 480
rect 6012 354 6040 16546
rect 7668 480 7696 16546
rect 9954 8936 10010 8945
rect 9954 8871 10010 8880
rect 8758 4856 8814 4865
rect 8758 4791 8814 4800
rect 8772 480 8800 4791
rect 9968 480 9996 8871
rect 10336 3466 10364 78066
rect 13082 77888 13138 77897
rect 13082 77823 13138 77832
rect 11058 76528 11114 76537
rect 11058 76463 11114 76472
rect 11072 16574 11100 76463
rect 11072 16546 11928 16574
rect 11152 3528 11204 3534
rect 11152 3470 11204 3476
rect 10324 3460 10376 3466
rect 10324 3402 10376 3408
rect 11164 480 11192 3470
rect 6430 354 6542 480
rect 6012 326 6542 354
rect 6430 -960 6542 326
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 11900 354 11928 16546
rect 13096 3534 13124 77823
rect 16580 73908 16632 73914
rect 16580 73850 16632 73856
rect 15200 18624 15252 18630
rect 15200 18566 15252 18572
rect 15212 16574 15240 18566
rect 16592 16574 16620 73850
rect 19340 39364 19392 39370
rect 19340 39306 19392 39312
rect 19352 16574 19380 39306
rect 23032 33114 23060 136614
rect 24136 132462 24164 213930
rect 29644 162920 29696 162926
rect 29644 162862 29696 162868
rect 24216 135312 24268 135318
rect 24216 135254 24268 135260
rect 24124 132456 24176 132462
rect 24124 132398 24176 132404
rect 24228 71738 24256 135254
rect 29656 133890 29684 162862
rect 29644 133884 29696 133890
rect 29644 133826 29696 133832
rect 40052 117298 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 234632 703582 235028 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 700398 73016 703520
rect 89180 702434 89208 703520
rect 88352 702406 89208 702434
rect 72976 700392 73028 700398
rect 72976 700334 73028 700340
rect 79324 292596 79376 292602
rect 79324 292538 79376 292544
rect 40040 117292 40092 117298
rect 40040 117234 40092 117240
rect 79336 79490 79364 292538
rect 88352 142934 88380 702406
rect 105464 699718 105492 703520
rect 137848 700398 137876 703520
rect 154132 700466 154160 703520
rect 170324 702434 170352 703520
rect 202800 703050 202828 703520
rect 201500 703044 201552 703050
rect 201500 702986 201552 702992
rect 202788 703044 202840 703050
rect 202788 702986 202840 702992
rect 169772 702406 170352 702434
rect 154120 700460 154172 700466
rect 154120 700402 154172 700408
rect 119344 700392 119396 700398
rect 119344 700334 119396 700340
rect 137836 700392 137888 700398
rect 137836 700334 137888 700340
rect 105452 699712 105504 699718
rect 105452 699654 105504 699660
rect 106924 699712 106976 699718
rect 106924 699654 106976 699660
rect 88340 142928 88392 142934
rect 88340 142870 88392 142876
rect 106936 115938 106964 699654
rect 118700 616888 118752 616894
rect 118700 616830 118752 616836
rect 116584 553444 116636 553450
rect 116584 553386 116636 553392
rect 106924 115932 106976 115938
rect 106924 115874 106976 115880
rect 116596 79830 116624 553386
rect 118608 404388 118660 404394
rect 118608 404330 118660 404336
rect 118516 351960 118568 351966
rect 118516 351902 118568 351908
rect 116676 345092 116728 345098
rect 116676 345034 116728 345040
rect 116584 79824 116636 79830
rect 116584 79766 116636 79772
rect 116688 79558 116716 345034
rect 118424 239420 118476 239426
rect 118424 239362 118476 239368
rect 118332 202156 118384 202162
rect 118332 202098 118384 202104
rect 118240 142860 118292 142866
rect 118240 142802 118292 142808
rect 118056 141500 118108 141506
rect 118056 141442 118108 141448
rect 117318 137592 117374 137601
rect 117318 137527 117374 137536
rect 117332 136678 117360 137527
rect 117320 136672 117372 136678
rect 117320 136614 117372 136620
rect 117318 136096 117374 136105
rect 117318 136031 117374 136040
rect 117332 135318 117360 136031
rect 117320 135312 117372 135318
rect 117320 135254 117372 135260
rect 117318 134600 117374 134609
rect 117318 134535 117374 134544
rect 117332 133958 117360 134535
rect 117320 133952 117372 133958
rect 117320 133894 117372 133900
rect 117412 133884 117464 133890
rect 117412 133826 117464 133832
rect 117424 133113 117452 133826
rect 117410 133104 117466 133113
rect 117410 133039 117466 133048
rect 117320 132456 117372 132462
rect 117320 132398 117372 132404
rect 117332 131617 117360 132398
rect 117318 131608 117374 131617
rect 117318 131543 117374 131552
rect 117320 131096 117372 131102
rect 117320 131038 117372 131044
rect 117332 130121 117360 131038
rect 117318 130112 117374 130121
rect 117318 130047 117374 130056
rect 117320 129736 117372 129742
rect 117320 129678 117372 129684
rect 117332 128625 117360 129678
rect 117318 128616 117374 128625
rect 117318 128551 117374 128560
rect 117320 128308 117372 128314
rect 117320 128250 117372 128256
rect 117332 127129 117360 128250
rect 117318 127120 117374 127129
rect 117318 127055 117374 127064
rect 117320 126948 117372 126954
rect 117320 126890 117372 126896
rect 117332 125633 117360 126890
rect 117318 125624 117374 125633
rect 117318 125559 117374 125568
rect 117320 124160 117372 124166
rect 117318 124128 117320 124137
rect 117372 124128 117374 124137
rect 117318 124063 117374 124072
rect 117320 122800 117372 122806
rect 117320 122742 117372 122748
rect 117332 122641 117360 122742
rect 117318 122632 117374 122641
rect 117318 122567 117374 122576
rect 117320 121440 117372 121446
rect 117320 121382 117372 121388
rect 117332 121145 117360 121382
rect 117318 121136 117374 121145
rect 117318 121071 117374 121080
rect 117320 120080 117372 120086
rect 117320 120022 117372 120028
rect 117332 119649 117360 120022
rect 117318 119640 117374 119649
rect 117318 119575 117374 119584
rect 117320 118652 117372 118658
rect 117320 118594 117372 118600
rect 117332 118153 117360 118594
rect 117318 118144 117374 118153
rect 117318 118079 117374 118088
rect 117320 117292 117372 117298
rect 117320 117234 117372 117240
rect 117332 116657 117360 117234
rect 117318 116648 117374 116657
rect 117318 116583 117374 116592
rect 117320 115932 117372 115938
rect 117320 115874 117372 115880
rect 117332 115161 117360 115874
rect 117318 115152 117374 115161
rect 117318 115087 117374 115096
rect 118068 113665 118096 141442
rect 118148 139460 118200 139466
rect 118148 139402 118200 139408
rect 118054 113656 118110 113665
rect 118054 113591 118110 113600
rect 118160 88233 118188 139402
rect 118252 89729 118280 142802
rect 118344 91225 118372 202098
rect 118436 92721 118464 239362
rect 118528 94217 118556 351902
rect 118620 95713 118648 404330
rect 118712 101697 118740 616830
rect 118792 275324 118844 275330
rect 118792 275266 118844 275272
rect 118804 112169 118832 275266
rect 118884 149728 118936 149734
rect 118884 149670 118936 149676
rect 118790 112160 118846 112169
rect 118790 112095 118846 112104
rect 118896 110673 118924 149670
rect 119160 141432 119212 141438
rect 119160 141374 119212 141380
rect 119068 140140 119120 140146
rect 119068 140082 119120 140088
rect 118976 140072 119028 140078
rect 118976 140014 119028 140020
rect 118882 110664 118938 110673
rect 118882 110599 118938 110608
rect 118988 104689 119016 140014
rect 119080 106185 119108 140082
rect 119172 107681 119200 141374
rect 119252 140208 119304 140214
rect 119252 140150 119304 140156
rect 119264 109177 119292 140150
rect 119250 109168 119306 109177
rect 119250 109103 119306 109112
rect 119158 107672 119214 107681
rect 119158 107607 119214 107616
rect 119066 106176 119122 106185
rect 119066 106111 119122 106120
rect 118974 104680 119030 104689
rect 118974 104615 119030 104624
rect 118698 101688 118754 101697
rect 118698 101623 118754 101632
rect 118606 95704 118662 95713
rect 118606 95639 118662 95648
rect 118514 94208 118570 94217
rect 118514 94143 118570 94152
rect 118422 92712 118478 92721
rect 118422 92647 118478 92656
rect 118330 91216 118386 91225
rect 118330 91151 118386 91160
rect 118238 89720 118294 89729
rect 118238 89655 118294 89664
rect 118146 88224 118202 88233
rect 118146 88159 118202 88168
rect 118422 86728 118478 86737
rect 118422 86663 118478 86672
rect 118330 82240 118386 82249
rect 118330 82175 118386 82184
rect 116676 79552 116728 79558
rect 116676 79494 116728 79500
rect 79324 79484 79376 79490
rect 79324 79426 79376 79432
rect 96620 78260 96672 78266
rect 96620 78202 96672 78208
rect 78680 78192 78732 78198
rect 78680 78134 78732 78140
rect 43444 78056 43496 78062
rect 43444 77998 43496 78004
rect 41420 76628 41472 76634
rect 41420 76570 41472 76576
rect 34520 76560 34572 76566
rect 34520 76502 34572 76508
rect 29000 73976 29052 73982
rect 29000 73918 29052 73924
rect 26238 73808 26294 73817
rect 26238 73743 26294 73752
rect 24216 71732 24268 71738
rect 24216 71674 24268 71680
rect 23020 33108 23072 33114
rect 23020 33050 23072 33056
rect 15212 16546 15976 16574
rect 16592 16546 17080 16574
rect 19352 16546 19472 16574
rect 14740 4888 14792 4894
rect 14740 4830 14792 4836
rect 13544 4820 13596 4826
rect 13544 4762 13596 4768
rect 13084 3528 13136 3534
rect 13084 3470 13136 3476
rect 13556 480 13584 4762
rect 14752 480 14780 4830
rect 15948 480 15976 16546
rect 17052 480 17080 16546
rect 18236 4140 18288 4146
rect 18236 4082 18288 4088
rect 18248 480 18276 4082
rect 19444 480 19472 16546
rect 25318 9072 25374 9081
rect 25318 9007 25374 9016
rect 24216 6248 24268 6254
rect 24216 6190 24268 6196
rect 23020 6180 23072 6186
rect 23020 6122 23072 6128
rect 20628 5160 20680 5166
rect 20628 5102 20680 5108
rect 20640 480 20668 5102
rect 21824 4956 21876 4962
rect 21824 4898 21876 4904
rect 21836 480 21864 4898
rect 23032 480 23060 6122
rect 24228 480 24256 6190
rect 25332 480 25360 9007
rect 12318 354 12430 480
rect 11900 326 12430 354
rect 12318 -960 12430 326
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 73743
rect 29012 16574 29040 73918
rect 29012 16546 30144 16574
rect 27710 7576 27766 7585
rect 27710 7511 27766 7520
rect 27724 480 27752 7511
rect 28908 5092 28960 5098
rect 28908 5034 28960 5040
rect 28920 480 28948 5034
rect 30116 480 30144 16546
rect 31300 7608 31352 7614
rect 31300 7550 31352 7556
rect 31312 480 31340 7550
rect 33600 5024 33652 5030
rect 33600 4966 33652 4972
rect 32404 3732 32456 3738
rect 32404 3674 32456 3680
rect 32416 480 32444 3674
rect 33612 480 33640 4966
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34532 354 34560 76502
rect 38660 44872 38712 44878
rect 38660 44814 38712 44820
rect 35900 18692 35952 18698
rect 35900 18634 35952 18640
rect 35912 16574 35940 18634
rect 38672 16574 38700 44814
rect 41432 16574 41460 76570
rect 42800 57248 42852 57254
rect 42800 57190 42852 57196
rect 35912 16546 36032 16574
rect 38672 16546 39160 16574
rect 41432 16546 41920 16574
rect 36004 480 36032 16546
rect 38384 8968 38436 8974
rect 38384 8910 38436 8916
rect 37188 3528 37240 3534
rect 37188 3470 37240 3476
rect 37200 480 37228 3470
rect 38396 480 38424 8910
rect 34766 354 34878 480
rect 34532 326 34878 354
rect 34766 -960 34878 326
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39132 354 39160 16546
rect 40684 6316 40736 6322
rect 40684 6258 40736 6264
rect 40696 480 40724 6258
rect 41892 480 41920 16546
rect 39550 354 39662 480
rect 39132 326 39662 354
rect 39550 -960 39662 326
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 42812 354 42840 57190
rect 43456 5166 43484 77998
rect 60738 75440 60794 75449
rect 60738 75375 60794 75384
rect 69020 75404 69072 75410
rect 51080 75336 51132 75342
rect 44178 75304 44234 75313
rect 51080 75278 51132 75284
rect 44178 75239 44234 75248
rect 46940 75268 46992 75274
rect 44192 16574 44220 75239
rect 46940 75210 46992 75216
rect 46952 16574 46980 75210
rect 48318 73944 48374 73953
rect 48318 73879 48374 73888
rect 48332 16574 48360 73879
rect 44192 16546 44312 16574
rect 46952 16546 47440 16574
rect 48332 16546 48544 16574
rect 43444 5160 43496 5166
rect 43444 5102 43496 5108
rect 44284 480 44312 16546
rect 45466 9208 45522 9217
rect 45466 9143 45522 9152
rect 45480 480 45508 9143
rect 46664 3596 46716 3602
rect 46664 3538 46716 3544
rect 46676 480 46704 3538
rect 43046 354 43158 480
rect 42812 326 43158 354
rect 43046 -960 43158 326
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47412 354 47440 16546
rect 47830 354 47942 480
rect 47412 326 47942 354
rect 48516 354 48544 16546
rect 50160 9036 50212 9042
rect 50160 8978 50212 8984
rect 50172 480 50200 8978
rect 48934 354 49046 480
rect 48516 326 49046 354
rect 47830 -960 47942 326
rect 48934 -960 49046 326
rect 50130 -960 50242 480
rect 51092 354 51120 75278
rect 57980 72548 58032 72554
rect 57980 72490 58032 72496
rect 53840 71052 53892 71058
rect 53840 70994 53892 71000
rect 53852 16574 53880 70994
rect 57992 16574 58020 72490
rect 60752 16574 60780 75375
rect 69020 75346 69072 75352
rect 64880 74044 64932 74050
rect 64880 73986 64932 73992
rect 63498 22672 63554 22681
rect 63498 22607 63554 22616
rect 63512 16574 63540 22607
rect 64892 16574 64920 73986
rect 69032 16574 69060 75346
rect 78692 16574 78720 78134
rect 91100 76832 91152 76838
rect 91100 76774 91152 76780
rect 84200 76696 84252 76702
rect 80058 76664 80114 76673
rect 84200 76638 84252 76644
rect 80058 76599 80114 76608
rect 80072 16574 80100 76599
rect 81440 75472 81492 75478
rect 81440 75414 81492 75420
rect 81452 16574 81480 75414
rect 82820 74112 82872 74118
rect 82820 74054 82872 74060
rect 82832 16574 82860 74054
rect 53852 16546 54984 16574
rect 57992 16546 58480 16574
rect 60752 16546 61608 16574
rect 63512 16546 64368 16574
rect 64892 16546 65104 16574
rect 69032 16546 69152 16574
rect 78692 16546 79272 16574
rect 80072 16546 80928 16574
rect 81452 16546 81664 16574
rect 82832 16546 83320 16574
rect 53748 9104 53800 9110
rect 53748 9046 53800 9052
rect 52552 6384 52604 6390
rect 52552 6326 52604 6332
rect 52564 480 52592 6326
rect 53760 480 53788 9046
rect 54956 480 54984 16546
rect 57244 9172 57296 9178
rect 57244 9114 57296 9120
rect 56048 6452 56100 6458
rect 56048 6394 56100 6400
rect 56060 480 56088 6394
rect 57256 480 57284 9114
rect 58452 480 58480 16546
rect 60830 9344 60886 9353
rect 60830 9279 60886 9288
rect 59636 3664 59688 3670
rect 59636 3606 59688 3612
rect 59648 480 59676 3606
rect 60844 480 60872 9279
rect 51326 354 51438 480
rect 51092 326 51438 354
rect 51326 -960 51438 326
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61580 354 61608 16546
rect 63222 6216 63278 6225
rect 63222 6151 63278 6160
rect 63236 480 63264 6151
rect 64340 480 64368 16546
rect 61998 354 62110 480
rect 61580 326 62110 354
rect 61998 -960 62110 326
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65076 354 65104 16546
rect 67640 10396 67692 10402
rect 67640 10338 67692 10344
rect 66720 7676 66772 7682
rect 66720 7618 66772 7624
rect 66732 480 66760 7618
rect 65494 354 65606 480
rect 65076 326 65606 354
rect 65494 -960 65606 326
rect 66690 -960 66802 480
rect 67652 354 67680 10338
rect 69124 480 69152 16546
rect 75000 10464 75052 10470
rect 75000 10406 75052 10412
rect 71504 10328 71556 10334
rect 71504 10270 71556 10276
rect 70308 5160 70360 5166
rect 70308 5102 70360 5108
rect 70320 480 70348 5102
rect 71516 480 71544 10270
rect 73804 6520 73856 6526
rect 73804 6462 73856 6468
rect 72608 3868 72660 3874
rect 72608 3810 72660 3816
rect 72620 480 72648 3810
rect 73816 480 73844 6462
rect 75012 480 75040 10406
rect 78586 9480 78642 9489
rect 78586 9415 78642 9424
rect 77392 6588 77444 6594
rect 77392 6530 77444 6536
rect 76196 3800 76248 3806
rect 76196 3742 76248 3748
rect 76208 480 76236 3742
rect 77404 480 77432 6530
rect 78600 480 78628 9415
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79244 354 79272 16546
rect 80900 480 80928 16546
rect 79662 354 79774 480
rect 79244 326 79774 354
rect 79662 -960 79774 326
rect 80858 -960 80970 480
rect 81636 354 81664 16546
rect 83292 480 83320 16546
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84212 354 84240 76638
rect 88340 22840 88392 22846
rect 88340 22782 88392 22788
rect 88352 16574 88380 22782
rect 91112 16574 91140 76774
rect 95238 21312 95294 21321
rect 95238 21247 95294 21256
rect 95252 16574 95280 21247
rect 96632 16574 96660 78202
rect 115938 76936 115994 76945
rect 115938 76871 115994 76880
rect 97998 76800 98054 76809
rect 97998 76735 98054 76744
rect 104900 76764 104952 76770
rect 98012 16574 98040 76735
rect 104900 76706 104952 76712
rect 104912 16574 104940 76706
rect 114560 74180 114612 74186
rect 114560 74122 114612 74128
rect 107660 72616 107712 72622
rect 107660 72558 107712 72564
rect 107672 16574 107700 72558
rect 111800 18760 111852 18766
rect 111800 18702 111852 18708
rect 111812 16574 111840 18702
rect 114572 16574 114600 74122
rect 115952 16574 115980 76871
rect 118344 22778 118372 82175
rect 118436 81161 118464 86663
rect 118606 85232 118662 85241
rect 118606 85167 118662 85176
rect 118514 83736 118570 83745
rect 118514 83671 118570 83680
rect 118422 81152 118478 81161
rect 118422 81087 118478 81096
rect 118528 46918 118556 83671
rect 118620 80986 118648 85167
rect 118608 80980 118660 80986
rect 118608 80922 118660 80928
rect 119356 78849 119384 700334
rect 120724 670744 120776 670750
rect 120724 670686 120776 670692
rect 119436 240168 119488 240174
rect 119436 240110 119488 240116
rect 119342 78840 119398 78849
rect 119342 78775 119398 78784
rect 119448 78577 119476 240110
rect 120736 103465 120764 670686
rect 120816 563100 120868 563106
rect 120816 563042 120868 563048
rect 120722 103456 120778 103465
rect 120722 103391 120778 103400
rect 120828 100745 120856 563042
rect 120908 510672 120960 510678
rect 120908 510614 120960 510620
rect 120814 100736 120870 100745
rect 120814 100671 120870 100680
rect 120920 98705 120948 510614
rect 121000 456816 121052 456822
rect 121000 456758 121052 456764
rect 120906 98696 120962 98705
rect 120906 98631 120962 98640
rect 121012 97209 121040 456758
rect 122104 165640 122156 165646
rect 122104 165582 122156 165588
rect 122116 139466 122144 165582
rect 169772 141506 169800 702406
rect 189080 700460 189132 700466
rect 189080 700402 189132 700408
rect 200764 700460 200816 700466
rect 200764 700402 200816 700408
rect 188344 305040 188396 305046
rect 188344 304982 188396 304988
rect 169760 141500 169812 141506
rect 169760 141442 169812 141448
rect 122104 139460 122156 139466
rect 122104 139402 122156 139408
rect 188356 139398 188384 304982
rect 188436 253972 188488 253978
rect 188436 253914 188488 253920
rect 188344 139392 188396 139398
rect 188344 139334 188396 139340
rect 188448 139330 188476 253914
rect 188436 139324 188488 139330
rect 188436 139266 188488 139272
rect 189092 114510 189120 700402
rect 189356 700392 189408 700398
rect 189356 700334 189408 700340
rect 199384 700392 199436 700398
rect 199384 700334 199436 700340
rect 189172 700324 189224 700330
rect 189172 700266 189224 700272
rect 189184 117298 189212 700266
rect 189264 670812 189316 670818
rect 189264 670754 189316 670760
rect 189276 118658 189304 670754
rect 189264 118652 189316 118658
rect 189264 118594 189316 118600
rect 189172 117292 189224 117298
rect 189172 117234 189224 117240
rect 189080 114504 189132 114510
rect 189080 114446 189132 114452
rect 120998 97200 121054 97209
rect 120998 97135 121054 97144
rect 179602 80744 179658 80753
rect 179602 80679 179658 80688
rect 179788 80708 179840 80714
rect 179512 80640 179564 80646
rect 179512 80582 179564 80588
rect 127808 80436 127860 80442
rect 127808 80378 127860 80384
rect 127820 79558 127848 80378
rect 129372 80300 129424 80306
rect 129372 80242 129424 80248
rect 129280 80164 129332 80170
rect 129280 80106 129332 80112
rect 127808 79552 127860 79558
rect 127808 79494 127860 79500
rect 126244 78736 126296 78742
rect 126244 78678 126296 78684
rect 119434 78568 119490 78577
rect 119434 78503 119490 78512
rect 120724 74248 120776 74254
rect 120724 74190 120776 74196
rect 118516 46912 118568 46918
rect 118516 46854 118568 46860
rect 118332 22772 118384 22778
rect 118332 22714 118384 22720
rect 117320 18896 117372 18902
rect 117320 18838 117372 18844
rect 88352 16546 89208 16574
rect 91112 16546 91600 16574
rect 95252 16546 95832 16574
rect 96632 16546 97488 16574
rect 98012 16546 98224 16574
rect 104912 16546 105768 16574
rect 107672 16546 108160 16574
rect 111812 16546 112392 16574
rect 114572 16546 114784 16574
rect 115952 16546 116440 16574
rect 85672 10532 85724 10538
rect 85672 10474 85724 10480
rect 85684 480 85712 10474
rect 87972 6656 88024 6662
rect 87972 6598 88024 6604
rect 86868 3936 86920 3942
rect 86868 3878 86920 3884
rect 86880 480 86908 3878
rect 87984 480 88012 6598
rect 89180 480 89208 16546
rect 90364 4004 90416 4010
rect 90364 3946 90416 3952
rect 90376 480 90404 3946
rect 91572 480 91600 16546
rect 92480 10600 92532 10606
rect 92480 10542 92532 10548
rect 84446 354 84558 480
rect 84212 326 84558 354
rect 84446 -960 84558 326
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92492 354 92520 10542
rect 95148 7744 95200 7750
rect 95148 7686 95200 7692
rect 92572 6724 92624 6730
rect 92572 6666 92624 6672
rect 92584 3738 92612 6666
rect 92572 3732 92624 3738
rect 92572 3674 92624 3680
rect 93952 3732 94004 3738
rect 93952 3674 94004 3680
rect 93964 480 93992 3674
rect 95160 480 95188 7686
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 95804 354 95832 16546
rect 97460 480 97488 16546
rect 96222 354 96334 480
rect 95804 326 96334 354
rect 96222 -960 96334 326
rect 97418 -960 97530 480
rect 98196 354 98224 16546
rect 102140 11756 102192 11762
rect 102140 11698 102192 11704
rect 99840 10736 99892 10742
rect 99840 10678 99892 10684
rect 99852 480 99880 10678
rect 101034 4992 101090 5001
rect 101034 4927 101090 4936
rect 101048 480 101076 4927
rect 102152 3466 102180 11698
rect 102232 7812 102284 7818
rect 102232 7754 102284 7760
rect 102140 3460 102192 3466
rect 102140 3402 102192 3408
rect 102244 480 102272 7754
rect 104532 5228 104584 5234
rect 104532 5170 104584 5176
rect 103336 3460 103388 3466
rect 103336 3402 103388 3408
rect 103348 480 103376 3402
rect 104544 480 104572 5170
rect 105740 480 105768 16546
rect 106464 10668 106516 10674
rect 106464 10610 106516 10616
rect 98614 354 98726 480
rect 98196 326 98726 354
rect 98614 -960 98726 326
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106476 354 106504 10610
rect 108132 480 108160 16546
rect 110512 8016 110564 8022
rect 110512 7958 110564 7964
rect 109316 7880 109368 7886
rect 109316 7822 109368 7828
rect 109328 480 109356 7822
rect 110524 480 110552 7958
rect 111616 7948 111668 7954
rect 111616 7890 111668 7896
rect 111628 480 111656 7890
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112364 354 112392 16546
rect 114006 10296 114062 10305
rect 114006 10231 114062 10240
rect 114020 480 114048 10231
rect 112782 354 112894 480
rect 112364 326 112894 354
rect 112782 -960 112894 326
rect 113978 -960 114090 480
rect 114756 354 114784 16546
rect 116412 480 116440 16546
rect 115174 354 115286 480
rect 114756 326 115286 354
rect 115174 -960 115286 326
rect 116370 -960 116482 480
rect 117332 354 117360 18838
rect 120080 18828 120132 18834
rect 120080 18770 120132 18776
rect 120092 16574 120120 18770
rect 120092 16546 120672 16574
rect 119894 7712 119950 7721
rect 119894 7647 119950 7656
rect 118790 3360 118846 3369
rect 118790 3295 118846 3304
rect 118804 480 118832 3295
rect 119908 480 119936 7647
rect 117566 354 117678 480
rect 117332 326 117678 354
rect 117566 -960 117678 326
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 120644 354 120672 16546
rect 120736 3670 120764 74190
rect 124220 51128 124272 51134
rect 124220 51070 124272 51076
rect 124232 16574 124260 51070
rect 124232 16546 124720 16574
rect 123484 8084 123536 8090
rect 123484 8026 123536 8032
rect 120724 3664 120776 3670
rect 120724 3606 120776 3612
rect 122288 3392 122340 3398
rect 122288 3334 122340 3340
rect 122300 480 122328 3334
rect 123496 480 123524 8026
rect 124692 480 124720 16546
rect 126256 5098 126284 78678
rect 126336 78668 126388 78674
rect 126336 78610 126388 78616
rect 126348 18698 126376 78610
rect 127624 78600 127676 78606
rect 127624 78542 127676 78548
rect 126980 76900 127032 76906
rect 126980 76842 127032 76848
rect 126336 18692 126388 18698
rect 126336 18634 126388 18640
rect 126992 11762 127020 76842
rect 127072 75540 127124 75546
rect 127072 75482 127124 75488
rect 126980 11756 127032 11762
rect 126980 11698 127032 11704
rect 127084 6914 127112 75482
rect 127636 51134 127664 78542
rect 129096 78464 129148 78470
rect 129096 78406 129148 78412
rect 129002 77208 129058 77217
rect 129002 77143 129058 77152
rect 128360 75608 128412 75614
rect 128360 75550 128412 75556
rect 127624 51128 127676 51134
rect 127624 51070 127676 51076
rect 128372 16574 128400 75550
rect 128372 16546 128952 16574
rect 128176 11756 128228 11762
rect 128176 11698 128228 11704
rect 126992 6886 127112 6914
rect 126888 5432 126940 5438
rect 126888 5374 126940 5380
rect 126244 5092 126296 5098
rect 126244 5034 126296 5040
rect 125876 4072 125928 4078
rect 125876 4014 125928 4020
rect 125888 480 125916 4014
rect 126900 3534 126928 5374
rect 126888 3528 126940 3534
rect 126888 3470 126940 3476
rect 126992 480 127020 6886
rect 128188 480 128216 11698
rect 121062 354 121174 480
rect 120644 326 121174 354
rect 121062 -960 121174 326
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 128924 354 128952 16546
rect 129016 3602 129044 77143
rect 129108 8022 129136 78406
rect 129188 77648 129240 77654
rect 129188 77590 129240 77596
rect 129200 18902 129228 77590
rect 129292 39370 129320 80106
rect 129384 57254 129412 80242
rect 130304 80158 130640 80186
rect 130016 78396 130068 78402
rect 130016 78338 130068 78344
rect 129648 78328 129700 78334
rect 129648 78270 129700 78276
rect 129554 77752 129610 77761
rect 129554 77687 129610 77696
rect 129372 57248 129424 57254
rect 129372 57190 129424 57196
rect 129280 39364 129332 39370
rect 129280 39306 129332 39312
rect 129188 18896 129240 18902
rect 129188 18838 129240 18844
rect 129568 14618 129596 77687
rect 129556 14612 129608 14618
rect 129556 14554 129608 14560
rect 129096 8016 129148 8022
rect 129096 7958 129148 7964
rect 129660 6798 129688 78270
rect 130028 69698 130056 78338
rect 130200 77376 130252 77382
rect 130200 77318 130252 77324
rect 130108 75676 130160 75682
rect 130108 75618 130160 75624
rect 130016 69692 130068 69698
rect 130016 69634 130068 69640
rect 130120 16574 130148 75618
rect 130212 72298 130240 77318
rect 130304 72486 130332 80158
rect 130476 80028 130528 80034
rect 130476 79970 130528 79976
rect 130488 79082 130516 79970
rect 130718 79966 130746 80036
rect 130810 79966 130838 80036
rect 130706 79960 130758 79966
rect 130706 79902 130758 79908
rect 130798 79960 130850 79966
rect 130798 79902 130850 79908
rect 130660 79824 130712 79830
rect 130660 79766 130712 79772
rect 130752 79824 130804 79830
rect 130752 79766 130804 79772
rect 130568 79756 130620 79762
rect 130568 79698 130620 79704
rect 130476 79076 130528 79082
rect 130476 79018 130528 79024
rect 130580 78985 130608 79698
rect 130566 78976 130622 78985
rect 130566 78911 130622 78920
rect 130568 77716 130620 77722
rect 130568 77658 130620 77664
rect 130476 77444 130528 77450
rect 130476 77386 130528 77392
rect 130488 73930 130516 77386
rect 130580 74066 130608 77658
rect 130672 75206 130700 79766
rect 130660 75200 130712 75206
rect 130660 75142 130712 75148
rect 130580 74038 130700 74066
rect 130488 73902 130608 73930
rect 130292 72480 130344 72486
rect 130292 72422 130344 72428
rect 130212 72270 130516 72298
rect 130384 72208 130436 72214
rect 130384 72150 130436 72156
rect 130120 16546 130332 16574
rect 129648 6792 129700 6798
rect 129648 6734 129700 6740
rect 129004 3596 129056 3602
rect 129004 3538 129056 3544
rect 130304 3482 130332 16546
rect 130396 3874 130424 72150
rect 130488 10538 130516 72270
rect 130580 10606 130608 73902
rect 130672 10742 130700 74038
rect 130764 73846 130792 79766
rect 130902 79744 130930 80036
rect 130856 79716 130930 79744
rect 130856 77994 130884 79716
rect 130994 79676 131022 80036
rect 130948 79648 131022 79676
rect 131086 79676 131114 80036
rect 131178 79744 131206 80036
rect 131270 79971 131298 80036
rect 131256 79962 131312 79971
rect 131362 79966 131390 80036
rect 131256 79897 131312 79906
rect 131350 79960 131402 79966
rect 131350 79902 131402 79908
rect 131454 79898 131482 80036
rect 131442 79892 131494 79898
rect 131442 79834 131494 79840
rect 131394 79792 131450 79801
rect 131178 79716 131252 79744
rect 131546 79778 131574 80036
rect 131450 79750 131574 79778
rect 131394 79727 131450 79736
rect 131086 79648 131160 79676
rect 130948 78130 130976 79648
rect 131132 78402 131160 79648
rect 131120 78396 131172 78402
rect 131120 78338 131172 78344
rect 130936 78124 130988 78130
rect 130936 78066 130988 78072
rect 131120 78124 131172 78130
rect 131120 78066 131172 78072
rect 130844 77988 130896 77994
rect 130844 77930 130896 77936
rect 130936 77988 130988 77994
rect 130936 77930 130988 77936
rect 130752 73840 130804 73846
rect 130752 73782 130804 73788
rect 130948 70394 130976 77930
rect 131028 75744 131080 75750
rect 131028 75686 131080 75692
rect 131040 75478 131068 75686
rect 131028 75472 131080 75478
rect 131028 75414 131080 75420
rect 131132 75274 131160 78066
rect 131224 78033 131252 79716
rect 131304 79688 131356 79694
rect 131638 79676 131666 80036
rect 131730 79971 131758 80036
rect 131716 79962 131772 79971
rect 131822 79966 131850 80036
rect 131716 79897 131772 79906
rect 131810 79960 131862 79966
rect 131914 79937 131942 80036
rect 131810 79902 131862 79908
rect 131900 79928 131956 79937
rect 131900 79863 131956 79872
rect 131764 79756 131816 79762
rect 131764 79698 131816 79704
rect 131304 79630 131356 79636
rect 131394 79656 131450 79665
rect 131210 78024 131266 78033
rect 131210 77959 131266 77968
rect 131316 77897 131344 79630
rect 131394 79591 131450 79600
rect 131592 79648 131666 79676
rect 131302 77888 131358 77897
rect 131302 77823 131358 77832
rect 131212 77784 131264 77790
rect 131212 77726 131264 77732
rect 131120 75268 131172 75274
rect 131120 75210 131172 75216
rect 130764 70366 130976 70394
rect 130764 11830 130792 70366
rect 130752 11824 130804 11830
rect 130752 11766 130804 11772
rect 130660 10736 130712 10742
rect 130660 10678 130712 10684
rect 130568 10600 130620 10606
rect 130568 10542 130620 10548
rect 130476 10532 130528 10538
rect 130476 10474 130528 10480
rect 131224 4826 131252 77726
rect 131408 77294 131436 79591
rect 131592 77790 131620 79648
rect 131672 79484 131724 79490
rect 131672 79426 131724 79432
rect 131684 78946 131712 79426
rect 131672 78940 131724 78946
rect 131672 78882 131724 78888
rect 131776 78656 131804 79698
rect 132006 79676 132034 80036
rect 132098 79966 132126 80036
rect 132190 79966 132218 80036
rect 132282 79966 132310 80036
rect 132374 79966 132402 80036
rect 132086 79960 132138 79966
rect 132086 79902 132138 79908
rect 132178 79960 132230 79966
rect 132178 79902 132230 79908
rect 132270 79960 132322 79966
rect 132270 79902 132322 79908
rect 132362 79960 132414 79966
rect 132362 79902 132414 79908
rect 132466 79778 132494 80036
rect 132558 79801 132586 80036
rect 132650 79966 132678 80036
rect 132638 79960 132690 79966
rect 132742 79937 132770 80036
rect 132638 79902 132690 79908
rect 132728 79928 132784 79937
rect 132728 79863 132784 79872
rect 132132 79756 132184 79762
rect 132132 79698 132184 79704
rect 132224 79756 132276 79762
rect 132224 79698 132276 79704
rect 132420 79750 132494 79778
rect 132544 79792 132600 79801
rect 131854 79656 131910 79665
rect 131854 79591 131910 79600
rect 131960 79648 132034 79676
rect 131684 78628 131804 78656
rect 131580 77784 131632 77790
rect 131580 77726 131632 77732
rect 131408 77266 131620 77294
rect 131592 77194 131620 77266
rect 131316 77166 131620 77194
rect 131316 4894 131344 77166
rect 131396 75336 131448 75342
rect 131396 75278 131448 75284
rect 131408 4962 131436 75278
rect 131580 75268 131632 75274
rect 131580 75210 131632 75216
rect 131488 75200 131540 75206
rect 131488 75142 131540 75148
rect 131500 6186 131528 75142
rect 131592 6254 131620 75210
rect 131684 18630 131712 78628
rect 131764 77308 131816 77314
rect 131764 77250 131816 77256
rect 131672 18624 131724 18630
rect 131672 18566 131724 18572
rect 131776 10402 131804 77250
rect 131868 73914 131896 79591
rect 131856 73908 131908 73914
rect 131856 73850 131908 73856
rect 131764 10396 131816 10402
rect 131764 10338 131816 10344
rect 131580 6248 131632 6254
rect 131580 6190 131632 6196
rect 131488 6180 131540 6186
rect 131488 6122 131540 6128
rect 131396 4956 131448 4962
rect 131396 4898 131448 4904
rect 131304 4888 131356 4894
rect 131304 4830 131356 4836
rect 131212 4820 131264 4826
rect 131212 4762 131264 4768
rect 131960 4146 131988 79648
rect 132144 78062 132172 79698
rect 132132 78056 132184 78062
rect 132132 77998 132184 78004
rect 132236 75342 132264 79698
rect 132316 79688 132368 79694
rect 132316 79630 132368 79636
rect 132224 75336 132276 75342
rect 132224 75278 132276 75284
rect 132328 75206 132356 79630
rect 132420 75274 132448 79750
rect 132834 79778 132862 80036
rect 132544 79727 132600 79736
rect 132696 79750 132862 79778
rect 132500 79688 132552 79694
rect 132500 79630 132552 79636
rect 132512 78713 132540 79630
rect 132696 78742 132724 79750
rect 132926 79744 132954 80036
rect 133018 79898 133046 80036
rect 133110 79937 133138 80036
rect 133096 79928 133152 79937
rect 133006 79892 133058 79898
rect 133096 79863 133152 79872
rect 133006 79834 133058 79840
rect 133202 79812 133230 80036
rect 133294 79903 133322 80036
rect 133386 79966 133414 80036
rect 133374 79960 133426 79966
rect 133478 79937 133506 80036
rect 133280 79894 133336 79903
rect 133374 79902 133426 79908
rect 133464 79928 133520 79937
rect 133570 79898 133598 80036
rect 133464 79863 133520 79872
rect 133558 79892 133610 79898
rect 133280 79829 133336 79838
rect 133558 79834 133610 79840
rect 133156 79784 133230 79812
rect 133418 79792 133474 79801
rect 132926 79716 133000 79744
rect 132776 79688 132828 79694
rect 132972 79676 133000 79716
rect 132828 79648 132908 79676
rect 132972 79648 133046 79676
rect 132776 79630 132828 79636
rect 132774 79520 132830 79529
rect 132774 79455 132830 79464
rect 132684 78736 132736 78742
rect 132498 78704 132554 78713
rect 132684 78678 132736 78684
rect 132498 78639 132554 78648
rect 132592 77036 132644 77042
rect 132592 76978 132644 76984
rect 132408 75268 132460 75274
rect 132408 75210 132460 75216
rect 132316 75200 132368 75206
rect 132316 75142 132368 75148
rect 132604 73982 132632 76978
rect 132684 75336 132736 75342
rect 132684 75278 132736 75284
rect 132592 73976 132644 73982
rect 132592 73918 132644 73924
rect 132696 6322 132724 75278
rect 132788 6730 132816 79455
rect 132880 7614 132908 79648
rect 133018 79506 133046 79648
rect 132972 79478 133046 79506
rect 132972 77042 133000 79478
rect 133050 78432 133106 78441
rect 133050 78367 133106 78376
rect 132960 77036 133012 77042
rect 132960 76978 133012 76984
rect 133064 76566 133092 78367
rect 133052 76560 133104 76566
rect 133052 76502 133104 76508
rect 133052 75268 133104 75274
rect 133052 75210 133104 75216
rect 132960 75200 133012 75206
rect 132960 75142 133012 75148
rect 132972 8974 133000 75142
rect 133064 44878 133092 75210
rect 133052 44872 133104 44878
rect 133052 44814 133104 44820
rect 132960 8968 133012 8974
rect 132960 8910 133012 8916
rect 132868 7608 132920 7614
rect 132868 7550 132920 7556
rect 132776 6724 132828 6730
rect 132776 6666 132828 6672
rect 132684 6316 132736 6322
rect 132684 6258 132736 6264
rect 133156 5030 133184 79784
rect 133662 79744 133690 80036
rect 133418 79727 133474 79736
rect 133236 79688 133288 79694
rect 133236 79630 133288 79636
rect 133248 78674 133276 79630
rect 133236 78668 133288 78674
rect 133236 78610 133288 78616
rect 133328 78668 133380 78674
rect 133328 78610 133380 78616
rect 133340 75206 133368 78610
rect 133328 75200 133380 75206
rect 133328 75142 133380 75148
rect 133432 70394 133460 79727
rect 133616 79716 133690 79744
rect 133512 79688 133564 79694
rect 133512 79630 133564 79636
rect 133524 76634 133552 79630
rect 133512 76628 133564 76634
rect 133512 76570 133564 76576
rect 133616 75274 133644 79716
rect 133754 79506 133782 80036
rect 133846 79966 133874 80036
rect 133938 79966 133966 80036
rect 134030 79971 134058 80036
rect 133834 79960 133886 79966
rect 133834 79902 133886 79908
rect 133926 79960 133978 79966
rect 133926 79902 133978 79908
rect 134016 79962 134072 79971
rect 134016 79897 134072 79906
rect 134122 79835 134150 80036
rect 133972 79824 134024 79830
rect 133972 79766 134024 79772
rect 134108 79826 134164 79835
rect 133754 79478 133828 79506
rect 133800 75342 133828 79478
rect 133880 79008 133932 79014
rect 133880 78950 133932 78956
rect 133892 78810 133920 78950
rect 133880 78804 133932 78810
rect 133880 78746 133932 78752
rect 133984 78674 134012 79766
rect 134108 79761 134164 79770
rect 134214 79676 134242 80036
rect 134306 79937 134334 80036
rect 134292 79928 134348 79937
rect 134292 79863 134348 79872
rect 134168 79648 134242 79676
rect 134064 79416 134116 79422
rect 134064 79358 134116 79364
rect 133880 78668 134012 78674
rect 133932 78646 134012 78668
rect 133880 78610 133932 78616
rect 134076 78520 134104 79358
rect 133892 78492 134104 78520
rect 133788 75336 133840 75342
rect 133788 75278 133840 75284
rect 133892 75274 133920 78492
rect 134064 78396 134116 78402
rect 134064 78338 134116 78344
rect 133970 78160 134026 78169
rect 133970 78095 133972 78104
rect 134024 78095 134026 78104
rect 133972 78066 134024 78072
rect 133604 75268 133656 75274
rect 133604 75210 133656 75216
rect 133880 75268 133932 75274
rect 133880 75210 133932 75216
rect 133880 73296 133932 73302
rect 133880 73238 133932 73244
rect 133340 70366 133460 70394
rect 133340 5438 133368 70366
rect 133328 5432 133380 5438
rect 133328 5374 133380 5380
rect 133144 5024 133196 5030
rect 133144 4966 133196 4972
rect 131948 4140 132000 4146
rect 131948 4082 132000 4088
rect 130384 3868 130436 3874
rect 130384 3810 130436 3816
rect 130304 3454 130608 3482
rect 130580 480 130608 3454
rect 131764 3460 131816 3466
rect 131764 3402 131816 3408
rect 131776 480 131804 3402
rect 132960 3120 133012 3126
rect 132960 3062 133012 3068
rect 132972 480 133000 3062
rect 129342 354 129454 480
rect 128924 326 129454 354
rect 129342 -960 129454 326
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 133892 354 133920 73238
rect 134076 6458 134104 78338
rect 134168 77217 134196 79648
rect 134398 79540 134426 80036
rect 134490 79898 134518 80036
rect 134478 79892 134530 79898
rect 134478 79834 134530 79840
rect 134582 79830 134610 80036
rect 134674 79830 134702 80036
rect 134570 79824 134622 79830
rect 134570 79766 134622 79772
rect 134662 79824 134714 79830
rect 134766 79812 134794 80036
rect 134858 79971 134886 80036
rect 134844 79962 134900 79971
rect 134844 79897 134900 79906
rect 134950 79898 134978 80036
rect 134938 79892 134990 79898
rect 134938 79834 134990 79840
rect 134766 79801 134840 79812
rect 134766 79792 134854 79801
rect 134766 79784 134798 79792
rect 134662 79766 134714 79772
rect 135042 79778 135070 80036
rect 135134 79966 135162 80036
rect 135226 79966 135254 80036
rect 135122 79960 135174 79966
rect 135122 79902 135174 79908
rect 135214 79960 135266 79966
rect 135214 79902 135266 79908
rect 134798 79727 134854 79736
rect 134996 79750 135070 79778
rect 135166 79792 135222 79801
rect 134890 79656 134946 79665
rect 134890 79591 134946 79600
rect 134524 79552 134576 79558
rect 134398 79512 134472 79540
rect 134248 79280 134300 79286
rect 134248 79222 134300 79228
rect 134260 79082 134288 79222
rect 134248 79076 134300 79082
rect 134248 79018 134300 79024
rect 134444 78033 134472 79512
rect 134524 79494 134576 79500
rect 134798 79520 134854 79529
rect 134430 78024 134486 78033
rect 134430 77959 134486 77968
rect 134536 77976 134564 79494
rect 134708 79484 134760 79490
rect 134798 79455 134854 79464
rect 134708 79426 134760 79432
rect 134616 79416 134668 79422
rect 134616 79358 134668 79364
rect 134628 78402 134656 79358
rect 134616 78396 134668 78402
rect 134616 78338 134668 78344
rect 134536 77948 134656 77976
rect 134524 77580 134576 77586
rect 134524 77522 134576 77528
rect 134154 77208 134210 77217
rect 134154 77143 134210 77152
rect 134156 75268 134208 75274
rect 134156 75210 134208 75216
rect 134248 75268 134300 75274
rect 134248 75210 134300 75216
rect 134168 9042 134196 75210
rect 134260 9110 134288 75210
rect 134340 75200 134392 75206
rect 134340 75142 134392 75148
rect 134352 9178 134380 75142
rect 134536 10470 134564 77522
rect 134628 75410 134656 77948
rect 134616 75404 134668 75410
rect 134616 75346 134668 75352
rect 134524 10464 134576 10470
rect 134524 10406 134576 10412
rect 134340 9172 134392 9178
rect 134340 9114 134392 9120
rect 134248 9104 134300 9110
rect 134248 9046 134300 9052
rect 134156 9036 134208 9042
rect 134156 8978 134208 8984
rect 134064 6452 134116 6458
rect 134064 6394 134116 6400
rect 134720 6390 134748 79426
rect 134812 75274 134840 79455
rect 134800 75268 134852 75274
rect 134800 75210 134852 75216
rect 134904 71058 134932 79591
rect 134996 75206 135024 79750
rect 135318 79778 135346 80036
rect 135410 79966 135438 80036
rect 135502 79971 135530 80036
rect 135398 79960 135450 79966
rect 135398 79902 135450 79908
rect 135488 79962 135544 79971
rect 135594 79966 135622 80036
rect 135686 79971 135714 80036
rect 135488 79897 135544 79906
rect 135582 79960 135634 79966
rect 135582 79902 135634 79908
rect 135672 79962 135728 79971
rect 135672 79897 135728 79906
rect 135778 79898 135806 80036
rect 135870 79898 135898 80036
rect 135962 79898 135990 80036
rect 136054 79898 136082 80036
rect 135766 79892 135818 79898
rect 135766 79834 135818 79840
rect 135858 79892 135910 79898
rect 135858 79834 135910 79840
rect 135950 79892 136002 79898
rect 135950 79834 136002 79840
rect 136042 79892 136094 79898
rect 136042 79834 136094 79840
rect 136146 79835 136174 80036
rect 136238 79966 136266 80036
rect 136226 79960 136278 79966
rect 136226 79902 136278 79908
rect 136132 79826 136188 79835
rect 136330 79830 136358 80036
rect 136422 79971 136450 80036
rect 136408 79962 136464 79971
rect 136514 79966 136542 80036
rect 136408 79897 136464 79906
rect 136502 79960 136554 79966
rect 136502 79902 136554 79908
rect 135222 79750 135346 79778
rect 135902 79792 135958 79801
rect 135720 79756 135772 79762
rect 135166 79727 135222 79736
rect 135720 79698 135772 79704
rect 135812 79756 135864 79762
rect 136132 79761 136188 79770
rect 136318 79824 136370 79830
rect 136318 79766 136370 79772
rect 136456 79824 136508 79830
rect 136456 79766 136508 79772
rect 135902 79727 135958 79736
rect 135812 79698 135864 79704
rect 135076 79688 135128 79694
rect 135076 79630 135128 79636
rect 135352 79688 135404 79694
rect 135352 79630 135404 79636
rect 134984 75200 135036 75206
rect 134984 75142 135036 75148
rect 135088 72554 135116 79630
rect 135168 79620 135220 79626
rect 135168 79562 135220 79568
rect 135180 74254 135208 79562
rect 135260 79076 135312 79082
rect 135260 79018 135312 79024
rect 135272 76702 135300 79018
rect 135260 76696 135312 76702
rect 135260 76638 135312 76644
rect 135364 75449 135392 79630
rect 135628 79620 135680 79626
rect 135628 79562 135680 79568
rect 135442 79520 135498 79529
rect 135442 79455 135498 79464
rect 135536 79484 135588 79490
rect 135456 78033 135484 79455
rect 135536 79426 135588 79432
rect 135442 78024 135498 78033
rect 135442 77959 135498 77968
rect 135548 75914 135576 79426
rect 135640 78033 135668 79562
rect 135626 78024 135682 78033
rect 135626 77959 135682 77968
rect 135456 75886 135576 75914
rect 135350 75440 135406 75449
rect 135350 75375 135406 75384
rect 135168 74248 135220 74254
rect 135168 74190 135220 74196
rect 135076 72548 135128 72554
rect 135076 72490 135128 72496
rect 134892 71052 134944 71058
rect 134892 70994 134944 71000
rect 135456 6526 135484 75886
rect 135536 75200 135588 75206
rect 135536 75142 135588 75148
rect 135548 6594 135576 75142
rect 135628 71800 135680 71806
rect 135628 71742 135680 71748
rect 135536 6588 135588 6594
rect 135536 6530 135588 6536
rect 135444 6520 135496 6526
rect 135444 6462 135496 6468
rect 134708 6384 134760 6390
rect 134708 6326 134760 6332
rect 135640 1986 135668 71742
rect 135732 7682 135760 79698
rect 135824 77314 135852 79698
rect 135812 77308 135864 77314
rect 135812 77250 135864 77256
rect 135916 64874 135944 79727
rect 136178 79656 136234 79665
rect 136088 79620 136140 79626
rect 136178 79591 136234 79600
rect 136088 79562 136140 79568
rect 135996 79552 136048 79558
rect 135996 79494 136048 79500
rect 136008 75478 136036 79494
rect 135996 75472 136048 75478
rect 135996 75414 136048 75420
rect 135996 75268 136048 75274
rect 135996 75210 136048 75216
rect 135824 64846 135944 64874
rect 135824 10334 135852 64846
rect 135812 10328 135864 10334
rect 135812 10270 135864 10276
rect 135720 7676 135772 7682
rect 135720 7618 135772 7624
rect 136008 3806 136036 75210
rect 136100 5166 136128 79562
rect 136192 74050 136220 79591
rect 136362 79520 136418 79529
rect 136272 79484 136324 79490
rect 136362 79455 136418 79464
rect 136272 79426 136324 79432
rect 136180 74044 136232 74050
rect 136180 73986 136232 73992
rect 136284 72214 136312 79426
rect 136376 77586 136404 79455
rect 136364 77580 136416 77586
rect 136364 77522 136416 77528
rect 136468 75274 136496 79766
rect 136606 79676 136634 80036
rect 136698 79971 136726 80036
rect 136684 79962 136740 79971
rect 136684 79897 136740 79906
rect 136790 79676 136818 80036
rect 136882 79966 136910 80036
rect 136870 79960 136922 79966
rect 136870 79902 136922 79908
rect 136974 79676 137002 80036
rect 137066 79966 137094 80036
rect 137054 79960 137106 79966
rect 137054 79902 137106 79908
rect 137158 79812 137186 80036
rect 137250 79966 137278 80036
rect 137238 79960 137290 79966
rect 137238 79902 137290 79908
rect 136560 79648 136634 79676
rect 136744 79648 136818 79676
rect 136928 79648 137002 79676
rect 137112 79784 137186 79812
rect 136456 75268 136508 75274
rect 136456 75210 136508 75216
rect 136560 75206 136588 79648
rect 136640 79552 136692 79558
rect 136640 79494 136692 79500
rect 136652 76673 136680 79494
rect 136744 78198 136772 79648
rect 136928 79422 136956 79648
rect 137008 79552 137060 79558
rect 137008 79494 137060 79500
rect 136916 79416 136968 79422
rect 136916 79358 136968 79364
rect 137020 78674 137048 79494
rect 137112 79082 137140 79784
rect 137342 79744 137370 80036
rect 137434 79898 137462 80036
rect 137526 79966 137554 80036
rect 137514 79960 137566 79966
rect 137514 79902 137566 79908
rect 137422 79892 137474 79898
rect 137422 79834 137474 79840
rect 137618 79812 137646 80036
rect 137710 79937 137738 80036
rect 137696 79928 137752 79937
rect 137696 79863 137752 79872
rect 137618 79784 137692 79812
rect 137296 79716 137370 79744
rect 137192 79688 137244 79694
rect 137192 79630 137244 79636
rect 137100 79076 137152 79082
rect 137100 79018 137152 79024
rect 136928 78646 137048 78674
rect 137100 78668 137152 78674
rect 136822 78432 136878 78441
rect 136822 78367 136878 78376
rect 136732 78192 136784 78198
rect 136732 78134 136784 78140
rect 136638 76664 136694 76673
rect 136638 76599 136694 76608
rect 136548 75200 136600 75206
rect 136548 75142 136600 75148
rect 136272 72208 136324 72214
rect 136272 72150 136324 72156
rect 136088 5160 136140 5166
rect 136088 5102 136140 5108
rect 135996 3800 136048 3806
rect 135996 3742 136048 3748
rect 136836 3738 136864 78367
rect 136928 74118 136956 78646
rect 137100 78610 137152 78616
rect 137008 78056 137060 78062
rect 137008 77998 137060 78004
rect 136916 74112 136968 74118
rect 136916 74054 136968 74060
rect 136916 73228 136968 73234
rect 136916 73170 136968 73176
rect 136824 3732 136876 3738
rect 136824 3674 136876 3680
rect 136456 3596 136508 3602
rect 136456 3538 136508 3544
rect 135272 1958 135668 1986
rect 135272 480 135300 1958
rect 136468 480 136496 3538
rect 136928 490 136956 73170
rect 137020 6662 137048 77998
rect 137112 7750 137140 78610
rect 137204 22846 137232 79630
rect 137192 22840 137244 22846
rect 137192 22782 137244 22788
rect 137100 7744 137152 7750
rect 137100 7686 137152 7692
rect 137008 6656 137060 6662
rect 137008 6598 137060 6604
rect 137296 3942 137324 79716
rect 137664 79608 137692 79784
rect 137802 79676 137830 80036
rect 137894 79937 137922 80036
rect 137986 79966 138014 80036
rect 138078 79966 138106 80036
rect 138170 79966 138198 80036
rect 137974 79960 138026 79966
rect 137880 79928 137936 79937
rect 137974 79902 138026 79908
rect 138066 79960 138118 79966
rect 138066 79902 138118 79908
rect 138158 79960 138210 79966
rect 138158 79902 138210 79908
rect 137880 79863 137936 79872
rect 138262 79812 138290 80036
rect 138216 79801 138290 79812
rect 138202 79792 138290 79801
rect 138258 79784 138290 79792
rect 138202 79727 138258 79736
rect 137928 79688 137980 79694
rect 137802 79648 137876 79676
rect 137572 79580 137692 79608
rect 137376 79552 137428 79558
rect 137376 79494 137428 79500
rect 137388 78062 137416 79494
rect 137468 79416 137520 79422
rect 137468 79358 137520 79364
rect 137376 78056 137428 78062
rect 137376 77998 137428 78004
rect 137480 75750 137508 79358
rect 137468 75744 137520 75750
rect 137468 75686 137520 75692
rect 137572 64874 137600 79580
rect 137742 79520 137798 79529
rect 137652 79484 137704 79490
rect 137742 79455 137798 79464
rect 137652 79426 137704 79432
rect 137664 77382 137692 79426
rect 137652 77376 137704 77382
rect 137652 77318 137704 77324
rect 137756 76838 137784 79455
rect 137848 77450 137876 79648
rect 137928 79630 137980 79636
rect 138112 79688 138164 79694
rect 138112 79630 138164 79636
rect 137940 78713 137968 79630
rect 138020 79620 138072 79626
rect 138020 79562 138072 79568
rect 137926 78704 137982 78713
rect 138032 78674 138060 79562
rect 137926 78639 137982 78648
rect 138020 78668 138072 78674
rect 138020 78610 138072 78616
rect 138124 78266 138152 79630
rect 138354 79540 138382 80036
rect 138446 79966 138474 80036
rect 138538 79966 138566 80036
rect 138630 79971 138658 80036
rect 138434 79960 138486 79966
rect 138434 79902 138486 79908
rect 138526 79960 138578 79966
rect 138526 79902 138578 79908
rect 138616 79962 138672 79971
rect 138616 79897 138672 79906
rect 138722 79898 138750 80036
rect 138814 79971 138842 80036
rect 138800 79962 138856 79971
rect 138906 79966 138934 80036
rect 138998 79966 139026 80036
rect 139090 79971 139118 80036
rect 138710 79892 138762 79898
rect 138800 79897 138856 79906
rect 138894 79960 138946 79966
rect 138894 79902 138946 79908
rect 138986 79960 139038 79966
rect 138986 79902 139038 79908
rect 139076 79962 139132 79971
rect 139076 79897 139132 79906
rect 138710 79834 138762 79840
rect 138434 79824 138486 79830
rect 138432 79792 138434 79801
rect 139182 79812 139210 80036
rect 139274 79966 139302 80036
rect 139366 79966 139394 80036
rect 139262 79960 139314 79966
rect 139262 79902 139314 79908
rect 139354 79960 139406 79966
rect 139354 79902 139406 79908
rect 138486 79792 138488 79801
rect 138432 79727 138488 79736
rect 138570 79792 138626 79801
rect 138570 79727 138626 79736
rect 138754 79792 138810 79801
rect 138754 79727 138810 79736
rect 139136 79784 139210 79812
rect 138480 79620 138532 79626
rect 138480 79562 138532 79568
rect 138354 79512 138428 79540
rect 138204 79484 138256 79490
rect 138204 79426 138256 79432
rect 138112 78260 138164 78266
rect 138112 78202 138164 78208
rect 137836 77444 137888 77450
rect 137836 77386 137888 77392
rect 137744 76832 137796 76838
rect 137744 76774 137796 76780
rect 138020 75132 138072 75138
rect 138020 75074 138072 75080
rect 137388 64846 137600 64874
rect 137388 4010 137416 64846
rect 138032 6914 138060 75074
rect 138216 7818 138244 79426
rect 138296 79212 138348 79218
rect 138296 79154 138348 79160
rect 138308 76770 138336 79154
rect 138400 77722 138428 79512
rect 138388 77716 138440 77722
rect 138388 77658 138440 77664
rect 138296 76764 138348 76770
rect 138296 76706 138348 76712
rect 138296 75268 138348 75274
rect 138296 75210 138348 75216
rect 138308 7954 138336 75210
rect 138388 75200 138440 75206
rect 138388 75142 138440 75148
rect 138296 7948 138348 7954
rect 138296 7890 138348 7896
rect 138400 7886 138428 75142
rect 138492 10674 138520 79562
rect 138584 77994 138612 79727
rect 138664 79552 138716 79558
rect 138664 79494 138716 79500
rect 138676 79098 138704 79494
rect 138768 79218 138796 79727
rect 138940 79688 138992 79694
rect 138940 79630 138992 79636
rect 138848 79416 138900 79422
rect 138848 79358 138900 79364
rect 138756 79212 138808 79218
rect 138756 79154 138808 79160
rect 138676 79070 138796 79098
rect 138664 79008 138716 79014
rect 138664 78950 138716 78956
rect 138676 78810 138704 78950
rect 138664 78804 138716 78810
rect 138664 78746 138716 78752
rect 138572 77988 138624 77994
rect 138572 77930 138624 77936
rect 138572 75336 138624 75342
rect 138572 75278 138624 75284
rect 138584 18766 138612 75278
rect 138768 70394 138796 79070
rect 138860 78470 138888 79358
rect 138848 78464 138900 78470
rect 138848 78406 138900 78412
rect 138952 72622 138980 79630
rect 139030 79520 139086 79529
rect 139030 79455 139086 79464
rect 139044 75206 139072 79455
rect 139136 79422 139164 79784
rect 139458 79778 139486 80036
rect 139550 79898 139578 80036
rect 139538 79892 139590 79898
rect 139538 79834 139590 79840
rect 139642 79830 139670 80036
rect 139412 79750 139486 79778
rect 139630 79824 139682 79830
rect 139630 79766 139682 79772
rect 139216 79688 139268 79694
rect 139216 79630 139268 79636
rect 139308 79688 139360 79694
rect 139412 79665 139440 79750
rect 139492 79688 139544 79694
rect 139308 79630 139360 79636
rect 139398 79656 139454 79665
rect 139124 79416 139176 79422
rect 139124 79358 139176 79364
rect 139124 79212 139176 79218
rect 139124 79154 139176 79160
rect 139032 75200 139084 75206
rect 139032 75142 139084 75148
rect 139136 75138 139164 79154
rect 139228 75274 139256 79630
rect 139320 75342 139348 79630
rect 139734 79676 139762 80036
rect 139826 79812 139854 80036
rect 139918 79971 139946 80036
rect 139904 79962 139960 79971
rect 140010 79966 140038 80036
rect 140102 79966 140130 80036
rect 140194 79966 140222 80036
rect 139904 79897 139960 79906
rect 139998 79960 140050 79966
rect 139998 79902 140050 79908
rect 140090 79960 140142 79966
rect 140090 79902 140142 79908
rect 140182 79960 140234 79966
rect 140182 79902 140234 79908
rect 140286 79903 140314 80036
rect 140272 79894 140328 79903
rect 140272 79829 140328 79838
rect 140378 79830 140406 80036
rect 140470 79898 140498 80036
rect 140458 79892 140510 79898
rect 140458 79834 140510 79840
rect 140366 79824 140418 79830
rect 139826 79784 139900 79812
rect 139544 79648 139624 79676
rect 139492 79630 139544 79636
rect 139398 79591 139454 79600
rect 139492 79552 139544 79558
rect 139492 79494 139544 79500
rect 139400 77784 139452 77790
rect 139400 77726 139452 77732
rect 139308 75336 139360 75342
rect 139308 75278 139360 75284
rect 139216 75268 139268 75274
rect 139216 75210 139268 75216
rect 139124 75132 139176 75138
rect 139124 75074 139176 75080
rect 138940 72616 138992 72622
rect 138940 72558 138992 72564
rect 139412 71806 139440 77726
rect 139504 76945 139532 79494
rect 139490 76936 139546 76945
rect 139490 76871 139546 76880
rect 139596 76820 139624 79648
rect 139688 79648 139762 79676
rect 139872 79665 139900 79784
rect 140134 79792 140190 79801
rect 140562 79812 140590 80036
rect 140654 79971 140682 80036
rect 140640 79962 140696 79971
rect 140640 79897 140696 79906
rect 140746 79898 140774 80036
rect 140734 79892 140786 79898
rect 140734 79834 140786 79840
rect 140562 79784 140636 79812
rect 140838 79801 140866 80036
rect 140930 79898 140958 80036
rect 141022 79898 141050 80036
rect 140918 79892 140970 79898
rect 140918 79834 140970 79840
rect 141010 79892 141062 79898
rect 141010 79834 141062 79840
rect 141114 79830 141142 80036
rect 141102 79824 141154 79830
rect 140366 79766 140418 79772
rect 140134 79727 140190 79736
rect 140228 79756 140280 79762
rect 139952 79688 140004 79694
rect 139858 79656 139914 79665
rect 139688 77654 139716 79648
rect 140004 79648 140084 79676
rect 139952 79630 140004 79636
rect 139858 79591 139914 79600
rect 139768 79416 139820 79422
rect 139768 79358 139820 79364
rect 139952 79416 140004 79422
rect 139952 79358 140004 79364
rect 139676 77648 139728 77654
rect 139676 77590 139728 77596
rect 139504 76792 139624 76820
rect 139504 74186 139532 76792
rect 139780 76752 139808 79358
rect 139860 79076 139912 79082
rect 139860 79018 139912 79024
rect 139596 76724 139808 76752
rect 139492 74180 139544 74186
rect 139492 74122 139544 74128
rect 139400 71800 139452 71806
rect 139400 71742 139452 71748
rect 138768 70366 139072 70394
rect 138572 18760 138624 18766
rect 138572 18702 138624 18708
rect 138480 10668 138532 10674
rect 138480 10610 138532 10616
rect 138388 7880 138440 7886
rect 138388 7822 138440 7828
rect 138204 7812 138256 7818
rect 138204 7754 138256 7760
rect 138032 6886 138888 6914
rect 137376 4004 137428 4010
rect 137376 3946 137428 3952
rect 137284 3936 137336 3942
rect 137284 3878 137336 3884
rect 134126 354 134238 480
rect 133892 326 134238 354
rect 134126 -960 134238 326
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 136928 462 137232 490
rect 138860 480 138888 6886
rect 139044 5234 139072 70366
rect 139596 8090 139624 76724
rect 139768 76152 139820 76158
rect 139768 76094 139820 76100
rect 139676 75404 139728 75410
rect 139676 75346 139728 75352
rect 139688 18834 139716 75346
rect 139676 18828 139728 18834
rect 139676 18770 139728 18776
rect 139584 8084 139636 8090
rect 139584 8026 139636 8032
rect 139032 5228 139084 5234
rect 139032 5170 139084 5176
rect 139780 3398 139808 76094
rect 139872 75313 139900 79018
rect 139964 76158 139992 79358
rect 139952 76152 140004 76158
rect 139952 76094 140004 76100
rect 139952 76016 140004 76022
rect 139952 75958 140004 75964
rect 139858 75304 139914 75313
rect 139858 75239 139914 75248
rect 139964 4078 139992 75958
rect 140056 75410 140084 79648
rect 140148 79082 140176 79727
rect 140608 79744 140636 79784
rect 140228 79698 140280 79704
rect 140516 79716 140636 79744
rect 140824 79792 140880 79801
rect 141102 79766 141154 79772
rect 140824 79727 140880 79736
rect 140136 79076 140188 79082
rect 140136 79018 140188 79024
rect 140240 76022 140268 79698
rect 140412 79688 140464 79694
rect 140318 79656 140374 79665
rect 140412 79630 140464 79636
rect 140318 79591 140374 79600
rect 140332 78606 140360 79591
rect 140320 78600 140372 78606
rect 140320 78542 140372 78548
rect 140228 76016 140280 76022
rect 140228 75958 140280 75964
rect 140228 75880 140280 75886
rect 140228 75822 140280 75828
rect 140044 75404 140096 75410
rect 140044 75346 140096 75352
rect 140044 75268 140096 75274
rect 140044 75210 140096 75216
rect 139952 4072 140004 4078
rect 139952 4014 140004 4020
rect 140056 3618 140084 75210
rect 140136 75200 140188 75206
rect 140136 75142 140188 75148
rect 139964 3590 140084 3618
rect 139964 3466 139992 3590
rect 140044 3528 140096 3534
rect 140044 3470 140096 3476
rect 139952 3460 140004 3466
rect 139952 3402 140004 3408
rect 139768 3392 139820 3398
rect 139768 3334 139820 3340
rect 140056 480 140084 3470
rect 140148 3126 140176 75142
rect 140240 3602 140268 75822
rect 140424 75546 140452 79630
rect 140516 76906 140544 79716
rect 141206 79676 141234 80036
rect 141298 79830 141326 80036
rect 141390 79937 141418 80036
rect 141376 79928 141432 79937
rect 141482 79898 141510 80036
rect 141574 79937 141602 80036
rect 141560 79928 141616 79937
rect 141376 79863 141432 79872
rect 141470 79892 141522 79898
rect 141666 79898 141694 80036
rect 141758 79971 141786 80036
rect 141744 79962 141800 79971
rect 141850 79966 141878 80036
rect 141560 79863 141616 79872
rect 141654 79892 141706 79898
rect 141744 79897 141800 79906
rect 141838 79960 141890 79966
rect 141838 79902 141890 79908
rect 141942 79903 141970 80036
rect 141470 79834 141522 79840
rect 141654 79834 141706 79840
rect 141928 79894 141984 79903
rect 141286 79824 141338 79830
rect 141928 79829 141984 79838
rect 141286 79766 141338 79772
rect 141698 79792 141754 79801
rect 141378 79756 141430 79762
rect 141430 79716 141510 79744
rect 141698 79727 141754 79736
rect 141792 79756 141844 79762
rect 141378 79698 141430 79704
rect 140594 79656 140650 79665
rect 140870 79656 140926 79665
rect 140650 79614 140728 79642
rect 140594 79591 140650 79600
rect 140596 79484 140648 79490
rect 140596 79426 140648 79432
rect 140608 77790 140636 79426
rect 140596 77784 140648 77790
rect 140596 77726 140648 77732
rect 140596 77104 140648 77110
rect 140596 77046 140648 77052
rect 140504 76900 140556 76906
rect 140504 76842 140556 76848
rect 140412 75540 140464 75546
rect 140412 75482 140464 75488
rect 140608 73302 140636 77046
rect 140700 75614 140728 79614
rect 140780 79620 140832 79626
rect 141206 79648 141280 79676
rect 140870 79591 140926 79600
rect 141056 79620 141108 79626
rect 140780 79562 140832 79568
rect 140792 75682 140820 79562
rect 140780 75676 140832 75682
rect 140780 75618 140832 75624
rect 140688 75608 140740 75614
rect 140688 75550 140740 75556
rect 140884 75274 140912 79591
rect 141056 79562 141108 79568
rect 140964 79552 141016 79558
rect 140964 79494 141016 79500
rect 140872 75268 140924 75274
rect 140872 75210 140924 75216
rect 140976 75206 141004 79494
rect 141068 77110 141096 79562
rect 141148 79416 141200 79422
rect 141148 79358 141200 79364
rect 141056 77104 141108 77110
rect 141056 77046 141108 77052
rect 140964 75200 141016 75206
rect 140964 75142 141016 75148
rect 141056 75200 141108 75206
rect 141056 75142 141108 75148
rect 140962 75032 141018 75041
rect 140962 74967 141018 74976
rect 140596 73296 140648 73302
rect 140596 73238 140648 73244
rect 140976 4146 141004 74967
rect 140964 4140 141016 4146
rect 140964 4082 141016 4088
rect 141068 3874 141096 75142
rect 141056 3868 141108 3874
rect 141056 3810 141108 3816
rect 140228 3596 140280 3602
rect 140228 3538 140280 3544
rect 141160 3534 141188 79358
rect 141252 75886 141280 79648
rect 141330 79656 141386 79665
rect 141482 79642 141510 79716
rect 141330 79591 141386 79600
rect 141436 79614 141510 79642
rect 141608 79620 141660 79626
rect 141344 79218 141372 79591
rect 141332 79212 141384 79218
rect 141332 79154 141384 79160
rect 141240 75880 141292 75886
rect 141240 75822 141292 75828
rect 141240 75744 141292 75750
rect 141240 75686 141292 75692
rect 141252 3738 141280 75686
rect 141332 75268 141384 75274
rect 141332 75210 141384 75216
rect 141344 44946 141372 75210
rect 141436 73234 141464 79614
rect 141608 79562 141660 79568
rect 141514 79520 141570 79529
rect 141514 79455 141570 79464
rect 141424 73228 141476 73234
rect 141424 73170 141476 73176
rect 141528 70394 141556 79455
rect 141620 75750 141648 79562
rect 141608 75744 141660 75750
rect 141608 75686 141660 75692
rect 141712 70394 141740 79727
rect 141792 79698 141844 79704
rect 141884 79756 141936 79762
rect 141884 79698 141936 79704
rect 141804 79665 141832 79698
rect 141790 79656 141846 79665
rect 141790 79591 141846 79600
rect 141790 78976 141846 78985
rect 141790 78911 141846 78920
rect 141804 75274 141832 78911
rect 141896 75274 141924 79698
rect 142034 79676 142062 80036
rect 142126 79744 142154 80036
rect 142218 79812 142246 80036
rect 142310 79937 142338 80036
rect 142402 79966 142430 80036
rect 142390 79960 142442 79966
rect 142296 79928 142352 79937
rect 142390 79902 142442 79908
rect 142296 79863 142352 79872
rect 142494 79812 142522 80036
rect 142218 79784 142384 79812
rect 142126 79716 142200 79744
rect 141988 79648 142062 79676
rect 141792 75268 141844 75274
rect 141792 75210 141844 75216
rect 141884 75268 141936 75274
rect 141884 75210 141936 75216
rect 141988 75206 142016 79648
rect 142068 76832 142120 76838
rect 142068 76774 142120 76780
rect 141976 75200 142028 75206
rect 141976 75142 142028 75148
rect 142080 71774 142108 76774
rect 142172 75313 142200 79716
rect 142252 79688 142304 79694
rect 142252 79630 142304 79636
rect 142158 75304 142214 75313
rect 142158 75239 142214 75248
rect 142080 71746 142200 71774
rect 141436 70366 141556 70394
rect 141620 70366 141740 70394
rect 141332 44940 141384 44946
rect 141332 44882 141384 44888
rect 141240 3732 141292 3738
rect 141240 3674 141292 3680
rect 141148 3528 141200 3534
rect 141148 3470 141200 3476
rect 140136 3120 140188 3126
rect 140136 3062 140188 3068
rect 137204 354 137232 462
rect 137622 354 137734 480
rect 137204 326 137734 354
rect 137622 -960 137734 326
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 354 141322 480
rect 141436 354 141464 70366
rect 141620 3602 141648 70366
rect 142172 3806 142200 71746
rect 142264 4962 142292 79630
rect 142356 75410 142384 79784
rect 142448 79784 142522 79812
rect 142448 76770 142476 79784
rect 142586 79744 142614 80036
rect 142540 79716 142614 79744
rect 142540 76838 142568 79716
rect 142678 79676 142706 80036
rect 142770 79778 142798 80036
rect 142862 79966 142890 80036
rect 142850 79960 142902 79966
rect 142850 79902 142902 79908
rect 142954 79898 142982 80036
rect 143046 79937 143074 80036
rect 143032 79928 143088 79937
rect 142942 79892 142994 79898
rect 143032 79863 143088 79872
rect 142942 79834 142994 79840
rect 142894 79792 142950 79801
rect 142770 79750 142844 79778
rect 142632 79648 142706 79676
rect 142528 76832 142580 76838
rect 142528 76774 142580 76780
rect 142436 76764 142488 76770
rect 142436 76706 142488 76712
rect 142632 76514 142660 79648
rect 142712 76900 142764 76906
rect 142712 76842 142764 76848
rect 142448 76486 142660 76514
rect 142344 75404 142396 75410
rect 142344 75346 142396 75352
rect 142344 75268 142396 75274
rect 142344 75210 142396 75216
rect 142356 5030 142384 75210
rect 142448 6254 142476 76486
rect 142528 75948 142580 75954
rect 142528 75890 142580 75896
rect 142540 15910 142568 75890
rect 142620 75404 142672 75410
rect 142620 75346 142672 75352
rect 142632 44198 142660 75346
rect 142724 51746 142752 76842
rect 142816 75954 142844 79750
rect 143138 79778 143166 80036
rect 143230 79966 143258 80036
rect 143218 79960 143270 79966
rect 143322 79937 143350 80036
rect 143218 79902 143270 79908
rect 143308 79928 143364 79937
rect 143308 79863 143364 79872
rect 143414 79812 143442 80036
rect 143506 79971 143534 80036
rect 143492 79962 143548 79971
rect 143492 79897 143548 79906
rect 143598 79812 143626 80036
rect 143414 79784 143488 79812
rect 142894 79727 142950 79736
rect 143000 79750 143166 79778
rect 142804 75948 142856 75954
rect 142804 75890 142856 75896
rect 142908 71774 142936 79727
rect 143000 76537 143028 79750
rect 143080 79688 143132 79694
rect 143080 79630 143132 79636
rect 143172 79688 143224 79694
rect 143172 79630 143224 79636
rect 143092 76906 143120 79630
rect 143080 76900 143132 76906
rect 143080 76842 143132 76848
rect 143184 76809 143212 79630
rect 143170 76800 143226 76809
rect 143080 76764 143132 76770
rect 143170 76735 143226 76744
rect 143080 76706 143132 76712
rect 142986 76528 143042 76537
rect 142986 76463 143042 76472
rect 142816 71746 142936 71774
rect 142816 69018 142844 71746
rect 143092 69766 143120 76706
rect 143460 76673 143488 79784
rect 143552 79784 143626 79812
rect 143446 76664 143502 76673
rect 143446 76599 143502 76608
rect 143552 75914 143580 79784
rect 143690 79744 143718 80036
rect 143782 79937 143810 80036
rect 143768 79928 143824 79937
rect 143874 79898 143902 80036
rect 143768 79863 143824 79872
rect 143862 79892 143914 79898
rect 143862 79834 143914 79840
rect 143644 79716 143718 79744
rect 143814 79792 143870 79801
rect 143966 79778 143994 80036
rect 144058 79801 144086 80036
rect 143814 79727 143870 79736
rect 143920 79750 143994 79778
rect 144044 79792 144100 79801
rect 143644 79665 143672 79716
rect 143630 79656 143686 79665
rect 143630 79591 143686 79600
rect 143630 79520 143686 79529
rect 143630 79455 143686 79464
rect 143644 76022 143672 79455
rect 143724 78532 143776 78538
rect 143724 78474 143776 78480
rect 143632 76016 143684 76022
rect 143632 75958 143684 75964
rect 143552 75886 143672 75914
rect 143080 69760 143132 69766
rect 143080 69702 143132 69708
rect 142804 69012 142856 69018
rect 142804 68954 142856 68960
rect 142712 51740 142764 51746
rect 142712 51682 142764 51688
rect 142896 44940 142948 44946
rect 142896 44882 142948 44888
rect 142802 44296 142858 44305
rect 142802 44231 142858 44240
rect 142620 44192 142672 44198
rect 142620 44134 142672 44140
rect 142528 15904 142580 15910
rect 142528 15846 142580 15852
rect 142436 6248 142488 6254
rect 142436 6190 142488 6196
rect 142344 5024 142396 5030
rect 142344 4966 142396 4972
rect 142252 4956 142304 4962
rect 142252 4898 142304 4904
rect 142160 3800 142212 3806
rect 142160 3742 142212 3748
rect 142436 3732 142488 3738
rect 142436 3674 142488 3680
rect 141608 3596 141660 3602
rect 141608 3538 141660 3544
rect 142448 480 142476 3674
rect 142816 3262 142844 44231
rect 142908 3330 142936 44882
rect 143644 4894 143672 75886
rect 143736 5166 143764 78474
rect 143828 5234 143856 79727
rect 143920 78266 143948 79750
rect 144150 79778 144178 80036
rect 144242 79898 144270 80036
rect 144334 79966 144362 80036
rect 144426 79971 144454 80036
rect 144322 79960 144374 79966
rect 144322 79902 144374 79908
rect 144412 79962 144468 79971
rect 144230 79892 144282 79898
rect 144412 79897 144468 79906
rect 144230 79834 144282 79840
rect 144150 79750 144224 79778
rect 144044 79727 144100 79736
rect 144000 79688 144052 79694
rect 144000 79630 144052 79636
rect 143908 78260 143960 78266
rect 143908 78202 143960 78208
rect 143906 78160 143962 78169
rect 143906 78095 143962 78104
rect 143816 5228 143868 5234
rect 143816 5170 143868 5176
rect 143724 5160 143776 5166
rect 143724 5102 143776 5108
rect 143632 4888 143684 4894
rect 143632 4830 143684 4836
rect 143920 4826 143948 78095
rect 144012 6186 144040 79630
rect 144196 78538 144224 79750
rect 144518 79744 144546 80036
rect 144610 79801 144638 80036
rect 144702 79966 144730 80036
rect 144690 79960 144742 79966
rect 144690 79902 144742 79908
rect 144380 79716 144546 79744
rect 144596 79792 144652 79801
rect 144794 79744 144822 80036
rect 144886 79966 144914 80036
rect 144874 79960 144926 79966
rect 144874 79902 144926 79908
rect 144978 79812 145006 80036
rect 144596 79727 144652 79736
rect 144748 79716 144822 79744
rect 144932 79784 145006 79812
rect 144276 79688 144328 79694
rect 144276 79630 144328 79636
rect 144184 78532 144236 78538
rect 144184 78474 144236 78480
rect 144092 78260 144144 78266
rect 144092 78202 144144 78208
rect 144104 63306 144132 78202
rect 144288 78130 144316 79630
rect 144276 78124 144328 78130
rect 144276 78066 144328 78072
rect 144380 77874 144408 79716
rect 144644 79688 144696 79694
rect 144458 79656 144514 79665
rect 144644 79630 144696 79636
rect 144458 79591 144514 79600
rect 144552 79620 144604 79626
rect 144288 77846 144408 77874
rect 144288 70394 144316 77846
rect 144368 77784 144420 77790
rect 144368 77726 144420 77732
rect 144380 71058 144408 77726
rect 144472 76226 144500 79591
rect 144552 79562 144604 79568
rect 144460 76220 144512 76226
rect 144460 76162 144512 76168
rect 144460 76016 144512 76022
rect 144460 75958 144512 75964
rect 144368 71052 144420 71058
rect 144368 70994 144420 71000
rect 144196 70366 144316 70394
rect 144196 69970 144224 70366
rect 144184 69964 144236 69970
rect 144184 69906 144236 69912
rect 144182 66192 144238 66201
rect 144182 66127 144238 66136
rect 144092 63300 144144 63306
rect 144092 63242 144144 63248
rect 144000 6180 144052 6186
rect 144000 6122 144052 6128
rect 143908 4820 143960 4826
rect 143908 4762 143960 4768
rect 144196 3670 144224 66127
rect 144276 44192 144328 44198
rect 144276 44134 144328 44140
rect 144184 3664 144236 3670
rect 144184 3606 144236 3612
rect 143540 3596 143592 3602
rect 143540 3538 143592 3544
rect 142896 3324 142948 3330
rect 142896 3266 142948 3272
rect 142804 3256 142856 3262
rect 142804 3198 142856 3204
rect 143552 480 143580 3538
rect 144288 3534 144316 44134
rect 144472 3738 144500 75958
rect 144460 3732 144512 3738
rect 144460 3674 144512 3680
rect 144276 3528 144328 3534
rect 144276 3470 144328 3476
rect 144564 3466 144592 79562
rect 144656 75585 144684 79630
rect 144748 76673 144776 79716
rect 144932 79665 144960 79784
rect 145070 79744 145098 80036
rect 145162 79801 145190 80036
rect 145024 79716 145098 79744
rect 145148 79792 145204 79801
rect 145148 79727 145204 79736
rect 145254 79744 145282 80036
rect 145346 79898 145374 80036
rect 145334 79892 145386 79898
rect 145334 79834 145386 79840
rect 145438 79778 145466 80036
rect 145530 79830 145558 80036
rect 145622 79903 145650 80036
rect 145608 79894 145664 79903
rect 145392 79750 145466 79778
rect 145518 79824 145570 79830
rect 145608 79829 145664 79838
rect 145714 79812 145742 80036
rect 145806 79966 145834 80036
rect 145794 79960 145846 79966
rect 145794 79902 145846 79908
rect 145714 79801 145788 79812
rect 145714 79792 145802 79801
rect 145714 79784 145746 79792
rect 145518 79766 145570 79772
rect 145254 79716 145328 79744
rect 144918 79656 144974 79665
rect 144828 79620 144880 79626
rect 145024 79626 145052 79716
rect 144918 79591 144974 79600
rect 145012 79620 145064 79626
rect 144828 79562 144880 79568
rect 145012 79562 145064 79568
rect 145104 79620 145156 79626
rect 145300 79608 145328 79716
rect 145104 79562 145156 79568
rect 145208 79580 145328 79608
rect 144840 78169 144868 79562
rect 145010 79520 145066 79529
rect 145010 79455 145066 79464
rect 144920 79076 144972 79082
rect 144920 79018 144972 79024
rect 144932 78946 144960 79018
rect 144920 78940 144972 78946
rect 144920 78882 144972 78888
rect 144826 78160 144882 78169
rect 144826 78095 144882 78104
rect 144734 76664 144790 76673
rect 144734 76599 144790 76608
rect 144642 75576 144698 75585
rect 144642 75511 144698 75520
rect 145024 31414 145052 79455
rect 145116 34270 145144 79562
rect 145208 34338 145236 79580
rect 145286 79520 145342 79529
rect 145286 79455 145342 79464
rect 145300 77654 145328 79455
rect 145288 77648 145340 77654
rect 145288 77590 145340 77596
rect 145392 77314 145420 79750
rect 145898 79778 145926 80036
rect 145990 79966 146018 80036
rect 145978 79960 146030 79966
rect 145978 79902 146030 79908
rect 146082 79778 146110 80036
rect 146174 79898 146202 80036
rect 146162 79892 146214 79898
rect 146162 79834 146214 79840
rect 146266 79778 146294 80036
rect 146358 79903 146386 80036
rect 146344 79894 146400 79903
rect 146344 79829 146400 79838
rect 145746 79727 145802 79736
rect 145852 79750 145926 79778
rect 146036 79750 146110 79778
rect 146220 79750 146294 79778
rect 145656 79688 145708 79694
rect 145656 79630 145708 79636
rect 145748 79688 145800 79694
rect 145748 79630 145800 79636
rect 145472 79620 145524 79626
rect 145472 79562 145524 79568
rect 145484 77353 145512 79562
rect 145562 79520 145618 79529
rect 145562 79455 145618 79464
rect 145470 77344 145526 77353
rect 145380 77308 145432 77314
rect 145470 77279 145526 77288
rect 145380 77250 145432 77256
rect 145288 75268 145340 75274
rect 145288 75210 145340 75216
rect 145196 34332 145248 34338
rect 145196 34274 145248 34280
rect 145104 34264 145156 34270
rect 145104 34206 145156 34212
rect 145300 34202 145328 75210
rect 145576 70394 145604 79455
rect 145668 75614 145696 79630
rect 145760 78334 145788 79630
rect 145748 78328 145800 78334
rect 145748 78270 145800 78276
rect 145748 76220 145800 76226
rect 145748 76162 145800 76168
rect 145656 75608 145708 75614
rect 145656 75550 145708 75556
rect 145760 75138 145788 76162
rect 145748 75132 145800 75138
rect 145748 75074 145800 75080
rect 145392 70366 145604 70394
rect 145392 67182 145420 70366
rect 145564 69012 145616 69018
rect 145564 68954 145616 68960
rect 145380 67176 145432 67182
rect 145380 67118 145432 67124
rect 145288 34196 145340 34202
rect 145288 34138 145340 34144
rect 145012 31408 145064 31414
rect 145012 31350 145064 31356
rect 144736 4140 144788 4146
rect 144736 4082 144788 4088
rect 144552 3460 144604 3466
rect 144552 3402 144604 3408
rect 144748 480 144776 4082
rect 145576 2990 145604 68954
rect 145852 68542 145880 79750
rect 145932 79688 145984 79694
rect 145932 79630 145984 79636
rect 145944 77178 145972 79630
rect 145932 77172 145984 77178
rect 145932 77114 145984 77120
rect 146036 75274 146064 79750
rect 146114 79656 146170 79665
rect 146114 79591 146170 79600
rect 146024 75268 146076 75274
rect 146024 75210 146076 75216
rect 146024 75132 146076 75138
rect 146024 75074 146076 75080
rect 145840 68536 145892 68542
rect 145840 68478 145892 68484
rect 145656 63300 145708 63306
rect 145656 63242 145708 63248
rect 145668 3398 145696 63242
rect 146036 3602 146064 75074
rect 146128 27266 146156 79591
rect 146220 77489 146248 79750
rect 146450 79744 146478 80036
rect 146542 79898 146570 80036
rect 146530 79892 146582 79898
rect 146530 79834 146582 79840
rect 146634 79778 146662 80036
rect 146726 79966 146754 80036
rect 146714 79960 146766 79966
rect 146714 79902 146766 79908
rect 146818 79898 146846 80036
rect 146806 79892 146858 79898
rect 146806 79834 146858 79840
rect 146634 79750 146800 79778
rect 146450 79716 146524 79744
rect 146300 79688 146352 79694
rect 146300 79630 146352 79636
rect 146206 77480 146262 77489
rect 146206 77415 146262 77424
rect 146116 27260 146168 27266
rect 146116 27202 146168 27208
rect 146312 4146 146340 79630
rect 146392 79620 146444 79626
rect 146392 79562 146444 79568
rect 146300 4140 146352 4146
rect 146300 4082 146352 4088
rect 146404 4078 146432 79562
rect 146496 77994 146524 79716
rect 146576 79688 146628 79694
rect 146576 79630 146628 79636
rect 146668 79688 146720 79694
rect 146668 79630 146720 79636
rect 146484 77988 146536 77994
rect 146484 77930 146536 77936
rect 146484 75200 146536 75206
rect 146484 75142 146536 75148
rect 146496 25974 146524 75142
rect 146588 27198 146616 79630
rect 146680 28762 146708 79630
rect 146772 75274 146800 79750
rect 146910 79744 146938 80036
rect 147002 79898 147030 80036
rect 146990 79892 147042 79898
rect 146990 79834 147042 79840
rect 147094 79744 147122 80036
rect 146864 79716 146938 79744
rect 147048 79716 147122 79744
rect 146760 75268 146812 75274
rect 146760 75210 146812 75216
rect 146760 75132 146812 75138
rect 146760 75074 146812 75080
rect 146772 32910 146800 75074
rect 146864 35630 146892 79716
rect 146944 79620 146996 79626
rect 146944 79562 146996 79568
rect 146956 78033 146984 79562
rect 146942 78024 146998 78033
rect 146942 77959 146998 77968
rect 146944 75268 146996 75274
rect 146944 75210 146996 75216
rect 146956 35698 146984 75210
rect 147048 75206 147076 79716
rect 147186 79676 147214 80036
rect 147278 79937 147306 80036
rect 147370 79966 147398 80036
rect 147358 79960 147410 79966
rect 147264 79928 147320 79937
rect 147358 79902 147410 79908
rect 147264 79863 147320 79872
rect 147312 79824 147364 79830
rect 147462 79778 147490 80036
rect 147554 79830 147582 80036
rect 147312 79766 147364 79772
rect 147140 79648 147214 79676
rect 147036 75200 147088 75206
rect 147036 75142 147088 75148
rect 147140 75138 147168 79648
rect 147220 79008 147272 79014
rect 147220 78950 147272 78956
rect 147232 78878 147260 78950
rect 147220 78872 147272 78878
rect 147220 78814 147272 78820
rect 147324 77489 147352 79766
rect 147416 79750 147490 79778
rect 147542 79824 147594 79830
rect 147542 79766 147594 79772
rect 147310 77480 147366 77489
rect 147310 77415 147366 77424
rect 147416 77353 147444 79750
rect 147494 79656 147550 79665
rect 147646 79642 147674 80036
rect 147738 79830 147766 80036
rect 147726 79824 147778 79830
rect 147726 79766 147778 79772
rect 147830 79676 147858 80036
rect 147922 79744 147950 80036
rect 148014 79937 148042 80036
rect 148000 79928 148056 79937
rect 148000 79863 148056 79872
rect 148106 79830 148134 80036
rect 148198 79971 148226 80036
rect 148184 79962 148240 79971
rect 148290 79966 148318 80036
rect 148382 79966 148410 80036
rect 148474 79966 148502 80036
rect 148566 79966 148594 80036
rect 148184 79897 148240 79906
rect 148278 79960 148330 79966
rect 148278 79902 148330 79908
rect 148370 79960 148422 79966
rect 148370 79902 148422 79908
rect 148462 79960 148514 79966
rect 148462 79902 148514 79908
rect 148554 79960 148606 79966
rect 148658 79937 148686 80036
rect 148554 79902 148606 79908
rect 148644 79928 148700 79937
rect 148750 79898 148778 80036
rect 148644 79863 148700 79872
rect 148738 79892 148790 79898
rect 148738 79834 148790 79840
rect 148094 79824 148146 79830
rect 148094 79766 148146 79772
rect 148232 79824 148284 79830
rect 148842 79812 148870 80036
rect 148934 79966 148962 80036
rect 148922 79960 148974 79966
rect 148922 79902 148974 79908
rect 148842 79801 148916 79812
rect 148842 79792 148930 79801
rect 148842 79784 148874 79792
rect 148232 79766 148284 79772
rect 147922 79716 148042 79744
rect 147494 79591 147550 79600
rect 147600 79614 147674 79642
rect 147784 79648 147858 79676
rect 148014 79676 148042 79716
rect 148014 79648 148088 79676
rect 147402 77344 147458 77353
rect 147220 77308 147272 77314
rect 147402 77279 147458 77288
rect 147220 77250 147272 77256
rect 147128 75132 147180 75138
rect 147128 75074 147180 75080
rect 146944 35692 146996 35698
rect 146944 35634 146996 35640
rect 146852 35624 146904 35630
rect 146852 35566 146904 35572
rect 146760 32904 146812 32910
rect 146760 32846 146812 32852
rect 146668 28756 146720 28762
rect 146668 28698 146720 28704
rect 147232 27334 147260 77250
rect 147508 75546 147536 79591
rect 147600 76401 147628 79614
rect 147680 79416 147732 79422
rect 147680 79358 147732 79364
rect 147692 79082 147720 79358
rect 147680 79076 147732 79082
rect 147680 79018 147732 79024
rect 147586 76392 147642 76401
rect 147586 76327 147642 76336
rect 147496 75540 147548 75546
rect 147496 75482 147548 75488
rect 147220 27328 147272 27334
rect 147220 27270 147272 27276
rect 146576 27192 146628 27198
rect 146576 27134 146628 27140
rect 146484 25968 146536 25974
rect 146484 25910 146536 25916
rect 146392 4072 146444 4078
rect 146392 4014 146444 4020
rect 147784 4010 147812 79648
rect 147864 79552 147916 79558
rect 147864 79494 147916 79500
rect 147956 79552 148008 79558
rect 147956 79494 148008 79500
rect 147876 77722 147904 79494
rect 147864 77716 147916 77722
rect 147864 77658 147916 77664
rect 147864 76764 147916 76770
rect 147864 76706 147916 76712
rect 147876 6730 147904 76706
rect 147968 76498 147996 79494
rect 147956 76492 148008 76498
rect 147956 76434 148008 76440
rect 147956 76356 148008 76362
rect 147956 76298 148008 76304
rect 147968 28626 147996 76298
rect 148060 28694 148088 79648
rect 148140 76492 148192 76498
rect 148140 76434 148192 76440
rect 148152 32842 148180 76434
rect 148244 34134 148272 79766
rect 148416 79756 148468 79762
rect 148416 79698 148468 79704
rect 148508 79756 148560 79762
rect 149026 79744 149054 80036
rect 149118 79778 149146 80036
rect 149210 79966 149238 80036
rect 149198 79960 149250 79966
rect 149302 79937 149330 80036
rect 149198 79902 149250 79908
rect 149288 79928 149344 79937
rect 149394 79898 149422 80036
rect 149486 79898 149514 80036
rect 149578 79898 149606 80036
rect 149670 79937 149698 80036
rect 149656 79928 149712 79937
rect 149288 79863 149344 79872
rect 149382 79892 149434 79898
rect 149382 79834 149434 79840
rect 149474 79892 149526 79898
rect 149474 79834 149526 79840
rect 149566 79892 149618 79898
rect 149656 79863 149712 79872
rect 149566 79834 149618 79840
rect 149762 79812 149790 80036
rect 149716 79784 149790 79812
rect 149716 79778 149744 79784
rect 149118 79750 149192 79778
rect 148874 79727 148930 79736
rect 148508 79698 148560 79704
rect 148980 79716 149054 79744
rect 148322 78432 148378 78441
rect 148322 78367 148378 78376
rect 148336 75682 148364 78367
rect 148428 76770 148456 79698
rect 148416 76764 148468 76770
rect 148416 76706 148468 76712
rect 148414 76664 148470 76673
rect 148414 76599 148470 76608
rect 148324 75676 148376 75682
rect 148324 75618 148376 75624
rect 148322 75440 148378 75449
rect 148322 75375 148378 75384
rect 148336 49026 148364 75375
rect 148428 61606 148456 76599
rect 148520 76362 148548 79698
rect 148600 79688 148652 79694
rect 148600 79630 148652 79636
rect 148876 79688 148928 79694
rect 148876 79630 148928 79636
rect 148508 76356 148560 76362
rect 148508 76298 148560 76304
rect 148612 74118 148640 79630
rect 148692 79620 148744 79626
rect 148692 79562 148744 79568
rect 148704 77217 148732 79562
rect 148784 79552 148836 79558
rect 148784 79494 148836 79500
rect 148690 77208 148746 77217
rect 148690 77143 148746 77152
rect 148600 74112 148652 74118
rect 148600 74054 148652 74060
rect 148796 73154 148824 79494
rect 148888 75177 148916 79630
rect 148980 76673 149008 79716
rect 149058 79520 149114 79529
rect 149058 79455 149114 79464
rect 148966 76664 149022 76673
rect 148966 76599 149022 76608
rect 148874 75168 148930 75177
rect 148874 75103 148930 75112
rect 148704 73126 148824 73154
rect 148704 64874 148732 73126
rect 148612 64846 148732 64874
rect 148416 61600 148468 61606
rect 148416 61542 148468 61548
rect 148324 49020 148376 49026
rect 148324 48962 148376 48968
rect 148232 34128 148284 34134
rect 148232 34070 148284 34076
rect 148140 32836 148192 32842
rect 148140 32778 148192 32784
rect 148048 28688 148100 28694
rect 148048 28630 148100 28636
rect 147956 28620 148008 28626
rect 147956 28562 148008 28568
rect 147864 6724 147916 6730
rect 147864 6666 147916 6672
rect 147772 4004 147824 4010
rect 147772 3946 147824 3952
rect 148612 3874 148640 64846
rect 149072 6526 149100 79455
rect 149164 76294 149192 79750
rect 149244 79756 149296 79762
rect 149244 79698 149296 79704
rect 149336 79756 149388 79762
rect 149336 79698 149388 79704
rect 149624 79750 149744 79778
rect 149152 76288 149204 76294
rect 149152 76230 149204 76236
rect 149152 76152 149204 76158
rect 149152 76094 149204 76100
rect 149164 6594 149192 76094
rect 149256 6662 149284 79698
rect 149348 76498 149376 79698
rect 149520 79688 149572 79694
rect 149520 79630 149572 79636
rect 149428 79620 149480 79626
rect 149428 79562 149480 79568
rect 149336 76492 149388 76498
rect 149336 76434 149388 76440
rect 149440 76158 149468 79562
rect 149428 76152 149480 76158
rect 149428 76094 149480 76100
rect 149428 75132 149480 75138
rect 149428 75074 149480 75080
rect 149336 75064 149388 75070
rect 149336 75006 149388 75012
rect 149244 6656 149296 6662
rect 149244 6598 149296 6604
rect 149152 6588 149204 6594
rect 149152 6530 149204 6536
rect 149060 6520 149112 6526
rect 149060 6462 149112 6468
rect 149348 6458 149376 75006
rect 149440 13530 149468 75074
rect 149532 29986 149560 79630
rect 149624 79529 149652 79750
rect 149854 79744 149882 80036
rect 149808 79716 149882 79744
rect 149946 79744 149974 80036
rect 150038 79971 150066 80036
rect 150024 79962 150080 79971
rect 150024 79897 150080 79906
rect 150130 79812 150158 80036
rect 150222 79971 150250 80036
rect 150208 79962 150264 79971
rect 150208 79897 150264 79906
rect 150314 79830 150342 80036
rect 150302 79824 150354 79830
rect 150130 79801 150204 79812
rect 150130 79792 150218 79801
rect 150130 79784 150162 79792
rect 149946 79716 150020 79744
rect 150302 79766 150354 79772
rect 150162 79727 150218 79736
rect 149702 79656 149758 79665
rect 149702 79591 149758 79600
rect 149610 79520 149666 79529
rect 149610 79455 149666 79464
rect 149612 79348 149664 79354
rect 149612 79290 149664 79296
rect 149624 78985 149652 79290
rect 149610 78976 149666 78985
rect 149610 78911 149666 78920
rect 149716 78606 149744 79591
rect 149704 78600 149756 78606
rect 149704 78542 149756 78548
rect 149808 76616 149836 79716
rect 149624 76588 149836 76616
rect 149520 29980 149572 29986
rect 149520 29922 149572 29928
rect 149624 29918 149652 76588
rect 149796 76492 149848 76498
rect 149796 76434 149848 76440
rect 149704 76288 149756 76294
rect 149704 76230 149756 76236
rect 149716 32774 149744 76230
rect 149808 34066 149836 76434
rect 149992 75138 150020 79716
rect 150164 79688 150216 79694
rect 150070 79656 150126 79665
rect 150406 79676 150434 80036
rect 150498 79830 150526 80036
rect 150590 79971 150618 80036
rect 150576 79962 150632 79971
rect 150576 79897 150632 79906
rect 150682 79830 150710 80036
rect 150774 79971 150802 80036
rect 150760 79962 150816 79971
rect 150866 79966 150894 80036
rect 150760 79897 150816 79906
rect 150854 79960 150906 79966
rect 150958 79937 150986 80036
rect 151050 79966 151078 80036
rect 151142 79971 151170 80036
rect 151038 79960 151090 79966
rect 150854 79902 150906 79908
rect 150944 79928 151000 79937
rect 151038 79902 151090 79908
rect 151128 79962 151184 79971
rect 151128 79897 151184 79906
rect 150944 79863 151000 79872
rect 150486 79824 150538 79830
rect 150486 79766 150538 79772
rect 150670 79824 150722 79830
rect 151084 79824 151136 79830
rect 150670 79766 150722 79772
rect 150806 79792 150862 79801
rect 150862 79750 150940 79778
rect 151084 79766 151136 79772
rect 150806 79727 150862 79736
rect 150164 79630 150216 79636
rect 150360 79648 150434 79676
rect 150716 79688 150768 79694
rect 150070 79591 150126 79600
rect 150084 75914 150112 79591
rect 150176 78713 150204 79630
rect 150254 79520 150310 79529
rect 150254 79455 150310 79464
rect 150162 78704 150218 78713
rect 150162 78639 150218 78648
rect 150084 75886 150204 75914
rect 149980 75132 150032 75138
rect 149980 75074 150032 75080
rect 150176 75070 150204 75886
rect 150164 75064 150216 75070
rect 150164 75006 150216 75012
rect 150268 74186 150296 79455
rect 150360 77081 150388 79648
rect 150716 79630 150768 79636
rect 150806 79656 150862 79665
rect 150624 79620 150676 79626
rect 150624 79562 150676 79568
rect 150532 79144 150584 79150
rect 150532 79086 150584 79092
rect 150544 78810 150572 79086
rect 150532 78804 150584 78810
rect 150532 78746 150584 78752
rect 150440 77240 150492 77246
rect 150440 77182 150492 77188
rect 150346 77072 150402 77081
rect 150346 77007 150402 77016
rect 150256 74180 150308 74186
rect 150256 74122 150308 74128
rect 149796 34060 149848 34066
rect 149796 34002 149848 34008
rect 149704 32768 149756 32774
rect 149704 32710 149756 32716
rect 149612 29912 149664 29918
rect 149612 29854 149664 29860
rect 149428 13524 149480 13530
rect 149428 13466 149480 13472
rect 149336 6452 149388 6458
rect 149336 6394 149388 6400
rect 150452 6390 150480 77182
rect 150532 76900 150584 76906
rect 150532 76842 150584 76848
rect 150544 8838 150572 76842
rect 150636 76752 150664 79562
rect 150728 76906 150756 79630
rect 150806 79591 150862 79600
rect 150820 77790 150848 79591
rect 150808 77784 150860 77790
rect 150808 77726 150860 77732
rect 150716 76900 150768 76906
rect 150716 76842 150768 76848
rect 150912 76820 150940 79750
rect 150992 79756 151044 79762
rect 150992 79698 151044 79704
rect 151004 77024 151032 79698
rect 151096 77246 151124 79766
rect 151234 79744 151262 80036
rect 151326 79778 151354 80036
rect 151418 79971 151446 80036
rect 151404 79962 151460 79971
rect 151404 79897 151460 79906
rect 151326 79750 151400 79778
rect 151188 79716 151262 79744
rect 151084 77240 151136 77246
rect 151084 77182 151136 77188
rect 151004 76996 151124 77024
rect 150912 76792 151032 76820
rect 150636 76724 150940 76752
rect 150622 76664 150678 76673
rect 150622 76599 150678 76608
rect 150636 8906 150664 76599
rect 150716 75948 150768 75954
rect 150716 75890 150768 75896
rect 150728 15026 150756 75890
rect 150808 75880 150860 75886
rect 150808 75822 150860 75828
rect 150820 29850 150848 75822
rect 150912 35562 150940 76724
rect 151004 74050 151032 76792
rect 151096 75954 151124 76996
rect 151084 75948 151136 75954
rect 151084 75890 151136 75896
rect 151188 75886 151216 79716
rect 151372 78130 151400 79750
rect 151510 79744 151538 80036
rect 151464 79716 151538 79744
rect 151602 79744 151630 80036
rect 151694 79971 151722 80036
rect 151680 79962 151736 79971
rect 151680 79897 151736 79906
rect 151786 79812 151814 80036
rect 151878 79966 151906 80036
rect 151866 79960 151918 79966
rect 151866 79902 151918 79908
rect 151970 79812 151998 80036
rect 151786 79801 151860 79812
rect 151786 79792 151874 79801
rect 151786 79784 151818 79792
rect 151602 79716 151768 79744
rect 151818 79727 151874 79736
rect 151924 79784 151998 79812
rect 151360 78124 151412 78130
rect 151360 78066 151412 78072
rect 151360 77988 151412 77994
rect 151360 77930 151412 77936
rect 151176 75880 151228 75886
rect 151176 75822 151228 75828
rect 150992 74044 151044 74050
rect 150992 73986 151044 73992
rect 151084 69760 151136 69766
rect 151084 69702 151136 69708
rect 150900 35556 150952 35562
rect 150900 35498 150952 35504
rect 150808 29844 150860 29850
rect 150808 29786 150860 29792
rect 150716 15020 150768 15026
rect 150716 14962 150768 14968
rect 150624 8900 150676 8906
rect 150624 8842 150676 8848
rect 150532 8832 150584 8838
rect 150532 8774 150584 8780
rect 150440 6384 150492 6390
rect 150440 6326 150492 6332
rect 147128 3868 147180 3874
rect 147128 3810 147180 3816
rect 148600 3868 148652 3874
rect 148600 3810 148652 3816
rect 146024 3596 146076 3602
rect 146024 3538 146076 3544
rect 145656 3392 145708 3398
rect 145656 3334 145708 3340
rect 145932 3324 145984 3330
rect 145932 3266 145984 3272
rect 145564 2984 145616 2990
rect 145564 2926 145616 2932
rect 145944 480 145972 3266
rect 147140 480 147168 3810
rect 151096 3602 151124 69702
rect 151372 64874 151400 77930
rect 151464 76974 151492 79716
rect 151634 79656 151690 79665
rect 151544 79620 151596 79626
rect 151634 79591 151690 79600
rect 151544 79562 151596 79568
rect 151452 76968 151504 76974
rect 151452 76910 151504 76916
rect 151556 73914 151584 79562
rect 151648 77858 151676 79591
rect 151636 77852 151688 77858
rect 151636 77794 151688 77800
rect 151740 76673 151768 79716
rect 151818 79656 151874 79665
rect 151818 79591 151874 79600
rect 151726 76664 151782 76673
rect 151726 76599 151782 76608
rect 151544 73908 151596 73914
rect 151544 73850 151596 73856
rect 151280 64846 151400 64874
rect 151084 3596 151136 3602
rect 151084 3538 151136 3544
rect 149520 3528 149572 3534
rect 149520 3470 149572 3476
rect 148324 3256 148376 3262
rect 148324 3198 148376 3204
rect 148336 480 148364 3198
rect 149532 480 149560 3470
rect 151280 3398 151308 64846
rect 151832 9654 151860 79591
rect 151924 78674 151952 79784
rect 152062 79744 152090 80036
rect 152016 79716 152090 79744
rect 151912 78668 151964 78674
rect 151912 78610 151964 78616
rect 151912 77308 151964 77314
rect 151912 77250 151964 77256
rect 151820 9648 151872 9654
rect 151820 9590 151872 9596
rect 151924 9586 151952 77250
rect 152016 75818 152044 79716
rect 152154 79676 152182 80036
rect 152246 79744 152274 80036
rect 152338 79898 152366 80036
rect 152430 79966 152458 80036
rect 152418 79960 152470 79966
rect 152522 79937 152550 80036
rect 152418 79902 152470 79908
rect 152508 79928 152564 79937
rect 152326 79892 152378 79898
rect 152508 79863 152564 79872
rect 152326 79834 152378 79840
rect 152418 79824 152470 79830
rect 152470 79772 152550 79778
rect 152418 79766 152550 79772
rect 152430 79750 152550 79766
rect 152246 79716 152320 79744
rect 152108 79648 152182 79676
rect 152004 75812 152056 75818
rect 152004 75754 152056 75760
rect 152004 75132 152056 75138
rect 152004 75074 152056 75080
rect 152016 20262 152044 75074
rect 152108 20330 152136 79648
rect 152292 76430 152320 79716
rect 152372 79688 152424 79694
rect 152522 79676 152550 79750
rect 152372 79630 152424 79636
rect 152476 79648 152550 79676
rect 152280 76424 152332 76430
rect 152280 76366 152332 76372
rect 152188 75880 152240 75886
rect 152188 75822 152240 75828
rect 152200 25906 152228 75822
rect 152280 75812 152332 75818
rect 152280 75754 152332 75760
rect 152292 27130 152320 75754
rect 152384 28558 152412 79630
rect 152476 33998 152504 79648
rect 152614 79608 152642 80036
rect 152706 79744 152734 80036
rect 152798 79812 152826 80036
rect 152890 79966 152918 80036
rect 152982 79966 153010 80036
rect 152878 79960 152930 79966
rect 152878 79902 152930 79908
rect 152970 79960 153022 79966
rect 153074 79937 153102 80036
rect 152970 79902 153022 79908
rect 153060 79928 153116 79937
rect 153060 79863 153116 79872
rect 153016 79824 153068 79830
rect 152798 79784 152964 79812
rect 152706 79716 152826 79744
rect 152614 79580 152688 79608
rect 152556 76424 152608 76430
rect 152556 76366 152608 76372
rect 152568 61538 152596 76366
rect 152660 75886 152688 79580
rect 152798 79540 152826 79716
rect 152752 79512 152826 79540
rect 152648 75880 152700 75886
rect 152648 75822 152700 75828
rect 152752 75138 152780 79512
rect 152936 77314 152964 79784
rect 153166 79778 153194 80036
rect 153016 79766 153068 79772
rect 153028 77353 153056 79766
rect 153120 79750 153194 79778
rect 153014 77344 153070 77353
rect 152924 77308 152976 77314
rect 153014 77279 153070 77288
rect 152924 77250 152976 77256
rect 153120 76945 153148 79750
rect 153258 79676 153286 80036
rect 153350 79971 153378 80036
rect 153336 79962 153392 79971
rect 153442 79966 153470 80036
rect 153336 79897 153392 79906
rect 153430 79960 153482 79966
rect 153534 79937 153562 80036
rect 153626 79966 153654 80036
rect 153718 79971 153746 80036
rect 153614 79960 153666 79966
rect 153430 79902 153482 79908
rect 153520 79928 153576 79937
rect 153614 79902 153666 79908
rect 153704 79962 153760 79971
rect 153704 79897 153760 79906
rect 153810 79898 153838 80036
rect 153902 79966 153930 80036
rect 153994 79966 154022 80036
rect 154086 79966 154114 80036
rect 154178 79971 154206 80036
rect 153890 79960 153942 79966
rect 153890 79902 153942 79908
rect 153982 79960 154034 79966
rect 153982 79902 154034 79908
rect 154074 79960 154126 79966
rect 154074 79902 154126 79908
rect 154164 79962 154220 79971
rect 153520 79863 153576 79872
rect 153798 79892 153850 79898
rect 154164 79897 154220 79906
rect 153798 79834 153850 79840
rect 154270 79830 154298 80036
rect 154362 79966 154390 80036
rect 154350 79960 154402 79966
rect 154350 79902 154402 79908
rect 154166 79824 154218 79830
rect 153382 79792 153438 79801
rect 154086 79772 154166 79778
rect 154086 79766 154218 79772
rect 154258 79824 154310 79830
rect 154258 79766 154310 79772
rect 153382 79727 153438 79736
rect 153844 79756 153896 79762
rect 153212 79648 153286 79676
rect 153212 77246 153240 79648
rect 153292 79552 153344 79558
rect 153292 79494 153344 79500
rect 153304 77489 153332 79494
rect 153396 78538 153424 79727
rect 154086 79750 154206 79766
rect 153896 79716 153976 79744
rect 153844 79698 153896 79704
rect 153752 79688 153804 79694
rect 153752 79630 153804 79636
rect 153842 79656 153898 79665
rect 153568 79620 153620 79626
rect 153568 79562 153620 79568
rect 153476 79484 153528 79490
rect 153476 79426 153528 79432
rect 153488 79286 153516 79426
rect 153476 79280 153528 79286
rect 153476 79222 153528 79228
rect 153384 78532 153436 78538
rect 153384 78474 153436 78480
rect 153290 77480 153346 77489
rect 153290 77415 153346 77424
rect 153474 77344 153530 77353
rect 153384 77308 153436 77314
rect 153474 77279 153530 77288
rect 153384 77250 153436 77256
rect 153200 77240 153252 77246
rect 153200 77182 153252 77188
rect 153106 76936 153162 76945
rect 153106 76871 153162 76880
rect 153290 76664 153346 76673
rect 153290 76599 153346 76608
rect 153200 75472 153252 75478
rect 153200 75414 153252 75420
rect 152740 75132 152792 75138
rect 152740 75074 152792 75080
rect 152556 61532 152608 61538
rect 152556 61474 152608 61480
rect 152464 33992 152516 33998
rect 152464 33934 152516 33940
rect 152372 28552 152424 28558
rect 152372 28494 152424 28500
rect 152280 27124 152332 27130
rect 152280 27066 152332 27072
rect 152188 25900 152240 25906
rect 152188 25842 152240 25848
rect 152096 20324 152148 20330
rect 152096 20266 152148 20272
rect 152004 20256 152056 20262
rect 152004 20198 152056 20204
rect 153212 10742 153240 75414
rect 153200 10736 153252 10742
rect 153200 10678 153252 10684
rect 153304 10606 153332 76599
rect 153396 10674 153424 77250
rect 153488 24410 153516 77279
rect 153580 31278 153608 79562
rect 153660 79552 153712 79558
rect 153660 79494 153712 79500
rect 153672 31346 153700 79494
rect 153764 79200 153792 79630
rect 153842 79591 153898 79600
rect 153856 79268 153884 79591
rect 153948 79370 153976 79716
rect 154086 79676 154114 79750
rect 154212 79688 154264 79694
rect 154086 79648 154160 79676
rect 153948 79342 154068 79370
rect 153856 79240 153976 79268
rect 153764 79172 153884 79200
rect 153752 77240 153804 77246
rect 153752 77182 153804 77188
rect 153764 33930 153792 77182
rect 153856 65958 153884 79172
rect 153948 72826 153976 79240
rect 154040 75478 154068 79342
rect 154132 77314 154160 79648
rect 154454 79676 154482 80036
rect 154546 79801 154574 80036
rect 154638 79937 154666 80036
rect 154624 79928 154680 79937
rect 154730 79898 154758 80036
rect 154822 79966 154850 80036
rect 154810 79960 154862 79966
rect 154810 79902 154862 79908
rect 154624 79863 154680 79872
rect 154718 79892 154770 79898
rect 154718 79834 154770 79840
rect 154914 79812 154942 80036
rect 154532 79792 154588 79801
rect 154532 79727 154588 79736
rect 154868 79784 154942 79812
rect 154408 79648 154482 79676
rect 154764 79688 154816 79694
rect 154408 79642 154436 79648
rect 154212 79630 154264 79636
rect 154120 77308 154172 77314
rect 154120 77250 154172 77256
rect 154224 76809 154252 79630
rect 154316 79614 154436 79642
rect 154764 79630 154816 79636
rect 154580 79620 154632 79626
rect 154316 77353 154344 79614
rect 154580 79562 154632 79568
rect 154396 79552 154448 79558
rect 154396 79494 154448 79500
rect 154488 79552 154540 79558
rect 154488 79494 154540 79500
rect 154302 77344 154358 77353
rect 154302 77279 154358 77288
rect 154210 76800 154266 76809
rect 154210 76735 154266 76744
rect 154028 75472 154080 75478
rect 154028 75414 154080 75420
rect 153936 72820 153988 72826
rect 153936 72762 153988 72768
rect 154408 72758 154436 79494
rect 154500 77489 154528 79494
rect 154486 77480 154542 77489
rect 154486 77415 154542 77424
rect 154592 77314 154620 79562
rect 154672 79552 154724 79558
rect 154672 79494 154724 79500
rect 154580 77308 154632 77314
rect 154580 77250 154632 77256
rect 154580 76356 154632 76362
rect 154580 76298 154632 76304
rect 154396 72752 154448 72758
rect 154396 72694 154448 72700
rect 153844 65952 153896 65958
rect 153844 65894 153896 65900
rect 153844 51740 153896 51746
rect 153844 51682 153896 51688
rect 153752 33924 153804 33930
rect 153752 33866 153804 33872
rect 153660 31340 153712 31346
rect 153660 31282 153712 31288
rect 153568 31272 153620 31278
rect 153568 31214 153620 31220
rect 153476 24404 153528 24410
rect 153476 24346 153528 24352
rect 153384 10668 153436 10674
rect 153384 10610 153436 10616
rect 153292 10600 153344 10606
rect 153292 10542 153344 10548
rect 151912 9580 151964 9586
rect 151912 9522 151964 9528
rect 151820 5024 151872 5030
rect 151820 4966 151872 4972
rect 151268 3392 151320 3398
rect 151268 3334 151320 3340
rect 150624 2984 150676 2990
rect 150624 2926 150676 2932
rect 150636 480 150664 2926
rect 151832 480 151860 4966
rect 153016 3596 153068 3602
rect 153016 3538 153068 3544
rect 153028 480 153056 3538
rect 153856 3262 153884 51682
rect 154592 12374 154620 76298
rect 154684 17474 154712 79494
rect 154776 77246 154804 79630
rect 154868 79529 154896 79784
rect 155006 79744 155034 80036
rect 155098 79937 155126 80036
rect 155084 79928 155140 79937
rect 155084 79863 155140 79872
rect 154960 79716 155034 79744
rect 154854 79520 154910 79529
rect 154854 79455 154910 79464
rect 154854 78160 154910 78169
rect 154854 78095 154910 78104
rect 154764 77240 154816 77246
rect 154764 77182 154816 77188
rect 154764 76628 154816 76634
rect 154764 76570 154816 76576
rect 154776 24342 154804 76570
rect 154868 25838 154896 78095
rect 154960 77994 154988 79716
rect 155190 79676 155218 80036
rect 155282 79966 155310 80036
rect 155270 79960 155322 79966
rect 155270 79902 155322 79908
rect 155374 79801 155402 80036
rect 155466 79830 155494 80036
rect 155454 79824 155506 79830
rect 155360 79792 155416 79801
rect 155454 79766 155506 79772
rect 155360 79727 155416 79736
rect 155316 79688 155368 79694
rect 155038 79656 155094 79665
rect 155190 79648 155264 79676
rect 155038 79591 155094 79600
rect 154948 77988 155000 77994
rect 154948 77930 155000 77936
rect 154948 77308 155000 77314
rect 154948 77250 155000 77256
rect 154960 28490 154988 77250
rect 155052 29782 155080 79591
rect 155130 79520 155186 79529
rect 155130 79455 155186 79464
rect 155144 35494 155172 79455
rect 155236 77450 155264 79648
rect 155558 79676 155586 80036
rect 155650 79744 155678 80036
rect 155742 79812 155770 80036
rect 155834 79971 155862 80036
rect 155820 79962 155876 79971
rect 155820 79897 155876 79906
rect 155926 79812 155954 80036
rect 155742 79784 155816 79812
rect 155650 79716 155724 79744
rect 155316 79630 155368 79636
rect 155512 79648 155586 79676
rect 155328 78266 155356 79630
rect 155406 79520 155462 79529
rect 155406 79455 155462 79464
rect 155316 78260 155368 78266
rect 155316 78202 155368 78208
rect 155316 78124 155368 78130
rect 155316 78066 155368 78072
rect 155224 77444 155276 77450
rect 155224 77386 155276 77392
rect 155222 77344 155278 77353
rect 155222 77279 155278 77288
rect 155236 65890 155264 77279
rect 155328 73982 155356 78066
rect 155420 74534 155448 79455
rect 155512 76362 155540 79648
rect 155696 78418 155724 79716
rect 155788 79529 155816 79784
rect 155880 79784 155954 79812
rect 155774 79520 155830 79529
rect 155774 79455 155830 79464
rect 155604 78390 155724 78418
rect 155774 78432 155830 78441
rect 155604 76634 155632 78390
rect 155774 78367 155830 78376
rect 155788 78334 155816 78367
rect 155776 78328 155828 78334
rect 155776 78270 155828 78276
rect 155776 77444 155828 77450
rect 155776 77386 155828 77392
rect 155592 76628 155644 76634
rect 155592 76570 155644 76576
rect 155500 76356 155552 76362
rect 155500 76298 155552 76304
rect 155420 74506 155724 74534
rect 155316 73976 155368 73982
rect 155316 73918 155368 73924
rect 155696 72622 155724 74506
rect 155788 72690 155816 77386
rect 155880 76673 155908 79784
rect 156018 79744 156046 80036
rect 156110 79966 156138 80036
rect 156098 79960 156150 79966
rect 156098 79902 156150 79908
rect 156202 79812 156230 80036
rect 156156 79801 156230 79812
rect 155972 79716 156046 79744
rect 156142 79792 156230 79801
rect 156198 79784 156230 79792
rect 156294 79744 156322 80036
rect 156386 79966 156414 80036
rect 156374 79960 156426 79966
rect 156374 79902 156426 79908
rect 156478 79898 156506 80036
rect 156570 79937 156598 80036
rect 156556 79928 156612 79937
rect 156466 79892 156518 79898
rect 156556 79863 156612 79872
rect 156466 79834 156518 79840
rect 156374 79824 156426 79830
rect 156426 79772 156460 79778
rect 156374 79766 156460 79772
rect 156386 79750 156460 79766
rect 156142 79727 156198 79736
rect 156248 79716 156322 79744
rect 155866 76664 155922 76673
rect 155972 76634 156000 79716
rect 156248 79665 156276 79716
rect 156234 79656 156290 79665
rect 156052 79620 156104 79626
rect 156052 79562 156104 79568
rect 156144 79620 156196 79626
rect 156234 79591 156290 79600
rect 156144 79562 156196 79568
rect 155866 76599 155922 76608
rect 155960 76628 156012 76634
rect 155960 76570 156012 76576
rect 155776 72684 155828 72690
rect 155776 72626 155828 72632
rect 155684 72616 155736 72622
rect 155684 72558 155736 72564
rect 155224 65884 155276 65890
rect 155224 65826 155276 65832
rect 155132 35488 155184 35494
rect 155132 35430 155184 35436
rect 155040 29776 155092 29782
rect 155040 29718 155092 29724
rect 154948 28484 155000 28490
rect 154948 28426 155000 28432
rect 154856 25832 154908 25838
rect 154856 25774 154908 25780
rect 154764 24336 154816 24342
rect 154764 24278 154816 24284
rect 154672 17468 154724 17474
rect 154672 17410 154724 17416
rect 156064 16574 156092 79562
rect 155972 16546 156092 16574
rect 154580 12368 154632 12374
rect 154580 12310 154632 12316
rect 155972 9518 156000 16546
rect 156156 15994 156184 79562
rect 156236 79552 156288 79558
rect 156236 79494 156288 79500
rect 156248 79014 156276 79494
rect 156236 79008 156288 79014
rect 156236 78950 156288 78956
rect 156432 77432 156460 79750
rect 156662 79676 156690 80036
rect 156754 79898 156782 80036
rect 156846 79966 156874 80036
rect 156938 79966 156966 80036
rect 156834 79960 156886 79966
rect 156834 79902 156886 79908
rect 156926 79960 156978 79966
rect 156926 79902 156978 79908
rect 156742 79892 156794 79898
rect 156742 79834 156794 79840
rect 156878 79792 156934 79801
rect 156788 79756 156840 79762
rect 156878 79727 156934 79736
rect 157030 79744 157058 80036
rect 157122 79971 157150 80036
rect 157108 79962 157164 79971
rect 157108 79897 157164 79906
rect 157214 79778 157242 80036
rect 157306 79898 157334 80036
rect 157294 79892 157346 79898
rect 157294 79834 157346 79840
rect 157214 79750 157288 79778
rect 156788 79698 156840 79704
rect 156510 79656 156566 79665
rect 156510 79591 156566 79600
rect 156616 79648 156690 79676
rect 156064 15966 156184 15994
rect 156248 77404 156460 77432
rect 156064 12034 156092 15966
rect 156144 15904 156196 15910
rect 156144 15846 156196 15852
rect 156052 12028 156104 12034
rect 156052 11970 156104 11976
rect 155960 9512 156012 9518
rect 155960 9454 156012 9460
rect 155408 6248 155460 6254
rect 155408 6190 155460 6196
rect 154212 3800 154264 3806
rect 154212 3742 154264 3748
rect 153844 3256 153896 3262
rect 153844 3198 153896 3204
rect 154224 480 154252 3742
rect 155420 480 155448 6190
rect 141210 326 141464 354
rect 141210 -960 141322 326
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156156 354 156184 15846
rect 156248 12170 156276 77404
rect 156326 77344 156382 77353
rect 156326 77279 156382 77288
rect 156236 12164 156288 12170
rect 156236 12106 156288 12112
rect 156340 12102 156368 77279
rect 156420 76628 156472 76634
rect 156420 76570 156472 76576
rect 156432 12306 156460 76570
rect 156420 12300 156472 12306
rect 156420 12242 156472 12248
rect 156524 12238 156552 79591
rect 156616 58682 156644 79648
rect 156696 79552 156748 79558
rect 156694 79520 156696 79529
rect 156748 79520 156750 79529
rect 156694 79455 156750 79464
rect 156696 78600 156748 78606
rect 156696 78542 156748 78548
rect 156708 77042 156736 78542
rect 156696 77036 156748 77042
rect 156696 76978 156748 76984
rect 156800 70394 156828 79698
rect 156892 76838 156920 79727
rect 157030 79716 157104 79744
rect 157076 78742 157104 79716
rect 157156 79620 157208 79626
rect 157156 79562 157208 79568
rect 157064 78736 157116 78742
rect 157064 78678 157116 78684
rect 157168 77489 157196 79562
rect 157260 77625 157288 79750
rect 157398 79608 157426 80036
rect 157490 79676 157518 80036
rect 157582 79812 157610 80036
rect 157674 79966 157702 80036
rect 157662 79960 157714 79966
rect 157662 79902 157714 79908
rect 157582 79784 157656 79812
rect 157490 79648 157564 79676
rect 157398 79580 157472 79608
rect 157338 79520 157394 79529
rect 157338 79455 157394 79464
rect 157246 77616 157302 77625
rect 157246 77551 157302 77560
rect 157154 77480 157210 77489
rect 157154 77415 157210 77424
rect 156880 76832 156932 76838
rect 156880 76774 156932 76780
rect 156800 70366 157012 70394
rect 156604 58676 156656 58682
rect 156604 58618 156656 58624
rect 156512 12232 156564 12238
rect 156512 12174 156564 12180
rect 156328 12096 156380 12102
rect 156328 12038 156380 12044
rect 156984 9450 157012 70366
rect 157352 10470 157380 79455
rect 157444 76906 157472 79580
rect 157536 77294 157564 79648
rect 157628 78962 157656 79784
rect 157766 79744 157794 80036
rect 157858 79937 157886 80036
rect 157844 79928 157900 79937
rect 157844 79863 157900 79872
rect 157950 79778 157978 80036
rect 158042 79966 158070 80036
rect 158030 79960 158082 79966
rect 158030 79902 158082 79908
rect 157950 79750 158024 79778
rect 157720 79716 157794 79744
rect 157720 79132 157748 79716
rect 157800 79620 157852 79626
rect 157800 79562 157852 79568
rect 157812 79286 157840 79562
rect 157800 79280 157852 79286
rect 157800 79222 157852 79228
rect 157720 79104 157932 79132
rect 157628 78934 157840 78962
rect 157708 78872 157760 78878
rect 157708 78814 157760 78820
rect 157536 77266 157656 77294
rect 157524 77036 157576 77042
rect 157524 76978 157576 76984
rect 157432 76900 157484 76906
rect 157432 76842 157484 76848
rect 157432 76764 157484 76770
rect 157432 76706 157484 76712
rect 157444 10538 157472 76706
rect 157536 13394 157564 76978
rect 157628 13462 157656 77266
rect 157720 33862 157748 78814
rect 157812 55894 157840 78934
rect 157904 75070 157932 79104
rect 157996 78878 158024 79750
rect 158134 79744 158162 80036
rect 158226 79898 158254 80036
rect 158318 79971 158346 80036
rect 158304 79962 158360 79971
rect 158214 79892 158266 79898
rect 158304 79897 158360 79906
rect 158410 79898 158438 80036
rect 158502 79966 158530 80036
rect 158490 79960 158542 79966
rect 158594 79937 158622 80036
rect 158490 79902 158542 79908
rect 158580 79928 158636 79937
rect 158214 79834 158266 79840
rect 158398 79892 158450 79898
rect 158580 79863 158636 79872
rect 158398 79834 158450 79840
rect 158352 79756 158404 79762
rect 158134 79716 158208 79744
rect 158076 79620 158128 79626
rect 158076 79562 158128 79568
rect 157984 78872 158036 78878
rect 157984 78814 158036 78820
rect 157984 78736 158036 78742
rect 157984 78678 158036 78684
rect 157892 75064 157944 75070
rect 157892 75006 157944 75012
rect 157996 70394 158024 78678
rect 158088 77042 158116 79562
rect 158076 77036 158128 77042
rect 158076 76978 158128 76984
rect 158180 76770 158208 79716
rect 158686 79744 158714 80036
rect 158778 79966 158806 80036
rect 158870 79966 158898 80036
rect 158766 79960 158818 79966
rect 158766 79902 158818 79908
rect 158858 79960 158910 79966
rect 158858 79902 158910 79908
rect 158812 79756 158864 79762
rect 158686 79716 158760 79744
rect 158352 79698 158404 79704
rect 158258 78976 158314 78985
rect 158258 78911 158314 78920
rect 158272 78878 158300 78911
rect 158260 78872 158312 78878
rect 158260 78814 158312 78820
rect 158364 78713 158392 79698
rect 158536 79620 158588 79626
rect 158536 79562 158588 79568
rect 158628 79620 158680 79626
rect 158628 79562 158680 79568
rect 158444 79552 158496 79558
rect 158444 79494 158496 79500
rect 158350 78704 158406 78713
rect 158350 78639 158406 78648
rect 158456 77518 158484 79494
rect 158444 77512 158496 77518
rect 158444 77454 158496 77460
rect 158260 76900 158312 76906
rect 158260 76842 158312 76848
rect 158168 76764 158220 76770
rect 158168 76706 158220 76712
rect 158272 73846 158300 76842
rect 158260 73840 158312 73846
rect 158260 73782 158312 73788
rect 158548 73778 158576 79562
rect 158640 77353 158668 79562
rect 158732 77450 158760 79716
rect 158962 79744 158990 80036
rect 158812 79698 158864 79704
rect 158916 79716 158990 79744
rect 158824 78130 158852 79698
rect 158812 78124 158864 78130
rect 158812 78066 158864 78072
rect 158720 77444 158772 77450
rect 158720 77386 158772 77392
rect 158626 77344 158682 77353
rect 158916 77314 158944 79716
rect 159054 79676 159082 80036
rect 159146 79898 159174 80036
rect 159134 79892 159186 79898
rect 159134 79834 159186 79840
rect 159238 79744 159266 80036
rect 159330 79937 159358 80036
rect 159316 79928 159372 79937
rect 159316 79863 159372 79872
rect 159008 79648 159082 79676
rect 159192 79716 159266 79744
rect 158626 77279 158682 77288
rect 158904 77308 158956 77314
rect 158904 77250 158956 77256
rect 158628 77240 158680 77246
rect 159008 77194 159036 79648
rect 159192 79218 159220 79716
rect 159422 79676 159450 80036
rect 159514 79898 159542 80036
rect 159502 79892 159554 79898
rect 159502 79834 159554 79840
rect 159606 79778 159634 80036
rect 159698 79966 159726 80036
rect 159686 79960 159738 79966
rect 159686 79902 159738 79908
rect 159790 79812 159818 80036
rect 159744 79784 159818 79812
rect 159606 79750 159680 79778
rect 159548 79688 159600 79694
rect 159422 79648 159496 79676
rect 159272 79620 159324 79626
rect 159272 79562 159324 79568
rect 159180 79212 159232 79218
rect 159180 79154 159232 79160
rect 159088 77308 159140 77314
rect 159088 77250 159140 77256
rect 158628 77182 158680 77188
rect 158536 73772 158588 73778
rect 158536 73714 158588 73720
rect 158640 71194 158668 77182
rect 158732 77166 159036 77194
rect 158628 71188 158680 71194
rect 158628 71130 158680 71136
rect 157996 70366 158392 70394
rect 157800 55888 157852 55894
rect 157800 55830 157852 55836
rect 157708 33856 157760 33862
rect 157708 33798 157760 33804
rect 158364 31210 158392 70366
rect 158352 31204 158404 31210
rect 158352 31146 158404 31152
rect 157616 13456 157668 13462
rect 157616 13398 157668 13404
rect 157524 13388 157576 13394
rect 157524 13330 157576 13336
rect 158732 11966 158760 77166
rect 158812 76628 158864 76634
rect 158812 76570 158864 76576
rect 158824 14958 158852 76570
rect 158904 76560 158956 76566
rect 158904 76502 158956 76508
rect 158916 26994 158944 76502
rect 158996 76492 159048 76498
rect 158996 76434 159048 76440
rect 159008 28354 159036 76434
rect 159100 28422 159128 77250
rect 159180 76696 159232 76702
rect 159180 76638 159232 76644
rect 159192 31142 159220 76638
rect 159284 67114 159312 79562
rect 159468 77840 159496 79648
rect 159548 79630 159600 79636
rect 159376 77812 159496 77840
rect 159376 76634 159404 77812
rect 159560 77738 159588 79630
rect 159468 77710 159588 77738
rect 159364 76628 159416 76634
rect 159364 76570 159416 76576
rect 159468 76566 159496 77710
rect 159652 77602 159680 79750
rect 159560 77574 159680 77602
rect 159456 76560 159508 76566
rect 159456 76502 159508 76508
rect 159560 76498 159588 77574
rect 159640 77444 159692 77450
rect 159640 77386 159692 77392
rect 159548 76492 159600 76498
rect 159548 76434 159600 76440
rect 159652 71126 159680 77386
rect 159744 76702 159772 79784
rect 159882 79744 159910 80036
rect 159974 79903 160002 80036
rect 159960 79894 160016 79903
rect 159960 79829 160016 79838
rect 160066 79778 160094 80036
rect 160158 79898 160186 80036
rect 160250 79937 160278 80036
rect 160236 79928 160292 79937
rect 160146 79892 160198 79898
rect 160236 79863 160292 79872
rect 160146 79834 160198 79840
rect 160342 79778 160370 80036
rect 160434 79898 160462 80036
rect 160422 79892 160474 79898
rect 160422 79834 160474 79840
rect 159836 79716 159910 79744
rect 160020 79750 160094 79778
rect 160296 79750 160370 79778
rect 159836 77654 159864 79716
rect 159914 79520 159970 79529
rect 159914 79455 159970 79464
rect 159928 79014 159956 79455
rect 159916 79008 159968 79014
rect 159916 78950 159968 78956
rect 159824 77648 159876 77654
rect 159824 77590 159876 77596
rect 160020 77353 160048 79750
rect 160296 79744 160324 79750
rect 160526 79744 160554 80036
rect 160618 79778 160646 80036
rect 160710 79898 160738 80036
rect 160802 79966 160830 80036
rect 160790 79960 160842 79966
rect 160790 79902 160842 79908
rect 160894 79898 160922 80036
rect 160698 79892 160750 79898
rect 160698 79834 160750 79840
rect 160882 79892 160934 79898
rect 160882 79834 160934 79840
rect 160618 79750 160692 79778
rect 160204 79716 160324 79744
rect 160480 79716 160554 79744
rect 160006 77344 160062 77353
rect 160006 77279 160062 77288
rect 160100 76764 160152 76770
rect 160100 76706 160152 76712
rect 159732 76696 159784 76702
rect 159732 76638 159784 76644
rect 159824 73772 159876 73778
rect 159824 73714 159876 73720
rect 159836 72486 159864 73714
rect 159824 72480 159876 72486
rect 159824 72422 159876 72428
rect 159640 71120 159692 71126
rect 159640 71062 159692 71068
rect 159272 67108 159324 67114
rect 159272 67050 159324 67056
rect 159362 65512 159418 65521
rect 159362 65447 159418 65456
rect 159180 31136 159232 31142
rect 159180 31078 159232 31084
rect 159088 28416 159140 28422
rect 159088 28358 159140 28364
rect 158996 28348 159048 28354
rect 158996 28290 159048 28296
rect 158904 26988 158956 26994
rect 158904 26930 158956 26936
rect 158812 14952 158864 14958
rect 158812 14894 158864 14900
rect 158720 11960 158772 11966
rect 158720 11902 158772 11908
rect 157432 10532 157484 10538
rect 157432 10474 157484 10480
rect 157340 10464 157392 10470
rect 157340 10406 157392 10412
rect 156972 9444 157024 9450
rect 156972 9386 157024 9392
rect 157800 4956 157852 4962
rect 157800 4898 157852 4904
rect 156420 3596 156472 3602
rect 156420 3538 156472 3544
rect 156432 3330 156460 3538
rect 156420 3324 156472 3330
rect 156420 3266 156472 3272
rect 157812 480 157840 4898
rect 159376 3806 159404 65447
rect 160112 9246 160140 76706
rect 160204 9382 160232 79716
rect 160284 79620 160336 79626
rect 160284 79562 160336 79568
rect 160296 77450 160324 79562
rect 160376 79552 160428 79558
rect 160376 79494 160428 79500
rect 160284 77444 160336 77450
rect 160284 77386 160336 77392
rect 160388 77330 160416 79494
rect 160296 77302 160416 77330
rect 160192 9376 160244 9382
rect 160192 9318 160244 9324
rect 160296 9314 160324 77302
rect 160376 77240 160428 77246
rect 160376 77182 160428 77188
rect 160388 76770 160416 77182
rect 160376 76764 160428 76770
rect 160376 76706 160428 76712
rect 160480 76650 160508 79716
rect 160664 79558 160692 79750
rect 160744 79756 160796 79762
rect 160744 79698 160796 79704
rect 160836 79756 160888 79762
rect 160986 79744 161014 80036
rect 161078 79966 161106 80036
rect 161066 79960 161118 79966
rect 161170 79937 161198 80036
rect 161066 79902 161118 79908
rect 161156 79928 161212 79937
rect 161156 79863 161212 79872
rect 161262 79812 161290 80036
rect 161354 79966 161382 80036
rect 161446 79966 161474 80036
rect 161342 79960 161394 79966
rect 161342 79902 161394 79908
rect 161434 79960 161486 79966
rect 161538 79937 161566 80036
rect 161434 79902 161486 79908
rect 161524 79928 161580 79937
rect 161524 79863 161580 79872
rect 161216 79801 161290 79812
rect 160836 79698 160888 79704
rect 160940 79716 161014 79744
rect 161202 79792 161290 79801
rect 161258 79784 161290 79792
rect 161630 79778 161658 80036
rect 161722 79898 161750 80036
rect 161710 79892 161762 79898
rect 161710 79834 161762 79840
rect 161202 79727 161258 79736
rect 161480 79756 161532 79762
rect 160652 79552 160704 79558
rect 160652 79494 160704 79500
rect 160756 76770 160784 79698
rect 160848 77246 160876 79698
rect 160836 77240 160888 77246
rect 160836 77182 160888 77188
rect 160744 76764 160796 76770
rect 160744 76706 160796 76712
rect 160480 76622 160600 76650
rect 160468 76560 160520 76566
rect 160468 76502 160520 76508
rect 160376 76492 160428 76498
rect 160376 76434 160428 76440
rect 160388 11898 160416 76434
rect 160480 14890 160508 76502
rect 160572 16182 160600 76622
rect 160744 76628 160796 76634
rect 160744 76570 160796 76576
rect 160652 76492 160704 76498
rect 160652 76434 160704 76440
rect 160560 16176 160612 16182
rect 160560 16118 160612 16124
rect 160664 16114 160692 76434
rect 160756 51746 160784 76570
rect 160940 76566 160968 79716
rect 161630 79750 161704 79778
rect 161480 79698 161532 79704
rect 161492 79642 161520 79698
rect 161020 79620 161072 79626
rect 161020 79562 161072 79568
rect 161112 79620 161164 79626
rect 161112 79562 161164 79568
rect 161296 79620 161348 79626
rect 161296 79562 161348 79568
rect 161400 79614 161520 79642
rect 161572 79688 161624 79694
rect 161572 79630 161624 79636
rect 161032 76634 161060 79562
rect 161124 77704 161152 79562
rect 161204 79552 161256 79558
rect 161308 79529 161336 79562
rect 161204 79494 161256 79500
rect 161294 79520 161350 79529
rect 161216 78062 161244 79494
rect 161294 79455 161350 79464
rect 161296 79212 161348 79218
rect 161296 79154 161348 79160
rect 161204 78056 161256 78062
rect 161204 77998 161256 78004
rect 161124 77676 161244 77704
rect 161112 77580 161164 77586
rect 161112 77522 161164 77528
rect 161124 77246 161152 77522
rect 161112 77240 161164 77246
rect 161112 77182 161164 77188
rect 161020 76628 161072 76634
rect 161020 76570 161072 76576
rect 160928 76560 160980 76566
rect 160834 76528 160890 76537
rect 160928 76502 160980 76508
rect 161216 76498 161244 77676
rect 161308 76770 161336 79154
rect 161296 76764 161348 76770
rect 161296 76706 161348 76712
rect 161400 76537 161428 79614
rect 161480 79552 161532 79558
rect 161480 79494 161532 79500
rect 161386 76528 161442 76537
rect 160834 76463 160890 76472
rect 161204 76492 161256 76498
rect 160848 61470 160876 76463
rect 161386 76463 161442 76472
rect 161204 76434 161256 76440
rect 160836 61464 160888 61470
rect 160836 61406 160888 61412
rect 160744 51740 160796 51746
rect 160744 51682 160796 51688
rect 160652 16108 160704 16114
rect 160652 16050 160704 16056
rect 160468 14884 160520 14890
rect 160468 14826 160520 14832
rect 160376 11892 160428 11898
rect 160376 11834 160428 11840
rect 161492 11830 161520 79494
rect 161584 77897 161612 79630
rect 161676 78010 161704 79750
rect 161814 79744 161842 80036
rect 161906 79898 161934 80036
rect 161894 79892 161946 79898
rect 161894 79834 161946 79840
rect 161998 79744 162026 80036
rect 161768 79716 161842 79744
rect 161952 79716 162026 79744
rect 162090 79744 162118 80036
rect 162182 79937 162210 80036
rect 162168 79928 162224 79937
rect 162168 79863 162224 79872
rect 162274 79744 162302 80036
rect 162366 79898 162394 80036
rect 162354 79892 162406 79898
rect 162354 79834 162406 79840
rect 162458 79744 162486 80036
rect 162550 79966 162578 80036
rect 162642 79966 162670 80036
rect 162734 79971 162762 80036
rect 162538 79960 162590 79966
rect 162538 79902 162590 79908
rect 162630 79960 162682 79966
rect 162630 79902 162682 79908
rect 162720 79962 162776 79971
rect 162826 79966 162854 80036
rect 162720 79897 162776 79906
rect 162814 79960 162866 79966
rect 162814 79902 162866 79908
rect 162584 79824 162636 79830
rect 162584 79766 162636 79772
rect 162090 79716 162164 79744
rect 161768 78198 161796 79716
rect 161846 79656 161902 79665
rect 161846 79591 161902 79600
rect 161756 78192 161808 78198
rect 161756 78134 161808 78140
rect 161676 77982 161796 78010
rect 161664 77920 161716 77926
rect 161570 77888 161626 77897
rect 161664 77862 161716 77868
rect 161570 77823 161626 77832
rect 161572 76628 161624 76634
rect 161572 76570 161624 76576
rect 161584 13326 161612 76570
rect 161572 13320 161624 13326
rect 161572 13262 161624 13268
rect 161676 13258 161704 77862
rect 161768 14822 161796 77982
rect 161860 17406 161888 79591
rect 161952 76634 161980 79716
rect 162136 79558 162164 79716
rect 162228 79716 162302 79744
rect 162412 79716 162486 79744
rect 162124 79552 162176 79558
rect 162124 79494 162176 79500
rect 162032 79212 162084 79218
rect 162032 79154 162084 79160
rect 162044 78305 162072 79154
rect 162228 79014 162256 79716
rect 162308 79620 162360 79626
rect 162308 79562 162360 79568
rect 162124 79008 162176 79014
rect 162124 78950 162176 78956
rect 162216 79008 162268 79014
rect 162216 78950 162268 78956
rect 162136 78690 162164 78950
rect 162136 78662 162256 78690
rect 162030 78296 162086 78305
rect 162030 78231 162086 78240
rect 162032 78192 162084 78198
rect 162032 78134 162084 78140
rect 161940 76628 161992 76634
rect 161940 76570 161992 76576
rect 161940 76492 161992 76498
rect 161940 76434 161992 76440
rect 161952 19038 161980 76434
rect 162044 32638 162072 78134
rect 162124 77852 162176 77858
rect 162124 77794 162176 77800
rect 162136 76634 162164 77794
rect 162124 76628 162176 76634
rect 162124 76570 162176 76576
rect 162228 76430 162256 78662
rect 162320 76498 162348 79562
rect 162412 79218 162440 79716
rect 162492 79620 162544 79626
rect 162492 79562 162544 79568
rect 162400 79212 162452 79218
rect 162400 79154 162452 79160
rect 162400 79008 162452 79014
rect 162400 78950 162452 78956
rect 162412 77926 162440 78950
rect 162400 77920 162452 77926
rect 162400 77862 162452 77868
rect 162400 77784 162452 77790
rect 162400 77726 162452 77732
rect 162308 76492 162360 76498
rect 162308 76434 162360 76440
rect 162216 76424 162268 76430
rect 162216 76366 162268 76372
rect 162032 32632 162084 32638
rect 162032 32574 162084 32580
rect 161940 19032 161992 19038
rect 161940 18974 161992 18980
rect 161848 17400 161900 17406
rect 161848 17342 161900 17348
rect 162412 15094 162440 77726
rect 162504 76129 162532 79562
rect 162596 78470 162624 79766
rect 162918 79744 162946 80036
rect 163010 79966 163038 80036
rect 162998 79960 163050 79966
rect 162998 79902 163050 79908
rect 163102 79898 163130 80036
rect 163194 79898 163222 80036
rect 163090 79892 163142 79898
rect 163090 79834 163142 79840
rect 163182 79892 163234 79898
rect 163182 79834 163234 79840
rect 163286 79778 163314 80036
rect 163378 79898 163406 80036
rect 163366 79892 163418 79898
rect 163366 79834 163418 79840
rect 163286 79750 163360 79778
rect 162918 79716 162992 79744
rect 162676 79620 162728 79626
rect 162676 79562 162728 79568
rect 162860 79620 162912 79626
rect 162860 79562 162912 79568
rect 162584 78464 162636 78470
rect 162584 78406 162636 78412
rect 162688 76265 162716 79562
rect 162768 79280 162820 79286
rect 162768 79222 162820 79228
rect 162780 79014 162808 79222
rect 162768 79008 162820 79014
rect 162768 78950 162820 78956
rect 162674 76256 162730 76265
rect 162674 76191 162730 76200
rect 162490 76120 162546 76129
rect 162490 76055 162546 76064
rect 162400 15088 162452 15094
rect 162400 15030 162452 15036
rect 161756 14816 161808 14822
rect 161756 14758 161808 14764
rect 162872 14754 162900 79562
rect 162964 76412 162992 79716
rect 163044 79688 163096 79694
rect 163228 79688 163280 79694
rect 163096 79648 163176 79676
rect 163044 79630 163096 79636
rect 163148 76616 163176 79648
rect 163228 79630 163280 79636
rect 163240 78441 163268 79630
rect 163226 78432 163282 78441
rect 163226 78367 163282 78376
rect 163148 76588 163268 76616
rect 162964 76384 163176 76412
rect 162952 75336 163004 75342
rect 162952 75278 163004 75284
rect 162860 14748 162912 14754
rect 162860 14690 162912 14696
rect 162964 14686 162992 75278
rect 163044 75200 163096 75206
rect 163044 75142 163096 75148
rect 163056 18970 163084 75142
rect 163148 21690 163176 76384
rect 163240 29714 163268 76588
rect 163332 76226 163360 79750
rect 163470 79608 163498 80036
rect 163424 79580 163498 79608
rect 163562 79608 163590 80036
rect 163654 79830 163682 80036
rect 163642 79824 163694 79830
rect 163746 79801 163774 80036
rect 163838 79812 163866 80036
rect 163930 79966 163958 80036
rect 163918 79960 163970 79966
rect 163918 79902 163970 79908
rect 164022 79812 164050 80036
rect 164114 79898 164142 80036
rect 164206 79903 164234 80036
rect 164102 79892 164154 79898
rect 164102 79834 164154 79840
rect 164192 79894 164248 79903
rect 164192 79829 164248 79838
rect 163642 79766 163694 79772
rect 163732 79792 163788 79801
rect 163838 79784 163912 79812
rect 163732 79727 163788 79736
rect 163780 79688 163832 79694
rect 163780 79630 163832 79636
rect 163688 79620 163740 79626
rect 163562 79580 163636 79608
rect 163320 76220 163372 76226
rect 163320 76162 163372 76168
rect 163320 75132 163372 75138
rect 163320 75074 163372 75080
rect 163332 32570 163360 75074
rect 163424 35222 163452 79580
rect 163504 76220 163556 76226
rect 163504 76162 163556 76168
rect 163516 64326 163544 76162
rect 163504 64320 163556 64326
rect 163504 64262 163556 64268
rect 163608 64258 163636 79580
rect 163688 79562 163740 79568
rect 163700 75138 163728 79562
rect 163688 75132 163740 75138
rect 163688 75074 163740 75080
rect 163792 69902 163820 79630
rect 163884 75206 163912 79784
rect 163976 79784 164050 79812
rect 163976 78713 164004 79784
rect 164298 79744 164326 80036
rect 164252 79716 164326 79744
rect 164056 79688 164108 79694
rect 164056 79630 164108 79636
rect 164068 78985 164096 79630
rect 164148 79620 164200 79626
rect 164148 79562 164200 79568
rect 164054 78976 164110 78985
rect 164054 78911 164110 78920
rect 163962 78704 164018 78713
rect 163962 78639 164018 78648
rect 164160 75342 164188 79562
rect 164252 77790 164280 79716
rect 164390 79676 164418 80036
rect 164482 79778 164510 80036
rect 164574 79898 164602 80036
rect 164666 79966 164694 80036
rect 164654 79960 164706 79966
rect 164654 79902 164706 79908
rect 164758 79898 164786 80036
rect 164562 79892 164614 79898
rect 164562 79834 164614 79840
rect 164746 79892 164798 79898
rect 164746 79834 164798 79840
rect 164482 79750 164556 79778
rect 164390 79648 164464 79676
rect 164332 79552 164384 79558
rect 164330 79520 164332 79529
rect 164384 79520 164386 79529
rect 164330 79455 164386 79464
rect 164332 79416 164384 79422
rect 164332 79358 164384 79364
rect 164344 79150 164372 79358
rect 164332 79144 164384 79150
rect 164332 79086 164384 79092
rect 164332 78192 164384 78198
rect 164332 78134 164384 78140
rect 164240 77784 164292 77790
rect 164240 77726 164292 77732
rect 164240 77376 164292 77382
rect 164240 77318 164292 77324
rect 164148 75336 164200 75342
rect 164148 75278 164200 75284
rect 163872 75200 163924 75206
rect 163872 75142 163924 75148
rect 163780 69896 163832 69902
rect 163780 69838 163832 69844
rect 163596 64252 163648 64258
rect 163596 64194 163648 64200
rect 163412 35216 163464 35222
rect 163412 35158 163464 35164
rect 163320 32564 163372 32570
rect 163320 32506 163372 32512
rect 163228 29708 163280 29714
rect 163228 29650 163280 29656
rect 163136 21684 163188 21690
rect 163136 21626 163188 21632
rect 163044 18964 163096 18970
rect 163044 18906 163096 18912
rect 162952 14680 163004 14686
rect 162952 14622 163004 14628
rect 161664 13252 161716 13258
rect 161664 13194 161716 13200
rect 161480 11824 161532 11830
rect 161480 11766 161532 11772
rect 160284 9308 160336 9314
rect 160284 9250 160336 9256
rect 160100 9240 160152 9246
rect 160100 9182 160152 9188
rect 164252 5098 164280 77318
rect 164344 9178 164372 78134
rect 164436 75410 164464 79648
rect 164424 75404 164476 75410
rect 164424 75346 164476 75352
rect 164424 75268 164476 75274
rect 164424 75210 164476 75216
rect 164436 18902 164464 75210
rect 164528 32502 164556 79750
rect 164850 79676 164878 80036
rect 164942 79744 164970 80036
rect 165034 79937 165062 80036
rect 165020 79928 165076 79937
rect 165020 79863 165076 79872
rect 165126 79744 165154 80036
rect 165218 79966 165246 80036
rect 165206 79960 165258 79966
rect 165206 79902 165258 79908
rect 165310 79898 165338 80036
rect 165298 79892 165350 79898
rect 165298 79834 165350 79840
rect 165402 79830 165430 80036
rect 165390 79824 165442 79830
rect 165494 79812 165522 80036
rect 165586 79937 165614 80036
rect 165678 79966 165706 80036
rect 165770 79966 165798 80036
rect 165666 79960 165718 79966
rect 165572 79928 165628 79937
rect 165666 79902 165718 79908
rect 165758 79960 165810 79966
rect 165758 79902 165810 79908
rect 165862 79898 165890 80036
rect 165954 79971 165982 80036
rect 165940 79962 165996 79971
rect 165572 79863 165628 79872
rect 165850 79892 165902 79898
rect 165940 79897 165996 79906
rect 166046 79898 166074 80036
rect 165850 79834 165902 79840
rect 166034 79892 166086 79898
rect 166034 79834 166086 79840
rect 165494 79801 165568 79812
rect 165494 79792 165582 79801
rect 165494 79784 165526 79792
rect 165390 79766 165442 79772
rect 165252 79756 165304 79762
rect 164942 79716 165062 79744
rect 165126 79716 165200 79744
rect 165034 79676 165062 79716
rect 164850 79648 164924 79676
rect 165034 79648 165108 79676
rect 164608 79620 164660 79626
rect 164608 79562 164660 79568
rect 164620 78198 164648 79562
rect 164792 79552 164844 79558
rect 164792 79494 164844 79500
rect 164608 78192 164660 78198
rect 164608 78134 164660 78140
rect 164608 77988 164660 77994
rect 164608 77930 164660 77936
rect 164516 32496 164568 32502
rect 164516 32438 164568 32444
rect 164620 32434 164648 77930
rect 164698 76256 164754 76265
rect 164698 76191 164754 76200
rect 164712 33794 164740 76191
rect 164804 65754 164832 79494
rect 164896 78198 164924 79648
rect 164976 79552 165028 79558
rect 164976 79494 165028 79500
rect 164884 78192 164936 78198
rect 164884 78134 164936 78140
rect 164884 78056 164936 78062
rect 164884 77998 164936 78004
rect 164896 75562 164924 77998
rect 164988 77994 165016 79494
rect 164976 77988 165028 77994
rect 164976 77930 165028 77936
rect 164896 75534 165016 75562
rect 164884 75404 164936 75410
rect 164884 75346 164936 75352
rect 164896 68474 164924 75346
rect 164988 73154 165016 75534
rect 165080 75274 165108 79648
rect 165172 77382 165200 79716
rect 166138 79778 166166 80036
rect 166230 79830 166258 80036
rect 166322 79898 166350 80036
rect 166414 79898 166442 80036
rect 166310 79892 166362 79898
rect 166310 79834 166362 79840
rect 166402 79892 166454 79898
rect 166402 79834 166454 79840
rect 165526 79727 165582 79736
rect 165896 79756 165948 79762
rect 165252 79698 165304 79704
rect 165896 79698 165948 79704
rect 165988 79756 166040 79762
rect 165988 79698 166040 79704
rect 166092 79750 166166 79778
rect 166218 79824 166270 79830
rect 166218 79766 166270 79772
rect 165264 78033 165292 79698
rect 165804 79688 165856 79694
rect 165804 79630 165856 79636
rect 165436 79620 165488 79626
rect 165436 79562 165488 79568
rect 165528 79620 165580 79626
rect 165528 79562 165580 79568
rect 165712 79620 165764 79626
rect 165712 79562 165764 79568
rect 165344 79552 165396 79558
rect 165344 79494 165396 79500
rect 165250 78024 165306 78033
rect 165250 77959 165306 77968
rect 165160 77376 165212 77382
rect 165160 77318 165212 77324
rect 165356 76702 165384 79494
rect 165448 78169 165476 79562
rect 165434 78160 165490 78169
rect 165434 78095 165490 78104
rect 165540 78033 165568 79562
rect 165620 79416 165672 79422
rect 165620 79358 165672 79364
rect 165632 79286 165660 79358
rect 165620 79280 165672 79286
rect 165620 79222 165672 79228
rect 165618 78976 165674 78985
rect 165618 78911 165674 78920
rect 165632 78810 165660 78911
rect 165620 78804 165672 78810
rect 165620 78746 165672 78752
rect 165526 78024 165582 78033
rect 165526 77959 165582 77968
rect 165618 77616 165674 77625
rect 165618 77551 165674 77560
rect 165436 77512 165488 77518
rect 165436 77454 165488 77460
rect 165344 76696 165396 76702
rect 165344 76638 165396 76644
rect 165068 75268 165120 75274
rect 165068 75210 165120 75216
rect 164988 73126 165292 73154
rect 164884 68468 164936 68474
rect 164884 68410 164936 68416
rect 164792 65748 164844 65754
rect 164792 65690 164844 65696
rect 165264 64394 165292 73126
rect 165448 72554 165476 77454
rect 165632 77382 165660 77551
rect 165620 77376 165672 77382
rect 165620 77318 165672 77324
rect 165620 76900 165672 76906
rect 165620 76842 165672 76848
rect 165436 72548 165488 72554
rect 165436 72490 165488 72496
rect 165252 64388 165304 64394
rect 165252 64330 165304 64336
rect 164700 33788 164752 33794
rect 164700 33730 164752 33736
rect 164608 32428 164660 32434
rect 164608 32370 164660 32376
rect 164424 18896 164476 18902
rect 164424 18838 164476 18844
rect 164332 9172 164384 9178
rect 164332 9114 164384 9120
rect 165632 6254 165660 76842
rect 165724 6322 165752 79562
rect 165816 77858 165844 79630
rect 165804 77852 165856 77858
rect 165804 77794 165856 77800
rect 165804 77716 165856 77722
rect 165804 77658 165856 77664
rect 165816 7750 165844 77658
rect 165908 77602 165936 79698
rect 166000 77722 166028 79698
rect 165988 77716 166040 77722
rect 165988 77658 166040 77664
rect 165908 77574 166028 77602
rect 165896 76696 165948 76702
rect 165896 76638 165948 76644
rect 165908 9042 165936 76638
rect 166000 9110 166028 77574
rect 166092 10334 166120 79750
rect 166506 79744 166534 80036
rect 166598 79801 166626 80036
rect 166690 79937 166718 80036
rect 166676 79928 166732 79937
rect 166782 79898 166810 80036
rect 166874 79966 166902 80036
rect 166862 79960 166914 79966
rect 166862 79902 166914 79908
rect 166676 79863 166732 79872
rect 166770 79892 166822 79898
rect 166770 79834 166822 79840
rect 166966 79812 166994 80036
rect 166460 79716 166534 79744
rect 166584 79792 166640 79801
rect 166920 79784 166994 79812
rect 166816 79756 166868 79762
rect 166584 79727 166640 79736
rect 166736 79716 166816 79744
rect 166172 79688 166224 79694
rect 166354 79656 166410 79665
rect 166224 79636 166304 79642
rect 166172 79630 166304 79636
rect 166184 79614 166304 79630
rect 166172 79552 166224 79558
rect 166172 79494 166224 79500
rect 166184 76906 166212 79494
rect 166172 76900 166224 76906
rect 166172 76842 166224 76848
rect 166172 76560 166224 76566
rect 166172 76502 166224 76508
rect 166184 20058 166212 76502
rect 166276 68406 166304 79614
rect 166354 79591 166410 79600
rect 166368 77518 166396 79591
rect 166460 78033 166488 79716
rect 166538 79656 166594 79665
rect 166538 79591 166594 79600
rect 166446 78024 166502 78033
rect 166446 77959 166502 77968
rect 166448 77852 166500 77858
rect 166448 77794 166500 77800
rect 166356 77512 166408 77518
rect 166356 77454 166408 77460
rect 166460 70394 166488 77794
rect 166552 76566 166580 79591
rect 166632 79552 166684 79558
rect 166632 79494 166684 79500
rect 166644 77353 166672 79494
rect 166736 77489 166764 79716
rect 166816 79698 166868 79704
rect 166816 79620 166868 79626
rect 166816 79562 166868 79568
rect 166828 78538 166856 79562
rect 166920 79370 166948 79784
rect 167058 79744 167086 80036
rect 167150 79898 167178 80036
rect 167138 79892 167190 79898
rect 167138 79834 167190 79840
rect 167242 79744 167270 80036
rect 167334 79937 167362 80036
rect 167426 79966 167454 80036
rect 167518 79966 167546 80036
rect 167414 79960 167466 79966
rect 167320 79928 167376 79937
rect 167414 79902 167466 79908
rect 167506 79960 167558 79966
rect 167506 79902 167558 79908
rect 167320 79863 167376 79872
rect 167368 79824 167420 79830
rect 167610 79812 167638 80036
rect 167368 79766 167420 79772
rect 167564 79784 167638 79812
rect 167058 79716 167132 79744
rect 166920 79342 167040 79370
rect 166908 79212 166960 79218
rect 166908 79154 166960 79160
rect 166816 78532 166868 78538
rect 166816 78474 166868 78480
rect 166920 78266 166948 79154
rect 166908 78260 166960 78266
rect 166908 78202 166960 78208
rect 166908 78124 166960 78130
rect 166908 78066 166960 78072
rect 166722 77480 166778 77489
rect 166722 77415 166778 77424
rect 166630 77344 166686 77353
rect 166630 77279 166686 77288
rect 166540 76560 166592 76566
rect 166540 76502 166592 76508
rect 166920 70394 166948 78066
rect 167012 77625 167040 79342
rect 167104 78266 167132 79716
rect 167196 79716 167270 79744
rect 167092 78260 167144 78266
rect 167092 78202 167144 78208
rect 166998 77616 167054 77625
rect 166998 77551 167054 77560
rect 167196 75914 167224 79716
rect 167276 79620 167328 79626
rect 167276 79562 167328 79568
rect 166368 70366 166488 70394
rect 166644 70366 166948 70394
rect 167012 75886 167224 75914
rect 166368 69834 166396 70366
rect 166356 69828 166408 69834
rect 166356 69770 166408 69776
rect 166264 68400 166316 68406
rect 166264 68342 166316 68348
rect 166644 62898 166672 70366
rect 166632 62892 166684 62898
rect 166632 62834 166684 62840
rect 166172 20052 166224 20058
rect 166172 19994 166224 20000
rect 166080 10328 166132 10334
rect 166080 10270 166132 10276
rect 165988 9104 166040 9110
rect 165988 9046 166040 9052
rect 165896 9036 165948 9042
rect 165896 8978 165948 8984
rect 165804 7744 165856 7750
rect 165804 7686 165856 7692
rect 167012 7614 167040 75886
rect 167184 75336 167236 75342
rect 167184 75278 167236 75284
rect 167092 75200 167144 75206
rect 167092 75142 167144 75148
rect 167104 16046 167132 75142
rect 167092 16040 167144 16046
rect 167092 15982 167144 15988
rect 167196 15978 167224 75278
rect 167288 20126 167316 79562
rect 167380 77858 167408 79766
rect 167460 79688 167512 79694
rect 167460 79630 167512 79636
rect 167368 77852 167420 77858
rect 167368 77794 167420 77800
rect 167368 75132 167420 75138
rect 167368 75074 167420 75080
rect 167380 21622 167408 75074
rect 167472 25634 167500 79630
rect 167564 78062 167592 79784
rect 167702 79744 167730 80036
rect 167656 79716 167730 79744
rect 167794 79744 167822 80036
rect 167886 79898 167914 80036
rect 167874 79892 167926 79898
rect 167874 79834 167926 79840
rect 167978 79830 168006 80036
rect 168070 79937 168098 80036
rect 168056 79928 168112 79937
rect 168162 79898 168190 80036
rect 168254 79937 168282 80036
rect 168346 79966 168374 80036
rect 168334 79960 168386 79966
rect 168240 79928 168296 79937
rect 168056 79863 168112 79872
rect 168150 79892 168202 79898
rect 168334 79902 168386 79908
rect 168438 79898 168466 80036
rect 168240 79863 168296 79872
rect 168426 79892 168478 79898
rect 168150 79834 168202 79840
rect 168426 79834 168478 79840
rect 168530 79830 168558 80036
rect 168622 79898 168650 80036
rect 168610 79892 168662 79898
rect 168610 79834 168662 79840
rect 168714 79830 168742 80036
rect 168806 79937 168834 80036
rect 168792 79928 168848 79937
rect 168792 79863 168848 79872
rect 167966 79824 168018 79830
rect 167966 79766 168018 79772
rect 168518 79824 168570 79830
rect 168518 79766 168570 79772
rect 168702 79824 168754 79830
rect 168898 79812 168926 80036
rect 168990 79971 169018 80036
rect 168976 79962 169032 79971
rect 168976 79897 169032 79906
rect 169082 79812 169110 80036
rect 169174 79966 169202 80036
rect 169162 79960 169214 79966
rect 169162 79902 169214 79908
rect 169266 79898 169294 80036
rect 169358 79966 169386 80036
rect 169450 79966 169478 80036
rect 169346 79960 169398 79966
rect 169346 79902 169398 79908
rect 169438 79960 169490 79966
rect 169438 79902 169490 79908
rect 169542 79903 169570 80036
rect 169254 79892 169306 79898
rect 169254 79834 169306 79840
rect 169528 79894 169584 79903
rect 169634 79898 169662 80036
rect 169528 79829 169584 79838
rect 169622 79892 169674 79898
rect 169622 79834 169674 79840
rect 168852 79801 168926 79812
rect 168702 79766 168754 79772
rect 168838 79792 168926 79801
rect 168196 79756 168248 79762
rect 167794 79716 167868 79744
rect 167552 78056 167604 78062
rect 167552 77998 167604 78004
rect 167552 77852 167604 77858
rect 167552 77794 167604 77800
rect 167564 67046 167592 77794
rect 167656 75138 167684 79716
rect 167736 79484 167788 79490
rect 167736 79426 167788 79432
rect 167748 79286 167776 79426
rect 167736 79280 167788 79286
rect 167736 79222 167788 79228
rect 167736 77580 167788 77586
rect 167736 77522 167788 77528
rect 167644 75132 167696 75138
rect 167644 75074 167696 75080
rect 167748 70394 167776 77522
rect 167840 75206 167868 79716
rect 168894 79784 168926 79792
rect 169036 79784 169110 79812
rect 168838 79727 168894 79736
rect 168196 79698 168248 79704
rect 167920 79620 167972 79626
rect 167920 79562 167972 79568
rect 168104 79620 168156 79626
rect 168104 79562 168156 79568
rect 167932 75342 167960 79562
rect 168116 78606 168144 79562
rect 168104 78600 168156 78606
rect 168104 78542 168156 78548
rect 168010 77888 168066 77897
rect 168010 77823 168066 77832
rect 168024 77586 168052 77823
rect 168012 77580 168064 77586
rect 168012 77522 168064 77528
rect 168012 77444 168064 77450
rect 168012 77386 168064 77392
rect 167920 75336 167972 75342
rect 167920 75278 167972 75284
rect 167828 75200 167880 75206
rect 167828 75142 167880 75148
rect 168024 70394 168052 77386
rect 168102 77344 168158 77353
rect 168102 77279 168158 77288
rect 168116 74254 168144 77279
rect 168208 75313 168236 79698
rect 168288 79688 168340 79694
rect 168932 79688 168984 79694
rect 168288 79630 168340 79636
rect 168654 79656 168710 79665
rect 168300 79529 168328 79630
rect 168564 79620 168616 79626
rect 168932 79630 168984 79636
rect 168654 79591 168710 79600
rect 168564 79562 168616 79568
rect 168380 79552 168432 79558
rect 168286 79520 168342 79529
rect 168380 79494 168432 79500
rect 168286 79455 168342 79464
rect 168288 79416 168340 79422
rect 168288 79358 168340 79364
rect 168300 79150 168328 79358
rect 168288 79144 168340 79150
rect 168288 79086 168340 79092
rect 168288 78736 168340 78742
rect 168288 78678 168340 78684
rect 168300 77654 168328 78678
rect 168288 77648 168340 77654
rect 168288 77590 168340 77596
rect 168392 76566 168420 79494
rect 168576 79370 168604 79562
rect 168484 79342 168604 79370
rect 168380 76560 168432 76566
rect 168380 76502 168432 76508
rect 168380 76356 168432 76362
rect 168380 76298 168432 76304
rect 168194 75304 168250 75313
rect 168194 75239 168250 75248
rect 168104 74248 168156 74254
rect 168104 74190 168156 74196
rect 167748 70366 167960 70394
rect 168024 70366 168236 70394
rect 167552 67040 167604 67046
rect 167552 66982 167604 66988
rect 167932 35426 167960 70366
rect 168208 64874 168236 70366
rect 168024 64846 168236 64874
rect 167920 35420 167972 35426
rect 167920 35362 167972 35368
rect 168024 27062 168052 64846
rect 168012 27056 168064 27062
rect 168012 26998 168064 27004
rect 167460 25628 167512 25634
rect 167460 25570 167512 25576
rect 167368 21616 167420 21622
rect 167368 21558 167420 21564
rect 167276 20120 167328 20126
rect 167276 20062 167328 20068
rect 167184 15972 167236 15978
rect 167184 15914 167236 15920
rect 168392 11762 168420 76298
rect 168484 13122 168512 79342
rect 168564 79280 168616 79286
rect 168564 79222 168616 79228
rect 168576 79014 168604 79222
rect 168564 79008 168616 79014
rect 168564 78950 168616 78956
rect 168668 78962 168696 79591
rect 168838 79520 168894 79529
rect 168838 79455 168894 79464
rect 168668 78934 168788 78962
rect 168562 78704 168618 78713
rect 168562 78639 168618 78648
rect 168576 17338 168604 78639
rect 168760 77994 168788 78934
rect 168748 77988 168800 77994
rect 168748 77930 168800 77936
rect 168852 76362 168880 79455
rect 168840 76356 168892 76362
rect 168840 76298 168892 76304
rect 168656 76152 168708 76158
rect 168656 76094 168708 76100
rect 168668 21554 168696 76094
rect 168748 75336 168800 75342
rect 168748 75278 168800 75284
rect 168656 21548 168708 21554
rect 168656 21490 168708 21496
rect 168760 21486 168788 75278
rect 168840 75268 168892 75274
rect 168840 75210 168892 75216
rect 168852 31074 168880 75210
rect 168944 62830 168972 79630
rect 169036 78130 169064 79784
rect 169208 79756 169260 79762
rect 169208 79698 169260 79704
rect 169300 79756 169352 79762
rect 169300 79698 169352 79704
rect 169484 79756 169536 79762
rect 169726 79744 169754 80036
rect 169484 79698 169536 79704
rect 169680 79716 169754 79744
rect 169818 79744 169846 80036
rect 169910 79898 169938 80036
rect 170002 79898 170030 80036
rect 169898 79892 169950 79898
rect 169898 79834 169950 79840
rect 169990 79892 170042 79898
rect 169990 79834 170042 79840
rect 170094 79830 170122 80036
rect 170082 79824 170134 79830
rect 170186 79812 170214 80036
rect 170278 79971 170306 80036
rect 170264 79962 170320 79971
rect 170370 79966 170398 80036
rect 170264 79897 170320 79906
rect 170358 79960 170410 79966
rect 170358 79902 170410 79908
rect 170186 79784 170352 79812
rect 170082 79766 170134 79772
rect 169818 79716 169892 79744
rect 169116 79688 169168 79694
rect 169116 79630 169168 79636
rect 169024 78124 169076 78130
rect 169024 78066 169076 78072
rect 169128 76158 169156 79630
rect 169116 76152 169168 76158
rect 169116 76094 169168 76100
rect 169220 75274 169248 79698
rect 169208 75268 169260 75274
rect 169208 75210 169260 75216
rect 169312 70394 169340 79698
rect 169392 79552 169444 79558
rect 169390 79520 169392 79529
rect 169444 79520 169446 79529
rect 169390 79455 169446 79464
rect 169392 79144 169444 79150
rect 169392 79086 169444 79092
rect 169404 78674 169432 79086
rect 169392 78668 169444 78674
rect 169392 78610 169444 78616
rect 169496 75342 169524 79698
rect 169574 79656 169630 79665
rect 169574 79591 169630 79600
rect 169588 75818 169616 79591
rect 169680 79529 169708 79716
rect 169760 79620 169812 79626
rect 169760 79562 169812 79568
rect 169666 79520 169722 79529
rect 169666 79455 169722 79464
rect 169668 79076 169720 79082
rect 169668 79018 169720 79024
rect 169680 78810 169708 79018
rect 169668 78804 169720 78810
rect 169668 78746 169720 78752
rect 169668 78124 169720 78130
rect 169668 78066 169720 78072
rect 169680 77790 169708 78066
rect 169668 77784 169720 77790
rect 169668 77726 169720 77732
rect 169772 77654 169800 79562
rect 169760 77648 169812 77654
rect 169760 77590 169812 77596
rect 169576 75812 169628 75818
rect 169576 75754 169628 75760
rect 169484 75336 169536 75342
rect 169484 75278 169536 75284
rect 169036 70366 169340 70394
rect 169036 69766 169064 70366
rect 169024 69760 169076 69766
rect 169024 69702 169076 69708
rect 168932 62824 168984 62830
rect 168932 62766 168984 62772
rect 168840 31068 168892 31074
rect 168840 31010 168892 31016
rect 168748 21480 168800 21486
rect 168748 21422 168800 21428
rect 168564 17332 168616 17338
rect 168564 17274 168616 17280
rect 168472 13116 168524 13122
rect 168472 13058 168524 13064
rect 168380 11756 168432 11762
rect 168380 11698 168432 11704
rect 169864 7682 169892 79716
rect 170128 79688 170180 79694
rect 170180 79648 170260 79676
rect 170128 79630 170180 79636
rect 169944 79552 169996 79558
rect 169944 79494 169996 79500
rect 170128 79552 170180 79558
rect 170128 79494 170180 79500
rect 169956 77858 169984 79494
rect 170036 78396 170088 78402
rect 170036 78338 170088 78344
rect 169944 77852 169996 77858
rect 169944 77794 169996 77800
rect 169942 77752 169998 77761
rect 169942 77687 169998 77696
rect 169956 19990 169984 77687
rect 170048 22982 170076 78338
rect 170140 77976 170168 79494
rect 170232 78130 170260 79648
rect 170220 78124 170272 78130
rect 170220 78066 170272 78072
rect 170140 77948 170260 77976
rect 170128 77852 170180 77858
rect 170128 77794 170180 77800
rect 170140 60110 170168 77794
rect 170232 65686 170260 77948
rect 170324 75274 170352 79784
rect 170462 79778 170490 80036
rect 170554 79971 170582 80036
rect 170540 79962 170596 79971
rect 170646 79966 170674 80036
rect 170540 79897 170596 79906
rect 170634 79960 170686 79966
rect 170738 79937 170766 80036
rect 170830 79966 170858 80036
rect 170922 79971 170950 80036
rect 170818 79960 170870 79966
rect 170634 79902 170686 79908
rect 170724 79928 170780 79937
rect 170818 79902 170870 79908
rect 170908 79962 170964 79971
rect 171014 79966 171042 80036
rect 170908 79897 170964 79906
rect 171002 79960 171054 79966
rect 171106 79937 171134 80036
rect 171002 79902 171054 79908
rect 171092 79928 171148 79937
rect 170724 79863 170780 79872
rect 171092 79863 171148 79872
rect 170588 79824 170640 79830
rect 170462 79762 170536 79778
rect 171048 79824 171100 79830
rect 170640 79784 170812 79812
rect 170588 79766 170640 79772
rect 170462 79756 170548 79762
rect 170462 79750 170496 79756
rect 170496 79698 170548 79704
rect 170494 79656 170550 79665
rect 170416 79614 170494 79642
rect 170416 78402 170444 79614
rect 170494 79591 170550 79600
rect 170588 79620 170640 79626
rect 170588 79562 170640 79568
rect 170496 79552 170548 79558
rect 170496 79494 170548 79500
rect 170404 78396 170456 78402
rect 170404 78338 170456 78344
rect 170508 78044 170536 79494
rect 170416 78016 170536 78044
rect 170312 75268 170364 75274
rect 170312 75210 170364 75216
rect 170416 70394 170444 78016
rect 170600 77976 170628 79562
rect 170680 79552 170732 79558
rect 170680 79494 170732 79500
rect 170692 78713 170720 79494
rect 170678 78704 170734 78713
rect 170678 78639 170734 78648
rect 170680 78124 170732 78130
rect 170680 78066 170732 78072
rect 170508 77948 170628 77976
rect 170508 75478 170536 77948
rect 170588 77852 170640 77858
rect 170588 77794 170640 77800
rect 170496 75472 170548 75478
rect 170496 75414 170548 75420
rect 170324 70366 170444 70394
rect 170324 66978 170352 70366
rect 170600 68338 170628 77794
rect 170692 75750 170720 78066
rect 170784 77625 170812 79784
rect 171048 79766 171100 79772
rect 170956 79688 171008 79694
rect 170862 79656 170918 79665
rect 170956 79630 171008 79636
rect 170862 79591 170918 79600
rect 170876 77858 170904 79591
rect 170968 79218 170996 79630
rect 171060 79529 171088 79766
rect 171198 79744 171226 80036
rect 171152 79716 171226 79744
rect 171290 79744 171318 80036
rect 171382 79966 171410 80036
rect 171370 79960 171422 79966
rect 171370 79902 171422 79908
rect 171474 79812 171502 80036
rect 171428 79784 171502 79812
rect 171290 79716 171364 79744
rect 171046 79520 171102 79529
rect 171046 79455 171102 79464
rect 170956 79212 171008 79218
rect 170956 79154 171008 79160
rect 171152 79098 171180 79716
rect 171336 79665 171364 79716
rect 171322 79656 171378 79665
rect 171322 79591 171378 79600
rect 171428 79506 171456 79784
rect 171566 79744 171594 80036
rect 171658 79801 171686 80036
rect 171750 79937 171778 80036
rect 171736 79928 171792 79937
rect 171842 79898 171870 80036
rect 171736 79863 171792 79872
rect 171830 79892 171882 79898
rect 171830 79834 171882 79840
rect 170968 79070 171180 79098
rect 171244 79478 171456 79506
rect 171520 79716 171594 79744
rect 171644 79792 171700 79801
rect 171644 79727 171700 79736
rect 171784 79756 171836 79762
rect 170968 78538 170996 79070
rect 171140 79008 171192 79014
rect 171140 78950 171192 78956
rect 171048 78940 171100 78946
rect 171048 78882 171100 78888
rect 170956 78532 171008 78538
rect 170956 78474 171008 78480
rect 170954 78296 171010 78305
rect 170954 78231 171010 78240
rect 170968 77897 170996 78231
rect 170954 77888 171010 77897
rect 170864 77852 170916 77858
rect 171060 77858 171088 78882
rect 170954 77823 171010 77832
rect 171048 77852 171100 77858
rect 170864 77794 170916 77800
rect 171048 77794 171100 77800
rect 170770 77616 170826 77625
rect 170770 77551 170826 77560
rect 171152 77194 171180 78950
rect 171060 77166 171180 77194
rect 171060 76906 171088 77166
rect 171140 77036 171192 77042
rect 171140 76978 171192 76984
rect 171048 76900 171100 76906
rect 171048 76842 171100 76848
rect 171152 76634 171180 76978
rect 171140 76628 171192 76634
rect 171140 76570 171192 76576
rect 170680 75744 170732 75750
rect 170680 75686 170732 75692
rect 170772 75268 170824 75274
rect 170772 75210 170824 75216
rect 170680 75064 170732 75070
rect 170680 75006 170732 75012
rect 170588 68332 170640 68338
rect 170588 68274 170640 68280
rect 170312 66972 170364 66978
rect 170312 66914 170364 66920
rect 170220 65680 170272 65686
rect 170220 65622 170272 65628
rect 170402 63608 170458 63617
rect 170402 63543 170458 63552
rect 170128 60104 170180 60110
rect 170128 60046 170180 60052
rect 170036 22976 170088 22982
rect 170036 22918 170088 22924
rect 169944 19984 169996 19990
rect 169944 19926 169996 19932
rect 169852 7676 169904 7682
rect 169852 7618 169904 7624
rect 167000 7608 167052 7614
rect 167000 7550 167052 7556
rect 165712 6316 165764 6322
rect 165712 6258 165764 6264
rect 165620 6248 165672 6254
rect 165620 6190 165672 6196
rect 164240 5092 164292 5098
rect 164240 5034 164292 5040
rect 162490 4992 162546 5001
rect 162490 4927 162546 4936
rect 159364 3800 159416 3806
rect 159364 3742 159416 3748
rect 160100 3732 160152 3738
rect 160100 3674 160152 3680
rect 158904 3256 158956 3262
rect 158904 3198 158956 3204
rect 158916 480 158944 3198
rect 160112 480 160140 3674
rect 161294 3496 161350 3505
rect 161294 3431 161350 3440
rect 161308 480 161336 3431
rect 162504 480 162532 4927
rect 167184 4888 167236 4894
rect 166078 4856 166134 4865
rect 167184 4830 167236 4836
rect 166078 4791 166134 4800
rect 164884 3664 164936 3670
rect 164884 3606 164936 3612
rect 163686 3360 163742 3369
rect 163686 3295 163742 3304
rect 163700 480 163728 3295
rect 164896 480 164924 3606
rect 166092 480 166120 4791
rect 167196 480 167224 4830
rect 169576 4820 169628 4826
rect 169576 4762 169628 4768
rect 168380 3528 168432 3534
rect 168380 3470 168432 3476
rect 168392 480 168420 3470
rect 169588 480 169616 4762
rect 170416 3534 170444 63543
rect 170692 3942 170720 75006
rect 170784 16574 170812 75210
rect 171140 75200 171192 75206
rect 171140 75142 171192 75148
rect 170784 16546 170904 16574
rect 170772 6180 170824 6186
rect 170772 6122 170824 6128
rect 170680 3936 170732 3942
rect 170680 3878 170732 3884
rect 170404 3528 170456 3534
rect 170404 3470 170456 3476
rect 170784 480 170812 6122
rect 170876 5030 170904 16546
rect 170864 5024 170916 5030
rect 170864 4966 170916 4972
rect 171152 4962 171180 75142
rect 171244 8974 171272 79478
rect 171416 79416 171468 79422
rect 171416 79358 171468 79364
rect 171428 79218 171456 79358
rect 171416 79212 171468 79218
rect 171416 79154 171468 79160
rect 171520 79014 171548 79716
rect 171934 79744 171962 80036
rect 172026 79830 172054 80036
rect 172014 79824 172066 79830
rect 172014 79766 172066 79772
rect 171784 79698 171836 79704
rect 171888 79716 171962 79744
rect 171690 79656 171746 79665
rect 171690 79591 171746 79600
rect 171600 79484 171652 79490
rect 171600 79426 171652 79432
rect 171508 79008 171560 79014
rect 171508 78950 171560 78956
rect 171612 78792 171640 79426
rect 171428 78764 171640 78792
rect 171324 78396 171376 78402
rect 171324 78338 171376 78344
rect 171336 15910 171364 78338
rect 171428 17270 171456 78764
rect 171704 78690 171732 79591
rect 171612 78662 171732 78690
rect 171508 78532 171560 78538
rect 171508 78474 171560 78480
rect 171520 75410 171548 78474
rect 171612 78402 171640 78662
rect 171600 78396 171652 78402
rect 171600 78338 171652 78344
rect 171598 78296 171654 78305
rect 171598 78231 171654 78240
rect 171508 75404 171560 75410
rect 171508 75346 171560 75352
rect 171508 75268 171560 75274
rect 171508 75210 171560 75216
rect 171520 22846 171548 75210
rect 171612 22914 171640 78231
rect 171692 77852 171744 77858
rect 171692 77794 171744 77800
rect 171704 61402 171732 77794
rect 171796 66910 171824 79698
rect 171888 79490 171916 79716
rect 172118 79676 172146 80036
rect 172210 79830 172238 80036
rect 172302 79830 172330 80036
rect 172198 79824 172250 79830
rect 172198 79766 172250 79772
rect 172290 79824 172342 79830
rect 172394 79801 172422 80036
rect 172486 79937 172514 80036
rect 172578 79966 172606 80036
rect 172566 79960 172618 79966
rect 172472 79928 172528 79937
rect 172670 79937 172698 80036
rect 172566 79902 172618 79908
rect 172656 79928 172712 79937
rect 172472 79863 172528 79872
rect 172656 79863 172712 79872
rect 172290 79766 172342 79772
rect 172380 79792 172436 79801
rect 172762 79778 172790 80036
rect 172854 79898 172882 80036
rect 172946 79937 172974 80036
rect 173038 79966 173066 80036
rect 173026 79960 173078 79966
rect 172932 79928 172988 79937
rect 172842 79892 172894 79898
rect 173026 79902 173078 79908
rect 172932 79863 172988 79872
rect 172842 79834 172894 79840
rect 172978 79792 173034 79801
rect 172762 79750 172836 79778
rect 172380 79727 172436 79736
rect 172118 79648 172376 79676
rect 171968 79620 172020 79626
rect 171968 79562 172020 79568
rect 171876 79484 171928 79490
rect 171876 79426 171928 79432
rect 171876 79280 171928 79286
rect 171876 79222 171928 79228
rect 171888 78878 171916 79222
rect 171876 78872 171928 78878
rect 171876 78814 171928 78820
rect 171876 77172 171928 77178
rect 171876 77114 171928 77120
rect 171888 76498 171916 77114
rect 171876 76492 171928 76498
rect 171876 76434 171928 76440
rect 171980 75274 172008 79562
rect 172152 79552 172204 79558
rect 172152 79494 172204 79500
rect 172244 79552 172296 79558
rect 172244 79494 172296 79500
rect 172060 79484 172112 79490
rect 172060 79426 172112 79432
rect 172072 79082 172100 79426
rect 172060 79076 172112 79082
rect 172060 79018 172112 79024
rect 172058 78704 172114 78713
rect 172058 78639 172114 78648
rect 172072 78305 172100 78639
rect 172058 78296 172114 78305
rect 172058 78231 172114 78240
rect 172164 77489 172192 79494
rect 172256 78169 172284 79494
rect 172242 78160 172298 78169
rect 172242 78095 172298 78104
rect 172150 77480 172206 77489
rect 172150 77415 172206 77424
rect 172060 76764 172112 76770
rect 172060 76706 172112 76712
rect 172072 76430 172100 76706
rect 172060 76424 172112 76430
rect 172060 76366 172112 76372
rect 172348 75914 172376 79648
rect 172428 79620 172480 79626
rect 172428 79562 172480 79568
rect 172440 77294 172468 79562
rect 172610 79520 172666 79529
rect 172610 79455 172666 79464
rect 172624 79150 172652 79455
rect 172612 79144 172664 79150
rect 172612 79086 172664 79092
rect 172612 78940 172664 78946
rect 172612 78882 172664 78888
rect 172624 77926 172652 78882
rect 172702 78704 172758 78713
rect 172702 78639 172758 78648
rect 172612 77920 172664 77926
rect 172612 77862 172664 77868
rect 172440 77266 172652 77294
rect 172256 75886 172376 75914
rect 171968 75268 172020 75274
rect 171968 75210 172020 75216
rect 172256 75206 172284 75886
rect 172624 75274 172652 77266
rect 172612 75268 172664 75274
rect 172612 75210 172664 75216
rect 172244 75200 172296 75206
rect 172244 75142 172296 75148
rect 172612 75132 172664 75138
rect 172612 75074 172664 75080
rect 171784 66904 171836 66910
rect 171784 66846 171836 66852
rect 171692 61396 171744 61402
rect 171692 61338 171744 61344
rect 171600 22908 171652 22914
rect 171600 22850 171652 22856
rect 171508 22840 171560 22846
rect 171508 22782 171560 22788
rect 171416 17264 171468 17270
rect 171416 17206 171468 17212
rect 171324 15904 171376 15910
rect 171324 15846 171376 15852
rect 172624 14482 172652 75074
rect 172716 18834 172744 78639
rect 172808 24206 172836 79750
rect 173130 79778 173158 80036
rect 173222 79966 173250 80036
rect 173210 79960 173262 79966
rect 173210 79902 173262 79908
rect 173034 79750 173158 79778
rect 172978 79727 173034 79736
rect 172888 79688 172940 79694
rect 173164 79688 173216 79694
rect 172888 79630 172940 79636
rect 172978 79656 173034 79665
rect 172900 25770 172928 79630
rect 172978 79591 173034 79600
rect 173162 79656 173164 79665
rect 173314 79676 173342 80036
rect 173406 79744 173434 80036
rect 173498 79898 173526 80036
rect 173590 79971 173618 80036
rect 173576 79962 173632 79971
rect 173486 79892 173538 79898
rect 173576 79897 173632 79906
rect 173486 79834 173538 79840
rect 173530 79792 173586 79801
rect 173406 79716 173480 79744
rect 173682 79778 173710 80036
rect 173586 79750 173710 79778
rect 173530 79727 173586 79736
rect 173216 79656 173218 79665
rect 173314 79648 173388 79676
rect 173162 79591 173218 79600
rect 172888 25764 172940 25770
rect 172888 25706 172940 25712
rect 172992 25566 173020 79591
rect 173164 79552 173216 79558
rect 173164 79494 173216 79500
rect 173070 78160 173126 78169
rect 173070 78095 173126 78104
rect 173084 77314 173112 78095
rect 173072 77308 173124 77314
rect 173072 77250 173124 77256
rect 173176 76430 173204 79494
rect 173256 79008 173308 79014
rect 173254 78976 173256 78985
rect 173308 78976 173310 78985
rect 173254 78911 173310 78920
rect 173164 76424 173216 76430
rect 173164 76366 173216 76372
rect 173072 75268 173124 75274
rect 173072 75210 173124 75216
rect 173084 28286 173112 75210
rect 173360 75138 173388 79648
rect 173452 75206 173480 79716
rect 173774 79676 173802 80036
rect 173866 79898 173894 80036
rect 173854 79892 173906 79898
rect 173854 79834 173906 79840
rect 173958 79744 173986 80036
rect 174050 79971 174078 80036
rect 174036 79962 174092 79971
rect 174036 79897 174092 79906
rect 174142 79812 174170 80036
rect 174234 79898 174262 80036
rect 174326 79898 174354 80036
rect 174222 79892 174274 79898
rect 174222 79834 174274 79840
rect 174314 79892 174366 79898
rect 174314 79834 174366 79840
rect 174096 79784 174170 79812
rect 173958 79716 174032 79744
rect 173530 79656 173586 79665
rect 173530 79591 173586 79600
rect 173636 79648 173802 79676
rect 173854 79688 173906 79694
rect 173440 75200 173492 75206
rect 173440 75142 173492 75148
rect 173348 75132 173400 75138
rect 173348 75074 173400 75080
rect 173544 70394 173572 79591
rect 173636 78985 173664 79648
rect 173854 79630 173906 79636
rect 173714 79520 173770 79529
rect 173866 79506 173894 79630
rect 173714 79455 173770 79464
rect 173820 79478 173894 79506
rect 173622 78976 173678 78985
rect 173622 78911 173678 78920
rect 173728 70394 173756 79455
rect 173820 78713 173848 79478
rect 173806 78704 173862 78713
rect 173806 78639 173862 78648
rect 173544 70366 173664 70394
rect 173728 70366 173848 70394
rect 173072 28280 173124 28286
rect 173072 28222 173124 28228
rect 172980 25560 173032 25566
rect 172980 25502 173032 25508
rect 172796 24200 172848 24206
rect 172796 24142 172848 24148
rect 172704 18828 172756 18834
rect 172704 18770 172756 18776
rect 172612 14476 172664 14482
rect 172612 14418 172664 14424
rect 171232 8968 171284 8974
rect 171232 8910 171284 8916
rect 173164 5228 173216 5234
rect 173164 5170 173216 5176
rect 171140 4956 171192 4962
rect 171140 4898 171192 4904
rect 171968 3596 172020 3602
rect 171968 3538 172020 3544
rect 171980 480 172008 3538
rect 173176 480 173204 5170
rect 173636 4894 173664 70366
rect 173820 64190 173848 70366
rect 173808 64184 173860 64190
rect 173808 64126 173860 64132
rect 174004 18766 174032 79716
rect 173992 18760 174044 18766
rect 173992 18702 174044 18708
rect 174096 18698 174124 79784
rect 174418 79778 174446 80036
rect 174510 79830 174538 80036
rect 174280 79750 174446 79778
rect 174498 79824 174550 79830
rect 174498 79766 174550 79772
rect 174176 79688 174228 79694
rect 174176 79630 174228 79636
rect 174084 18692 174136 18698
rect 174084 18634 174136 18640
rect 174188 18630 174216 79630
rect 174280 21418 174308 79750
rect 174360 79688 174412 79694
rect 174360 79630 174412 79636
rect 174452 79688 174504 79694
rect 174602 79676 174630 80036
rect 174694 79812 174722 80036
rect 174786 79966 174814 80036
rect 174774 79960 174826 79966
rect 174774 79902 174826 79908
rect 174694 79784 174768 79812
rect 174452 79630 174504 79636
rect 174556 79648 174630 79676
rect 174372 75274 174400 79630
rect 174360 75268 174412 75274
rect 174360 75210 174412 75216
rect 174360 75132 174412 75138
rect 174360 75074 174412 75080
rect 174372 24138 174400 75074
rect 174464 29646 174492 79630
rect 174556 65618 174584 79648
rect 174636 78668 174688 78674
rect 174636 78610 174688 78616
rect 174544 65612 174596 65618
rect 174544 65554 174596 65560
rect 174648 65550 174676 78610
rect 174740 77294 174768 79784
rect 174878 79778 174906 80036
rect 174970 79801 174998 80036
rect 174832 79750 174906 79778
rect 174956 79792 175012 79801
rect 174832 78674 174860 79750
rect 175062 79778 175090 80036
rect 175154 79966 175182 80036
rect 175142 79960 175194 79966
rect 175246 79937 175274 80036
rect 175142 79902 175194 79908
rect 175232 79928 175288 79937
rect 175338 79898 175366 80036
rect 175430 79966 175458 80036
rect 175418 79960 175470 79966
rect 175522 79937 175550 80036
rect 175614 79966 175642 80036
rect 175602 79960 175654 79966
rect 175418 79902 175470 79908
rect 175508 79928 175564 79937
rect 175232 79863 175288 79872
rect 175326 79892 175378 79898
rect 175602 79902 175654 79908
rect 175508 79863 175564 79872
rect 175326 79834 175378 79840
rect 175062 79750 175136 79778
rect 174956 79727 175012 79736
rect 174912 79688 174964 79694
rect 174912 79630 174964 79636
rect 175004 79688 175056 79694
rect 175004 79630 175056 79636
rect 174924 78674 174952 79630
rect 175016 78713 175044 79630
rect 175108 78985 175136 79750
rect 175464 79756 175516 79762
rect 175464 79698 175516 79704
rect 175556 79756 175608 79762
rect 175556 79698 175608 79704
rect 175186 79656 175242 79665
rect 175186 79591 175188 79600
rect 175240 79591 175242 79600
rect 175372 79620 175424 79626
rect 175188 79562 175240 79568
rect 175372 79562 175424 79568
rect 175280 79348 175332 79354
rect 175280 79290 175332 79296
rect 175292 79257 175320 79290
rect 175278 79248 175334 79257
rect 175278 79183 175334 79192
rect 175094 78976 175150 78985
rect 175094 78911 175150 78920
rect 175002 78704 175058 78713
rect 174820 78668 174872 78674
rect 174820 78610 174872 78616
rect 174912 78668 174964 78674
rect 175002 78639 175058 78648
rect 175188 78668 175240 78674
rect 174912 78610 174964 78616
rect 175188 78610 175240 78616
rect 174740 77266 174860 77294
rect 174728 75268 174780 75274
rect 174728 75210 174780 75216
rect 174740 69698 174768 75210
rect 174832 70394 174860 77266
rect 175096 75812 175148 75818
rect 175096 75754 175148 75760
rect 175004 75744 175056 75750
rect 175004 75686 175056 75692
rect 175016 75410 175044 75686
rect 175108 75478 175136 75754
rect 175096 75472 175148 75478
rect 175096 75414 175148 75420
rect 175004 75404 175056 75410
rect 175004 75346 175056 75352
rect 175200 75138 175228 78610
rect 175278 77888 175334 77897
rect 175278 77823 175334 77832
rect 175188 75132 175240 75138
rect 175188 75074 175240 75080
rect 175292 72894 175320 77823
rect 175280 72888 175332 72894
rect 175280 72830 175332 72836
rect 175280 71052 175332 71058
rect 175280 70994 175332 71000
rect 174832 70366 174952 70394
rect 174728 69692 174780 69698
rect 174728 69634 174780 69640
rect 174636 65544 174688 65550
rect 174636 65486 174688 65492
rect 174452 29640 174504 29646
rect 174452 29582 174504 29588
rect 174360 24132 174412 24138
rect 174360 24074 174412 24080
rect 174268 21412 174320 21418
rect 174268 21354 174320 21360
rect 174176 18624 174228 18630
rect 174176 18566 174228 18572
rect 174268 5160 174320 5166
rect 174268 5102 174320 5108
rect 173624 4888 173676 4894
rect 173624 4830 173676 4836
rect 174280 480 174308 5102
rect 174924 4826 174952 70366
rect 175292 16574 175320 70994
rect 175384 26926 175412 79562
rect 175476 78713 175504 79698
rect 175568 78985 175596 79698
rect 175706 79608 175734 80036
rect 175798 79801 175826 80036
rect 175890 79898 175918 80036
rect 175982 79966 176010 80036
rect 175970 79960 176022 79966
rect 175970 79902 176022 79908
rect 176074 79898 176102 80036
rect 175878 79892 175930 79898
rect 175878 79834 175930 79840
rect 176062 79892 176114 79898
rect 176062 79834 176114 79840
rect 176166 79830 176194 80036
rect 176258 79898 176286 80036
rect 176246 79892 176298 79898
rect 176246 79834 176298 79840
rect 176154 79824 176206 79830
rect 175784 79792 175840 79801
rect 176154 79766 176206 79772
rect 176350 79778 176378 80036
rect 176442 79898 176470 80036
rect 176534 79971 176562 80036
rect 176520 79962 176576 79971
rect 176626 79966 176654 80036
rect 176718 79966 176746 80036
rect 176430 79892 176482 79898
rect 176520 79897 176576 79906
rect 176614 79960 176666 79966
rect 176614 79902 176666 79908
rect 176706 79960 176758 79966
rect 176810 79937 176838 80036
rect 176706 79902 176758 79908
rect 176796 79928 176852 79937
rect 176796 79863 176852 79872
rect 176430 79834 176482 79840
rect 176752 79824 176804 79830
rect 176750 79792 176752 79801
rect 176902 79812 176930 80036
rect 176804 79792 176806 79801
rect 176350 79750 176516 79778
rect 175784 79727 175840 79736
rect 176062 79688 176114 79694
rect 176114 79648 176194 79676
rect 176488 79665 176516 79750
rect 176568 79756 176620 79762
rect 176750 79727 176806 79736
rect 176856 79784 176930 79812
rect 176994 79812 177022 80036
rect 177086 79966 177114 80036
rect 177178 79966 177206 80036
rect 177074 79960 177126 79966
rect 177074 79902 177126 79908
rect 177166 79960 177218 79966
rect 177166 79902 177218 79908
rect 177270 79898 177298 80036
rect 177362 79937 177390 80036
rect 177348 79928 177404 79937
rect 177258 79892 177310 79898
rect 177348 79863 177404 79872
rect 177258 79834 177310 79840
rect 176994 79784 177068 79812
rect 176568 79698 176620 79704
rect 176062 79630 176114 79636
rect 175924 79620 175976 79626
rect 175706 79580 175780 79608
rect 175648 79212 175700 79218
rect 175648 79154 175700 79160
rect 175660 79121 175688 79154
rect 175646 79112 175702 79121
rect 175646 79047 175702 79056
rect 175554 78976 175610 78985
rect 175554 78911 175610 78920
rect 175462 78704 175518 78713
rect 175462 78639 175518 78648
rect 175752 78402 175780 79580
rect 175924 79562 175976 79568
rect 175740 78396 175792 78402
rect 175740 78338 175792 78344
rect 175830 78160 175886 78169
rect 175936 78130 175964 79562
rect 176166 79540 176194 79648
rect 176474 79656 176530 79665
rect 176474 79591 176530 79600
rect 176120 79512 176194 79540
rect 175830 78095 175886 78104
rect 175924 78124 175976 78130
rect 175844 78010 175872 78095
rect 175924 78066 175976 78072
rect 175844 77982 175964 78010
rect 175832 77376 175884 77382
rect 175832 77318 175884 77324
rect 175844 73098 175872 77318
rect 175832 73092 175884 73098
rect 175832 73034 175884 73040
rect 175936 64874 175964 77982
rect 176120 75914 176148 79512
rect 176290 79384 176346 79393
rect 176200 79348 176252 79354
rect 176290 79319 176292 79328
rect 176200 79290 176252 79296
rect 176344 79319 176346 79328
rect 176292 79290 176344 79296
rect 176212 79218 176240 79290
rect 176200 79212 176252 79218
rect 176200 79154 176252 79160
rect 176580 78674 176608 79698
rect 176660 79688 176712 79694
rect 176856 79676 176884 79784
rect 176660 79630 176712 79636
rect 176810 79648 176884 79676
rect 176672 79393 176700 79630
rect 176810 79608 176838 79648
rect 176810 79580 176884 79608
rect 176658 79384 176714 79393
rect 176658 79319 176714 79328
rect 176752 79144 176804 79150
rect 176752 79086 176804 79092
rect 176200 78668 176252 78674
rect 176200 78610 176252 78616
rect 176568 78668 176620 78674
rect 176568 78610 176620 78616
rect 176028 75886 176148 75914
rect 176028 73166 176056 75886
rect 176106 75712 176162 75721
rect 176106 75647 176162 75656
rect 176016 73160 176068 73166
rect 176016 73102 176068 73108
rect 176120 72978 176148 75647
rect 176212 73302 176240 78610
rect 176476 78600 176528 78606
rect 176476 78542 176528 78548
rect 176292 77580 176344 77586
rect 176292 77522 176344 77528
rect 176200 73296 176252 73302
rect 176200 73238 176252 73244
rect 176200 73092 176252 73098
rect 176200 73034 176252 73040
rect 175752 64846 175964 64874
rect 176028 72950 176148 72978
rect 175372 26920 175424 26926
rect 175372 26862 175424 26868
rect 175292 16546 175504 16574
rect 174912 4820 174964 4826
rect 174912 4762 174964 4768
rect 175476 480 175504 16546
rect 175752 3505 175780 64846
rect 176028 3738 176056 72950
rect 176108 72888 176160 72894
rect 176108 72830 176160 72836
rect 176120 7818 176148 72830
rect 176212 35358 176240 73034
rect 176200 35352 176252 35358
rect 176200 35294 176252 35300
rect 176304 35290 176332 77522
rect 176384 77308 176436 77314
rect 176384 77250 176436 77256
rect 176396 60042 176424 77250
rect 176488 71058 176516 78542
rect 176764 77314 176792 79086
rect 176856 77858 176884 79580
rect 177040 78538 177068 79784
rect 177304 79688 177356 79694
rect 177304 79630 177356 79636
rect 177454 79642 177482 80036
rect 177546 79966 177574 80036
rect 177638 79966 177666 80036
rect 177534 79960 177586 79966
rect 177534 79902 177586 79908
rect 177626 79960 177678 79966
rect 177626 79902 177678 79908
rect 177580 79824 177632 79830
rect 177730 79812 177758 80036
rect 177822 79937 177850 80036
rect 177914 79966 177942 80036
rect 177902 79960 177954 79966
rect 177808 79928 177864 79937
rect 177902 79902 177954 79908
rect 177808 79863 177864 79872
rect 177730 79801 177804 79812
rect 177730 79792 177818 79801
rect 177730 79784 177762 79792
rect 177580 79766 177632 79772
rect 177120 79620 177172 79626
rect 177120 79562 177172 79568
rect 177212 79620 177264 79626
rect 177212 79562 177264 79568
rect 177132 78606 177160 79562
rect 177224 78849 177252 79562
rect 177210 78840 177266 78849
rect 177210 78775 177266 78784
rect 177120 78600 177172 78606
rect 177120 78542 177172 78548
rect 177028 78532 177080 78538
rect 177028 78474 177080 78480
rect 176934 78432 176990 78441
rect 176934 78367 176990 78376
rect 176948 78169 176976 78367
rect 176934 78160 176990 78169
rect 176934 78095 176990 78104
rect 176844 77852 176896 77858
rect 176844 77794 176896 77800
rect 177316 77790 177344 79630
rect 177454 79614 177528 79642
rect 177500 78849 177528 79614
rect 177592 79393 177620 79766
rect 177762 79727 177818 79736
rect 177856 79756 177908 79762
rect 178006 79744 178034 80036
rect 178098 79966 178126 80036
rect 178086 79960 178138 79966
rect 178086 79902 178138 79908
rect 178190 79898 178218 80036
rect 178178 79892 178230 79898
rect 178178 79834 178230 79840
rect 178086 79824 178138 79830
rect 178282 79812 178310 80036
rect 178374 79937 178402 80036
rect 178360 79928 178416 79937
rect 178360 79863 178416 79872
rect 178282 79784 178356 79812
rect 178138 79772 178218 79778
rect 178086 79766 178218 79772
rect 178098 79750 178218 79766
rect 177856 79698 177908 79704
rect 177960 79716 178034 79744
rect 177672 79688 177724 79694
rect 177764 79688 177816 79694
rect 177672 79630 177724 79636
rect 177762 79656 177764 79665
rect 177816 79656 177818 79665
rect 177578 79384 177634 79393
rect 177578 79319 177634 79328
rect 177684 78985 177712 79630
rect 177762 79591 177818 79600
rect 177868 79268 177896 79698
rect 177960 79626 177988 79716
rect 178190 79676 178218 79750
rect 178144 79648 178218 79676
rect 177948 79620 178000 79626
rect 177948 79562 178000 79568
rect 178040 79620 178092 79626
rect 178040 79562 178092 79568
rect 177868 79240 177988 79268
rect 178052 79257 178080 79562
rect 178144 79354 178172 79648
rect 178224 79484 178276 79490
rect 178224 79426 178276 79432
rect 178132 79348 178184 79354
rect 178132 79290 178184 79296
rect 178236 79257 178264 79426
rect 177670 78976 177726 78985
rect 177670 78911 177726 78920
rect 177486 78840 177542 78849
rect 177486 78775 177542 78784
rect 177856 78736 177908 78742
rect 177856 78678 177908 78684
rect 177672 78464 177724 78470
rect 177578 78432 177634 78441
rect 177672 78406 177724 78412
rect 177578 78367 177634 78376
rect 177488 78328 177540 78334
rect 177488 78270 177540 78276
rect 177396 77920 177448 77926
rect 177396 77862 177448 77868
rect 177304 77784 177356 77790
rect 177304 77726 177356 77732
rect 177212 77716 177264 77722
rect 177212 77658 177264 77664
rect 176752 77308 176804 77314
rect 176752 77250 176804 77256
rect 176752 75676 176804 75682
rect 176752 75618 176804 75624
rect 176566 74488 176622 74497
rect 176566 74423 176622 74432
rect 176476 71052 176528 71058
rect 176476 70994 176528 71000
rect 176384 60036 176436 60042
rect 176384 59978 176436 59984
rect 176292 35284 176344 35290
rect 176292 35226 176344 35232
rect 176108 7812 176160 7818
rect 176108 7754 176160 7760
rect 176580 6186 176608 74423
rect 176764 16574 176792 75618
rect 177224 44878 177252 77658
rect 177304 77648 177356 77654
rect 177304 77590 177356 77596
rect 177212 44872 177264 44878
rect 177212 44814 177264 44820
rect 176764 16546 177252 16574
rect 176568 6180 176620 6186
rect 176568 6122 176620 6128
rect 176016 3732 176068 3738
rect 176016 3674 176068 3680
rect 175738 3496 175794 3505
rect 175738 3431 175794 3440
rect 176660 3460 176712 3466
rect 176660 3402 176712 3408
rect 176672 480 176700 3402
rect 177224 3074 177252 16546
rect 177316 3602 177344 77590
rect 177408 3670 177436 77862
rect 177500 8770 177528 78270
rect 177592 24274 177620 78367
rect 177684 77568 177712 78406
rect 177684 77540 177804 77568
rect 177672 77444 177724 77450
rect 177672 77386 177724 77392
rect 177580 24268 177632 24274
rect 177580 24210 177632 24216
rect 177488 8764 177540 8770
rect 177488 8706 177540 8712
rect 177396 3664 177448 3670
rect 177396 3606 177448 3612
rect 177304 3596 177356 3602
rect 177304 3538 177356 3544
rect 177684 3194 177712 77386
rect 177776 25702 177804 77540
rect 177868 77450 177896 78678
rect 177960 78470 177988 79240
rect 178038 79248 178094 79257
rect 178038 79183 178094 79192
rect 178222 79248 178278 79257
rect 178328 79218 178356 79784
rect 178466 79778 178494 80036
rect 178558 79898 178586 80036
rect 178546 79892 178598 79898
rect 178546 79834 178598 79840
rect 178650 79812 178678 80036
rect 178742 79966 178770 80036
rect 178730 79960 178782 79966
rect 178730 79902 178782 79908
rect 178650 79784 178724 79812
rect 178466 79750 178540 79778
rect 178512 79744 178540 79750
rect 178512 79716 178632 79744
rect 178408 79688 178460 79694
rect 178408 79630 178460 79636
rect 178222 79183 178278 79192
rect 178316 79212 178368 79218
rect 178316 79154 178368 79160
rect 178420 78810 178448 79630
rect 178500 79620 178552 79626
rect 178500 79562 178552 79568
rect 178512 78878 178540 79562
rect 178604 79014 178632 79716
rect 178696 79642 178724 79784
rect 178834 79642 178862 80036
rect 178926 79898 178954 80036
rect 178914 79892 178966 79898
rect 178914 79834 178966 79840
rect 179018 79830 179046 80036
rect 179006 79824 179058 79830
rect 179006 79766 179058 79772
rect 179110 79778 179138 80036
rect 179202 79966 179230 80036
rect 179190 79960 179242 79966
rect 179190 79902 179242 79908
rect 179110 79762 179184 79778
rect 179110 79756 179196 79762
rect 179110 79750 179144 79756
rect 179294 79744 179322 80036
rect 179144 79698 179196 79704
rect 179248 79716 179322 79744
rect 179386 79744 179414 80036
rect 179524 79966 179552 80582
rect 179616 80170 179644 80679
rect 179788 80650 179840 80656
rect 179696 80436 179748 80442
rect 179696 80378 179748 80384
rect 179604 80164 179656 80170
rect 179604 80106 179656 80112
rect 179708 80034 179736 80378
rect 179696 80028 179748 80034
rect 179696 79970 179748 79976
rect 179512 79960 179564 79966
rect 179512 79902 179564 79908
rect 179696 79892 179748 79898
rect 179696 79834 179748 79840
rect 179386 79716 179460 79744
rect 178696 79614 178770 79642
rect 178834 79614 178908 79642
rect 178742 79506 178770 79614
rect 178696 79478 178770 79506
rect 178696 79286 178724 79478
rect 178880 79422 178908 79614
rect 179144 79620 179196 79626
rect 179144 79562 179196 79568
rect 178868 79416 178920 79422
rect 178868 79358 178920 79364
rect 178684 79280 178736 79286
rect 178684 79222 178736 79228
rect 179156 79121 179184 79562
rect 179142 79112 179198 79121
rect 179142 79047 179198 79056
rect 178592 79008 178644 79014
rect 178592 78950 178644 78956
rect 178500 78872 178552 78878
rect 178500 78814 178552 78820
rect 179248 78810 179276 79716
rect 178408 78804 178460 78810
rect 178408 78746 178460 78752
rect 178592 78804 178644 78810
rect 178592 78746 178644 78752
rect 179236 78804 179288 78810
rect 179236 78746 179288 78752
rect 177948 78464 178000 78470
rect 177948 78406 178000 78412
rect 177856 77444 177908 77450
rect 177856 77386 177908 77392
rect 178132 77444 178184 77450
rect 178132 77386 178184 77392
rect 177856 77308 177908 77314
rect 177856 77250 177908 77256
rect 177764 25696 177816 25702
rect 177764 25638 177816 25644
rect 177868 16574 177896 77250
rect 177948 73296 178000 73302
rect 177948 73238 178000 73244
rect 177960 33114 177988 73238
rect 178040 69964 178092 69970
rect 178040 69906 178092 69912
rect 177948 33108 178000 33114
rect 177948 33050 178000 33056
rect 178052 16574 178080 69906
rect 178144 32706 178172 77386
rect 178604 70394 178632 78746
rect 179432 77450 179460 79716
rect 179708 78305 179736 79834
rect 179800 79762 179828 80650
rect 180248 80572 180300 80578
rect 180248 80514 180300 80520
rect 179878 80472 179934 80481
rect 179878 80407 179934 80416
rect 179892 80102 179920 80407
rect 180062 80336 180118 80345
rect 180062 80271 180118 80280
rect 179972 80232 180024 80238
rect 179972 80174 180024 80180
rect 179880 80096 179932 80102
rect 179880 80038 179932 80044
rect 179788 79756 179840 79762
rect 179788 79698 179840 79704
rect 179984 79694 180012 80174
rect 179972 79688 180024 79694
rect 179972 79630 180024 79636
rect 179786 79520 179842 79529
rect 179786 79455 179842 79464
rect 179800 79354 179828 79455
rect 179788 79348 179840 79354
rect 179788 79290 179840 79296
rect 180076 79218 180104 80271
rect 180260 80170 180288 80514
rect 180706 80200 180762 80209
rect 180156 80164 180208 80170
rect 180156 80106 180208 80112
rect 180248 80164 180300 80170
rect 180706 80135 180762 80144
rect 180248 80106 180300 80112
rect 180168 79286 180196 80106
rect 180246 80064 180302 80073
rect 180246 79999 180302 80008
rect 180156 79280 180208 79286
rect 180156 79222 180208 79228
rect 180064 79212 180116 79218
rect 180064 79154 180116 79160
rect 180260 78713 180288 79999
rect 180720 79150 180748 80135
rect 180708 79144 180760 79150
rect 180708 79086 180760 79092
rect 180246 78704 180302 78713
rect 180246 78639 180302 78648
rect 189368 78470 189396 700334
rect 198004 700324 198056 700330
rect 198004 700266 198056 700272
rect 196624 683188 196676 683194
rect 196624 683130 196676 683136
rect 191104 643136 191156 643142
rect 191104 643078 191156 643084
rect 190460 618316 190512 618322
rect 190460 618258 190512 618264
rect 189448 409896 189500 409902
rect 189448 409838 189500 409844
rect 189460 126177 189488 409838
rect 189724 149116 189776 149122
rect 189724 149058 189776 149064
rect 189632 148368 189684 148374
rect 189632 148310 189684 148316
rect 189538 137048 189594 137057
rect 189538 136983 189594 136992
rect 189446 126168 189502 126177
rect 189446 126103 189502 126112
rect 189448 118652 189500 118658
rect 189448 118594 189500 118600
rect 189460 118561 189488 118594
rect 189446 118552 189502 118561
rect 189446 118487 189502 118496
rect 189448 117292 189500 117298
rect 189448 117234 189500 117240
rect 189460 117201 189488 117234
rect 189446 117192 189502 117201
rect 189446 117127 189502 117136
rect 189448 114504 189500 114510
rect 189448 114446 189500 114452
rect 189460 114209 189488 114446
rect 189446 114200 189502 114209
rect 189446 114135 189502 114144
rect 189356 78464 189408 78470
rect 189356 78406 189408 78412
rect 187608 78396 187660 78402
rect 187608 78338 187660 78344
rect 179694 78296 179750 78305
rect 186148 78266 186452 78282
rect 179694 78231 179750 78240
rect 186136 78260 186464 78266
rect 186188 78254 186412 78260
rect 186136 78202 186188 78208
rect 186412 78202 186464 78208
rect 187620 78198 187648 78338
rect 180156 78192 180208 78198
rect 187608 78192 187660 78198
rect 180156 78134 180208 78140
rect 180246 78160 180302 78169
rect 179420 77444 179472 77450
rect 179420 77386 179472 77392
rect 178684 76492 178736 76498
rect 178684 76434 178736 76440
rect 178236 70366 178632 70394
rect 178236 45558 178264 70366
rect 178224 45552 178276 45558
rect 178224 45494 178276 45500
rect 178132 32700 178184 32706
rect 178132 32642 178184 32648
rect 177868 16546 177988 16574
rect 178052 16546 178632 16574
rect 177960 3466 177988 16546
rect 177948 3460 178000 3466
rect 177948 3402 178000 3408
rect 177672 3188 177724 3194
rect 177672 3130 177724 3136
rect 177224 3046 177896 3074
rect 177868 480 177896 3046
rect 156574 354 156686 480
rect 156156 326 156686 354
rect 156574 -960 156686 326
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 178604 354 178632 16546
rect 178696 3330 178724 76434
rect 180062 76392 180118 76401
rect 180062 76327 180118 76336
rect 178684 3324 178736 3330
rect 178684 3266 178736 3272
rect 180076 3262 180104 76327
rect 180168 10402 180196 78134
rect 187608 78134 187660 78140
rect 180246 78095 180302 78104
rect 180260 13190 180288 78095
rect 181444 77512 181496 77518
rect 181444 77454 181496 77460
rect 180798 75576 180854 75585
rect 180798 75511 180854 75520
rect 180812 16574 180840 75511
rect 180812 16546 181024 16574
rect 180248 13184 180300 13190
rect 180248 13126 180300 13132
rect 180156 10396 180208 10402
rect 180156 10338 180208 10344
rect 180248 3800 180300 3806
rect 180248 3742 180300 3748
rect 180064 3256 180116 3262
rect 180064 3198 180116 3204
rect 180260 480 180288 3742
rect 179022 354 179134 480
rect 178604 326 179134 354
rect 179022 -960 179134 326
rect 180218 -960 180330 480
rect 180996 354 181024 16546
rect 181456 14550 181484 77454
rect 186320 77240 186372 77246
rect 186320 77182 186372 77188
rect 185584 74248 185636 74254
rect 185584 74190 185636 74196
rect 182178 69592 182234 69601
rect 182178 69527 182234 69536
rect 181444 14544 181496 14550
rect 181444 14486 181496 14492
rect 181414 354 181526 480
rect 180996 326 181526 354
rect 182192 354 182220 69527
rect 185032 31408 185084 31414
rect 185032 31350 185084 31356
rect 183558 25664 183614 25673
rect 183558 25599 183614 25608
rect 183572 16574 183600 25599
rect 183572 16546 183784 16574
rect 183756 480 183784 16546
rect 185044 6914 185072 31350
rect 184952 6886 185072 6914
rect 184952 480 184980 6886
rect 185596 3806 185624 74190
rect 186332 16574 186360 77182
rect 187700 34332 187752 34338
rect 187700 34274 187752 34280
rect 187712 16574 187740 34274
rect 189552 23050 189580 136983
rect 189644 124001 189672 148310
rect 189736 133657 189764 149058
rect 189722 133648 189778 133657
rect 189722 133583 189778 133592
rect 189630 123992 189686 124001
rect 189630 123927 189686 123936
rect 190472 119649 190500 618258
rect 190552 357468 190604 357474
rect 190552 357410 190604 357416
rect 190564 127129 190592 357410
rect 190736 201544 190788 201550
rect 190736 201486 190788 201492
rect 190644 138032 190696 138038
rect 190644 137974 190696 137980
rect 190656 134609 190684 137974
rect 190642 134600 190698 134609
rect 190642 134535 190698 134544
rect 190644 134496 190696 134502
rect 190644 134438 190696 134444
rect 190550 127120 190606 127129
rect 190550 127055 190606 127064
rect 190458 119640 190514 119649
rect 190458 119575 190514 119584
rect 189724 111852 189776 111858
rect 189724 111794 189776 111800
rect 189736 79558 189764 111794
rect 189724 79552 189776 79558
rect 189724 79494 189776 79500
rect 190656 65822 190684 134438
rect 190748 131617 190776 201486
rect 190920 144220 190972 144226
rect 190920 144162 190972 144168
rect 190828 142928 190880 142934
rect 190828 142870 190880 142876
rect 190734 131608 190790 131617
rect 190734 131543 190790 131552
rect 190840 115161 190868 142870
rect 190932 122641 190960 144162
rect 191010 136096 191066 136105
rect 191010 136031 191066 136040
rect 191024 134502 191052 136031
rect 191012 134496 191064 134502
rect 191012 134438 191064 134444
rect 190918 122632 190974 122641
rect 190918 122567 190974 122576
rect 190826 115152 190882 115161
rect 190826 115087 190882 115096
rect 191116 77790 191144 643078
rect 193864 630692 193916 630698
rect 193864 630634 193916 630640
rect 192484 590708 192536 590714
rect 192484 590650 192536 590656
rect 191840 565888 191892 565894
rect 191840 565830 191892 565836
rect 191852 121145 191880 565830
rect 191932 139392 191984 139398
rect 191932 139334 191984 139340
rect 191944 128625 191972 139334
rect 192024 139324 192076 139330
rect 192024 139266 192076 139272
rect 192036 130121 192064 139266
rect 192022 130112 192078 130121
rect 192022 130047 192078 130056
rect 191930 128616 191986 128625
rect 191930 128551 191986 128560
rect 191838 121136 191894 121145
rect 191838 121071 191894 121080
rect 192208 101788 192260 101794
rect 192208 101730 192260 101736
rect 192220 101697 192248 101730
rect 192206 101688 192262 101697
rect 192206 101623 192262 101632
rect 192208 100428 192260 100434
rect 192208 100370 192260 100376
rect 192220 100201 192248 100370
rect 192206 100192 192262 100201
rect 192206 100127 192262 100136
rect 192208 98864 192260 98870
rect 192208 98806 192260 98812
rect 192220 98705 192248 98806
rect 192206 98696 192262 98705
rect 192206 98631 192262 98640
rect 192496 78606 192524 590650
rect 192576 536852 192628 536858
rect 192576 536794 192628 536800
rect 192484 78600 192536 78606
rect 192484 78542 192536 78548
rect 192588 78538 192616 536794
rect 192668 418192 192720 418198
rect 192668 418134 192720 418140
rect 192680 95713 192708 418134
rect 192760 378208 192812 378214
rect 192760 378150 192812 378156
rect 192666 95704 192722 95713
rect 192666 95639 192722 95648
rect 192666 83736 192722 83745
rect 192666 83671 192722 83680
rect 192576 78532 192628 78538
rect 192576 78474 192628 78480
rect 191104 77784 191156 77790
rect 191104 77726 191156 77732
rect 191840 75608 191892 75614
rect 191840 75550 191892 75556
rect 190644 65816 190696 65822
rect 190644 65758 190696 65764
rect 190460 27328 190512 27334
rect 190460 27270 190512 27276
rect 189540 23044 189592 23050
rect 189540 22986 189592 22992
rect 186332 16546 186912 16574
rect 187712 16546 188568 16574
rect 185584 3800 185636 3806
rect 185584 3742 185636 3748
rect 186136 3188 186188 3194
rect 186136 3130 186188 3136
rect 186148 480 186176 3130
rect 182518 354 182630 480
rect 182192 326 182630 354
rect 181414 -960 181526 326
rect 182518 -960 182630 326
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 186884 354 186912 16546
rect 188540 480 188568 16546
rect 189724 6792 189776 6798
rect 189724 6734 189776 6740
rect 189736 480 189764 6734
rect 187302 354 187414 480
rect 186884 326 187414 354
rect 187302 -960 187414 326
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190472 354 190500 27270
rect 191852 16574 191880 75550
rect 192680 60722 192708 83671
rect 192772 79286 192800 378150
rect 192852 271924 192904 271930
rect 192852 271866 192904 271872
rect 192864 93854 192892 271866
rect 193128 113144 193180 113150
rect 193128 113086 193180 113092
rect 193140 112169 193168 113086
rect 193126 112160 193182 112169
rect 193126 112095 193182 112104
rect 193128 111784 193180 111790
rect 193128 111726 193180 111732
rect 193140 110673 193168 111726
rect 193126 110664 193182 110673
rect 193126 110599 193182 110608
rect 193036 110424 193088 110430
rect 193036 110366 193088 110372
rect 193048 109177 193076 110366
rect 193034 109168 193090 109177
rect 193034 109103 193090 109112
rect 193036 108996 193088 109002
rect 193036 108938 193088 108944
rect 193048 107681 193076 108938
rect 193034 107672 193090 107681
rect 193034 107607 193090 107616
rect 193128 106208 193180 106214
rect 193126 106176 193128 106185
rect 193180 106176 193182 106185
rect 193126 106111 193182 106120
rect 193128 104712 193180 104718
rect 193126 104680 193128 104689
rect 193180 104680 193182 104689
rect 193126 104615 193182 104624
rect 193128 103216 193180 103222
rect 193126 103184 193128 103193
rect 193180 103184 193182 103193
rect 193126 103119 193182 103128
rect 193876 101794 193904 630634
rect 193956 576904 194008 576910
rect 193956 576846 194008 576852
rect 193864 101788 193916 101794
rect 193864 101730 193916 101736
rect 193968 100434 193996 576846
rect 194048 524476 194100 524482
rect 194048 524418 194100 524424
rect 193956 100428 194008 100434
rect 193956 100370 194008 100376
rect 194060 98870 194088 524418
rect 196636 103222 196664 683130
rect 196716 191888 196768 191894
rect 196716 191830 196768 191836
rect 196624 103216 196676 103222
rect 196624 103158 196676 103164
rect 194048 98864 194100 98870
rect 194048 98806 194100 98812
rect 193128 97980 193180 97986
rect 193128 97922 193180 97928
rect 193140 97209 193168 97922
rect 193126 97200 193182 97209
rect 193126 97135 193182 97144
rect 193128 95192 193180 95198
rect 193128 95134 193180 95140
rect 193140 94217 193168 95134
rect 193126 94208 193182 94217
rect 193126 94143 193182 94152
rect 192864 93826 192984 93854
rect 192850 82240 192906 82249
rect 192850 82175 192906 82184
rect 192864 81462 192892 82175
rect 192852 81456 192904 81462
rect 192852 81398 192904 81404
rect 192760 79280 192812 79286
rect 192760 79222 192812 79228
rect 192956 79218 192984 93826
rect 193128 93832 193180 93838
rect 193128 93774 193180 93780
rect 193140 92721 193168 93774
rect 193126 92712 193182 92721
rect 193126 92647 193182 92656
rect 193128 92472 193180 92478
rect 193128 92414 193180 92420
rect 193140 91225 193168 92414
rect 193126 91216 193182 91225
rect 193126 91151 193182 91160
rect 193126 89720 193182 89729
rect 193126 89655 193128 89664
rect 193180 89655 193182 89664
rect 193128 89626 193180 89632
rect 193128 88324 193180 88330
rect 193128 88266 193180 88272
rect 193140 88233 193168 88266
rect 193126 88224 193182 88233
rect 193126 88159 193182 88168
rect 193128 86964 193180 86970
rect 193128 86906 193180 86912
rect 193140 86737 193168 86906
rect 193126 86728 193182 86737
rect 193126 86663 193182 86672
rect 193128 85536 193180 85542
rect 193128 85478 193180 85484
rect 193140 85241 193168 85478
rect 193126 85232 193182 85241
rect 193126 85167 193182 85176
rect 196728 80617 196756 191830
rect 196900 151836 196952 151842
rect 196900 151778 196952 151784
rect 196912 81025 196940 151778
rect 198016 104718 198044 700266
rect 199396 106214 199424 700334
rect 200776 109002 200804 700402
rect 200764 108996 200816 109002
rect 200764 108938 200816 108944
rect 199384 106208 199436 106214
rect 199384 106150 199436 106156
rect 198004 104712 198056 104718
rect 198004 104654 198056 104660
rect 196898 81016 196954 81025
rect 196898 80951 196954 80960
rect 196714 80608 196770 80617
rect 196714 80543 196770 80552
rect 192944 79212 192996 79218
rect 192944 79154 192996 79160
rect 201512 79150 201540 702986
rect 218992 700670 219020 703520
rect 207664 700664 207716 700670
rect 207664 700606 207716 700612
rect 218980 700664 219032 700670
rect 218980 700606 219032 700612
rect 206284 700596 206336 700602
rect 206284 700538 206336 700544
rect 203524 700528 203576 700534
rect 203524 700470 203576 700476
rect 203536 110430 203564 700470
rect 206296 111790 206324 700538
rect 207676 113150 207704 700606
rect 234632 275330 234660 703582
rect 235000 703474 235028 703582
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299492 703582 299980 703610
rect 235184 703474 235212 703520
rect 235000 703446 235212 703474
rect 267660 697610 267688 703520
rect 283852 700602 283880 703520
rect 283840 700596 283892 700602
rect 283840 700538 283892 700544
rect 266360 697604 266412 697610
rect 266360 697546 266412 697552
rect 267648 697604 267700 697610
rect 267648 697546 267700 697552
rect 234620 275324 234672 275330
rect 234620 275266 234672 275272
rect 207664 113144 207716 113150
rect 207664 113086 207716 113092
rect 206284 111784 206336 111790
rect 206284 111726 206336 111732
rect 203524 110424 203576 110430
rect 203524 110366 203576 110372
rect 266372 79665 266400 697546
rect 280804 298172 280856 298178
rect 280804 298114 280856 298120
rect 280816 239426 280844 298114
rect 280804 239420 280856 239426
rect 280804 239362 280856 239368
rect 280804 205692 280856 205698
rect 280804 205634 280856 205640
rect 280816 142866 280844 205634
rect 299492 149734 299520 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429212 703582 429700 703610
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 332520 703050 332548 703520
rect 331220 703044 331272 703050
rect 331220 702986 331272 702992
rect 332508 703044 332560 703050
rect 332508 702986 332560 702992
rect 299480 149728 299532 149734
rect 299480 149670 299532 149676
rect 280804 142860 280856 142866
rect 280804 142802 280856 142808
rect 292580 80300 292632 80306
rect 292580 80242 292632 80248
rect 266358 79656 266414 79665
rect 266358 79591 266414 79600
rect 201500 79144 201552 79150
rect 201500 79086 201552 79092
rect 274640 79076 274692 79082
rect 274640 79018 274692 79024
rect 268384 78260 268436 78266
rect 268384 78202 268436 78208
rect 260102 78024 260158 78033
rect 260102 77959 260158 77968
rect 233238 77208 233294 77217
rect 233238 77143 233294 77152
rect 201500 75540 201552 75546
rect 201500 75482 201552 75488
rect 195980 68536 196032 68542
rect 195980 68478 196032 68484
rect 193220 67176 193272 67182
rect 193220 67118 193272 67124
rect 192668 60716 192720 60722
rect 192668 60658 192720 60664
rect 191852 16546 192064 16574
rect 192036 480 192064 16546
rect 193232 480 193260 67118
rect 194600 34264 194652 34270
rect 194600 34206 194652 34212
rect 193312 27260 193364 27266
rect 193312 27202 193364 27208
rect 193324 16574 193352 27202
rect 194612 16574 194640 34206
rect 195992 16574 196020 68478
rect 200118 62792 200174 62801
rect 200118 62727 200174 62736
rect 198740 34196 198792 34202
rect 198740 34138 198792 34144
rect 193324 16546 194456 16574
rect 194612 16546 195192 16574
rect 195992 16546 196848 16574
rect 194428 480 194456 16546
rect 190798 354 190910 480
rect 190472 326 190910 354
rect 190798 -960 190910 326
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195164 354 195192 16546
rect 196820 480 196848 16546
rect 197912 3324 197964 3330
rect 197912 3266 197964 3272
rect 197924 480 197952 3266
rect 195582 354 195694 480
rect 195164 326 195694 354
rect 195582 -960 195694 326
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 198752 354 198780 34138
rect 200132 16574 200160 62727
rect 200132 16546 200344 16574
rect 200316 480 200344 16546
rect 201512 4146 201540 75482
rect 202144 74180 202196 74186
rect 202144 74122 202196 74128
rect 201590 24440 201646 24449
rect 201590 24375 201646 24384
rect 201500 4140 201552 4146
rect 201500 4082 201552 4088
rect 201604 3482 201632 24375
rect 201512 3454 201632 3482
rect 201512 480 201540 3454
rect 202156 3330 202184 74122
rect 230480 74112 230532 74118
rect 230480 74054 230532 74060
rect 223580 61600 223632 61606
rect 223580 61542 223632 61548
rect 205640 35692 205692 35698
rect 205640 35634 205692 35640
rect 204260 27192 204312 27198
rect 204260 27134 204312 27140
rect 204272 16574 204300 27134
rect 205652 16574 205680 35634
rect 209872 35624 209924 35630
rect 209872 35566 209924 35572
rect 208400 28756 208452 28762
rect 208400 28698 208452 28704
rect 208412 16574 208440 28698
rect 204272 16546 205128 16574
rect 205652 16546 206232 16574
rect 208412 16546 208624 16574
rect 202696 4140 202748 4146
rect 202696 4082 202748 4088
rect 202144 3324 202196 3330
rect 202144 3266 202196 3272
rect 202708 480 202736 4082
rect 203892 3392 203944 3398
rect 203892 3334 203944 3340
rect 203904 480 203932 3334
rect 205100 480 205128 16546
rect 206204 480 206232 16546
rect 207388 4140 207440 4146
rect 207388 4082 207440 4088
rect 207400 480 207428 4082
rect 208596 480 208624 16546
rect 209884 6914 209912 35566
rect 212540 32904 212592 32910
rect 212540 32846 212592 32852
rect 211160 25968 211212 25974
rect 211160 25910 211212 25916
rect 211172 16574 211200 25910
rect 212552 16574 212580 32846
rect 219440 32836 219492 32842
rect 219440 32778 219492 32784
rect 215298 28248 215354 28257
rect 215298 28183 215354 28192
rect 211172 16546 211752 16574
rect 212552 16546 213408 16574
rect 209792 6886 209912 6914
rect 209792 480 209820 6886
rect 210976 4072 211028 4078
rect 210976 4014 211028 4020
rect 210988 480 211016 4014
rect 199078 354 199190 480
rect 198752 326 199190 354
rect 199078 -960 199190 326
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 211724 354 211752 16546
rect 213380 480 213408 16546
rect 214470 3768 214526 3777
rect 214470 3703 214526 3712
rect 214484 480 214512 3703
rect 212142 354 212254 480
rect 211724 326 212254 354
rect 212142 -960 212254 326
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215312 354 215340 28183
rect 216678 18728 216734 18737
rect 216678 18663 216734 18672
rect 216692 16574 216720 18663
rect 219452 16574 219480 32778
rect 222200 28688 222252 28694
rect 222200 28630 222252 28636
rect 222212 16574 222240 28630
rect 216692 16546 216904 16574
rect 219452 16546 220032 16574
rect 222212 16546 222792 16574
rect 216876 480 216904 16546
rect 218058 3632 218114 3641
rect 218058 3567 218114 3576
rect 218072 480 218100 3567
rect 219256 3256 219308 3262
rect 219256 3198 219308 3204
rect 219268 480 219296 3198
rect 215638 354 215750 480
rect 215312 326 215750 354
rect 215638 -960 215750 326
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220004 354 220032 16546
rect 221556 4004 221608 4010
rect 221556 3946 221608 3952
rect 221568 480 221596 3946
rect 222764 480 222792 16546
rect 220422 354 220534 480
rect 220004 326 220534 354
rect 220422 -960 220534 326
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223592 354 223620 61542
rect 226340 49020 226392 49026
rect 226340 48962 226392 48968
rect 225144 3868 225196 3874
rect 225144 3810 225196 3816
rect 225156 480 225184 3810
rect 226352 480 226380 48962
rect 226432 34128 226484 34134
rect 226432 34070 226484 34076
rect 226444 16574 226472 34070
rect 229100 28620 229152 28626
rect 229100 28562 229152 28568
rect 228364 20120 228416 20126
rect 228364 20062 228416 20068
rect 226444 16546 227576 16574
rect 227548 480 227576 16546
rect 228376 3874 228404 20062
rect 229112 16574 229140 28562
rect 230492 16574 230520 74054
rect 233252 16574 233280 77143
rect 240140 77104 240192 77110
rect 240140 77046 240192 77052
rect 253938 77072 253994 77081
rect 237380 32768 237432 32774
rect 237380 32710 237432 32716
rect 235998 29608 236054 29617
rect 235998 29543 236054 29552
rect 236012 16574 236040 29543
rect 237392 16574 237420 32710
rect 229112 16546 229416 16574
rect 230492 16546 231072 16574
rect 233252 16546 233464 16574
rect 236012 16546 236592 16574
rect 237392 16546 237696 16574
rect 228732 6724 228784 6730
rect 228732 6666 228784 6672
rect 228364 3868 228416 3874
rect 228364 3810 228416 3816
rect 228744 480 228772 6666
rect 223918 354 224030 480
rect 223592 326 224030 354
rect 223918 -960 224030 326
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229388 354 229416 16546
rect 231044 480 231072 16546
rect 232226 6080 232282 6089
rect 232226 6015 232282 6024
rect 232240 480 232268 6015
rect 233436 480 233464 16546
rect 235814 6896 235870 6905
rect 235814 6831 235870 6840
rect 234618 5264 234674 5273
rect 234618 5199 234674 5208
rect 234632 480 234660 5199
rect 235828 480 235856 6831
rect 229806 354 229918 480
rect 229388 326 229918 354
rect 229806 -960 229918 326
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236564 354 236592 16546
rect 236982 354 237094 480
rect 236564 326 237094 354
rect 237668 354 237696 16546
rect 239312 6656 239364 6662
rect 239312 6598 239364 6604
rect 239324 480 239352 6598
rect 238086 354 238198 480
rect 237668 326 238198 354
rect 236982 -960 237094 326
rect 238086 -960 238198 326
rect 239282 -960 239394 480
rect 240152 354 240180 77046
rect 253938 77007 253994 77016
rect 251178 73944 251234 73953
rect 251178 73879 251234 73888
rect 241520 34060 241572 34066
rect 241520 34002 241572 34008
rect 241532 16574 241560 34002
rect 242900 29980 242952 29986
rect 242900 29922 242952 29928
rect 241532 16546 241744 16574
rect 241716 480 241744 16546
rect 242912 3398 242940 29922
rect 247040 29912 247092 29918
rect 247040 29854 247092 29860
rect 247052 16574 247080 29854
rect 247052 16546 247632 16574
rect 242992 6588 243044 6594
rect 242992 6530 243044 6536
rect 242900 3392 242952 3398
rect 242900 3334 242952 3340
rect 243004 3210 243032 6530
rect 246396 6520 246448 6526
rect 246396 6462 246448 6468
rect 244096 3392 244148 3398
rect 244096 3334 244148 3340
rect 242912 3182 243032 3210
rect 242912 480 242940 3182
rect 244108 480 244136 3334
rect 245200 3324 245252 3330
rect 245200 3266 245252 3272
rect 245212 480 245240 3266
rect 246408 480 246436 6462
rect 247604 480 247632 16546
rect 248420 13524 248472 13530
rect 248420 13466 248472 13472
rect 240478 354 240590 480
rect 240152 326 240590 354
rect 240478 -960 240590 326
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248432 354 248460 13466
rect 249984 6452 250036 6458
rect 249984 6394 250036 6400
rect 249996 480 250024 6394
rect 251192 4010 251220 73879
rect 253952 16574 253980 77007
rect 259460 74044 259512 74050
rect 259460 73986 259512 73992
rect 255320 35556 255372 35562
rect 255320 35498 255372 35504
rect 255332 16574 255360 35498
rect 253952 16546 254256 16574
rect 255332 16546 255912 16574
rect 251270 7576 251326 7585
rect 251270 7511 251326 7520
rect 251180 4004 251232 4010
rect 251180 3946 251232 3952
rect 251284 3482 251312 7511
rect 253478 6760 253534 6769
rect 253478 6695 253534 6704
rect 252376 4004 252428 4010
rect 252376 3946 252428 3952
rect 251192 3454 251312 3482
rect 251192 480 251220 3454
rect 252388 480 252416 3946
rect 253492 480 253520 6695
rect 248758 354 248870 480
rect 248432 326 248870 354
rect 248758 -960 248870 326
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254228 354 254256 16546
rect 255884 480 255912 16546
rect 256700 15088 256752 15094
rect 256700 15030 256752 15036
rect 254646 354 254758 480
rect 254228 326 254758 354
rect 254646 -960 254758 326
rect 255842 -960 255954 480
rect 256712 354 256740 15030
rect 258264 8832 258316 8838
rect 258264 8774 258316 8780
rect 258276 480 258304 8774
rect 259472 480 259500 73986
rect 260116 20126 260144 77959
rect 260840 77036 260892 77042
rect 260840 76978 260892 76984
rect 260104 20120 260156 20126
rect 260104 20062 260156 20068
rect 260852 16574 260880 76978
rect 267740 76968 267792 76974
rect 267740 76910 267792 76916
rect 266360 73976 266412 73982
rect 266360 73918 266412 73924
rect 264980 29844 265032 29850
rect 264980 29786 265032 29792
rect 260852 16546 261800 16574
rect 260656 6384 260708 6390
rect 260656 6326 260708 6332
rect 260668 480 260696 6326
rect 261772 480 261800 16546
rect 262496 15020 262548 15026
rect 262496 14962 262548 14968
rect 257038 354 257150 480
rect 256712 326 257150 354
rect 257038 -960 257150 326
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262508 354 262536 14962
rect 264152 8900 264204 8906
rect 264152 8842 264204 8848
rect 264164 480 264192 8842
rect 262926 354 263038 480
rect 262508 326 263038 354
rect 262926 -960 263038 326
rect 264122 -960 264234 480
rect 264992 354 265020 29786
rect 266372 16574 266400 73918
rect 267752 16574 267780 76910
rect 268396 20194 268424 78202
rect 273260 73908 273312 73914
rect 273260 73850 273312 73856
rect 271878 30968 271934 30977
rect 271878 30903 271934 30912
rect 269118 20224 269174 20233
rect 268384 20188 268436 20194
rect 269118 20159 269174 20168
rect 268384 20130 268436 20136
rect 269132 16574 269160 20159
rect 271892 16574 271920 30903
rect 266372 16546 266584 16574
rect 267752 16546 268424 16574
rect 269132 16546 270080 16574
rect 271892 16546 272472 16574
rect 266556 480 266584 16546
rect 267740 8764 267792 8770
rect 267740 8706 267792 8712
rect 267752 480 267780 8706
rect 265318 354 265430 480
rect 264992 326 265430 354
rect 265318 -960 265430 326
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268396 354 268424 16546
rect 270052 480 270080 16546
rect 271234 9208 271290 9217
rect 271234 9143 271290 9152
rect 271248 480 271276 9143
rect 272444 480 272472 16546
rect 268814 354 268926 480
rect 268396 326 268926 354
rect 268814 -960 268926 326
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273272 354 273300 73850
rect 274652 16574 274680 79018
rect 289818 76936 289874 76945
rect 289818 76871 289874 76880
rect 287058 73808 287114 73817
rect 287058 73743 287114 73752
rect 277400 61532 277452 61538
rect 277400 61474 277452 61480
rect 276020 27124 276072 27130
rect 276020 27066 276072 27072
rect 274652 16546 274864 16574
rect 274836 480 274864 16546
rect 276032 480 276060 27066
rect 276112 20324 276164 20330
rect 276112 20266 276164 20272
rect 276124 16574 276152 20266
rect 277412 16574 277440 61474
rect 280160 33992 280212 33998
rect 280160 33934 280212 33940
rect 278780 28552 278832 28558
rect 278780 28494 278832 28500
rect 278792 16574 278820 28494
rect 280172 16574 280200 33934
rect 285678 26888 285734 26897
rect 285678 26823 285734 26832
rect 282920 25900 282972 25906
rect 282920 25842 282972 25848
rect 282932 16574 282960 25842
rect 284300 20256 284352 20262
rect 284300 20198 284352 20204
rect 276124 16546 276704 16574
rect 277412 16546 278360 16574
rect 278792 16546 279096 16574
rect 280172 16546 280752 16574
rect 282932 16546 283144 16574
rect 273598 354 273710 480
rect 273272 326 273710 354
rect 273598 -960 273710 326
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 276676 354 276704 16546
rect 278332 480 278360 16546
rect 277094 354 277206 480
rect 276676 326 277206 354
rect 277094 -960 277206 326
rect 278290 -960 278402 480
rect 279068 354 279096 16546
rect 280724 480 280752 16546
rect 281908 9648 281960 9654
rect 281908 9590 281960 9596
rect 281920 480 281948 9590
rect 283116 480 283144 16546
rect 284312 480 284340 20198
rect 285692 16574 285720 26823
rect 287072 16574 287100 73743
rect 285692 16546 286640 16574
rect 287072 16546 287376 16574
rect 285404 9580 285456 9586
rect 285404 9522 285456 9528
rect 285416 480 285444 9522
rect 286612 480 286640 16546
rect 279486 354 279598 480
rect 279068 326 279598 354
rect 279486 -960 279598 326
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287348 354 287376 16546
rect 288990 10432 289046 10441
rect 288990 10367 289046 10376
rect 289004 480 289032 10367
rect 287766 354 287878 480
rect 287348 326 287878 354
rect 287766 -960 287878 326
rect 288962 -960 289074 480
rect 289832 354 289860 76871
rect 291200 33924 291252 33930
rect 291200 33866 291252 33872
rect 291212 16574 291240 33866
rect 291212 16546 291424 16574
rect 291396 480 291424 16546
rect 292592 480 292620 80242
rect 316040 80232 316092 80238
rect 316040 80174 316092 80180
rect 313280 78940 313332 78946
rect 313280 78882 313332 78888
rect 303618 76800 303674 76809
rect 303618 76735 303674 76744
rect 293960 72820 294012 72826
rect 293960 72762 294012 72768
rect 292672 31340 292724 31346
rect 292672 31282 292724 31288
rect 292684 16574 292712 31282
rect 293972 16574 294000 72762
rect 300860 72752 300912 72758
rect 300860 72694 300912 72700
rect 295340 65952 295392 65958
rect 295340 65894 295392 65900
rect 295352 16574 295380 65894
rect 299480 31272 299532 31278
rect 299480 31214 299532 31220
rect 296720 24404 296772 24410
rect 296720 24346 296772 24352
rect 296732 16574 296760 24346
rect 292684 16546 293264 16574
rect 293972 16546 294920 16574
rect 295352 16546 295656 16574
rect 296732 16546 297312 16574
rect 290158 354 290270 480
rect 289832 326 290270 354
rect 290158 -960 290270 326
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293236 354 293264 16546
rect 294892 480 294920 16546
rect 293654 354 293766 480
rect 293236 326 293766 354
rect 293654 -960 293766 326
rect 294850 -960 294962 480
rect 295628 354 295656 16546
rect 297284 480 297312 16546
rect 298100 10736 298152 10742
rect 298100 10678 298152 10684
rect 296046 354 296158 480
rect 295628 326 296158 354
rect 296046 -960 296158 326
rect 297242 -960 297354 480
rect 298112 354 298140 10678
rect 299492 3398 299520 31214
rect 300872 16574 300900 72694
rect 303632 16574 303660 76735
rect 309140 71188 309192 71194
rect 309140 71130 309192 71136
rect 307760 65884 307812 65890
rect 307760 65826 307812 65832
rect 306378 55856 306434 55865
rect 306378 55791 306434 55800
rect 300872 16546 301544 16574
rect 303632 16546 303936 16574
rect 299664 10668 299716 10674
rect 299664 10610 299716 10616
rect 299480 3392 299532 3398
rect 299480 3334 299532 3340
rect 299676 480 299704 10610
rect 300768 3392 300820 3398
rect 300768 3334 300820 3340
rect 300780 480 300808 3334
rect 298438 354 298550 480
rect 298112 326 298550 354
rect 298438 -960 298550 326
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301516 354 301544 16546
rect 303160 10600 303212 10606
rect 303160 10542 303212 10548
rect 303172 480 303200 10542
rect 301934 354 302046 480
rect 301516 326 302046 354
rect 301934 -960 302046 326
rect 303130 -960 303242 480
rect 303908 354 303936 16546
rect 305550 16144 305606 16153
rect 305550 16079 305606 16088
rect 305564 480 305592 16079
rect 304326 354 304438 480
rect 303908 326 304438 354
rect 304326 -960 304438 326
rect 305522 -960 305634 480
rect 306392 354 306420 55791
rect 307772 3398 307800 65826
rect 309152 16574 309180 71130
rect 311900 35488 311952 35494
rect 311900 35430 311952 35436
rect 310520 28484 310572 28490
rect 310520 28426 310572 28432
rect 310532 16574 310560 28426
rect 311912 16574 311940 35430
rect 313292 16574 313320 78882
rect 314660 25832 314712 25838
rect 314660 25774 314712 25780
rect 309152 16546 309824 16574
rect 310532 16546 311480 16574
rect 311912 16546 312216 16574
rect 313292 16546 313872 16574
rect 307942 6624 307998 6633
rect 307942 6559 307998 6568
rect 307760 3392 307812 3398
rect 307760 3334 307812 3340
rect 307956 480 307984 6559
rect 309048 3392 309100 3398
rect 309048 3334 309100 3340
rect 309060 480 309088 3334
rect 306718 354 306830 480
rect 306392 326 306830 354
rect 306718 -960 306830 326
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 309796 354 309824 16546
rect 311452 480 311480 16546
rect 310214 354 310326 480
rect 309796 326 310326 354
rect 310214 -960 310326 326
rect 311410 -960 311522 480
rect 312188 354 312216 16546
rect 313844 480 313872 16546
rect 312606 354 312718 480
rect 312188 326 312718 354
rect 312606 -960 312718 326
rect 313802 -960 313914 480
rect 314672 354 314700 25774
rect 316052 3398 316080 80174
rect 331232 79529 331260 702986
rect 348804 700534 348832 703520
rect 364996 702434 365024 703520
rect 364352 702406 365024 702434
rect 348792 700528 348844 700534
rect 348792 700470 348844 700476
rect 362224 311908 362276 311914
rect 362224 311850 362276 311856
rect 360844 244316 360896 244322
rect 360844 244258 360896 244264
rect 360856 202162 360884 244258
rect 360844 202156 360896 202162
rect 360844 202098 360896 202104
rect 358084 178084 358136 178090
rect 358084 178026 358136 178032
rect 358096 88330 358124 178026
rect 362236 93838 362264 311850
rect 364352 140214 364380 702406
rect 366364 364404 366416 364410
rect 366364 364346 366416 364352
rect 364340 140208 364392 140214
rect 364340 140150 364392 140156
rect 366376 95198 366404 364346
rect 366364 95192 366416 95198
rect 366364 95134 366416 95140
rect 362224 93832 362276 93838
rect 362224 93774 362276 93780
rect 358084 88324 358136 88330
rect 358084 88266 358136 88272
rect 347044 81456 347096 81462
rect 347044 81398 347096 81404
rect 331218 79520 331274 79529
rect 331218 79455 331274 79464
rect 337384 78192 337436 78198
rect 337384 78134 337436 78140
rect 327080 76900 327132 76906
rect 327080 76842 327132 76848
rect 324318 76664 324374 76673
rect 324318 76599 324374 76608
rect 316132 72684 316184 72690
rect 316132 72626 316184 72632
rect 316144 16574 316172 72626
rect 322940 72616 322992 72622
rect 322940 72558 322992 72564
rect 317420 29776 317472 29782
rect 317420 29718 317472 29724
rect 317432 16574 317460 29718
rect 321560 24336 321612 24342
rect 321560 24278 321612 24284
rect 318800 17468 318852 17474
rect 318800 17410 318852 17416
rect 318812 16574 318840 17410
rect 321572 16574 321600 24278
rect 316144 16546 316264 16574
rect 317432 16546 318104 16574
rect 318812 16546 319760 16574
rect 321572 16546 322152 16574
rect 316040 3392 316092 3398
rect 316040 3334 316092 3340
rect 316236 480 316264 16546
rect 317328 3392 317380 3398
rect 317328 3334 317380 3340
rect 317340 480 317368 3334
rect 314998 354 315110 480
rect 314672 326 315110 354
rect 314998 -960 315110 326
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 354 318104 16546
rect 319732 480 319760 16546
rect 320456 12368 320508 12374
rect 320456 12310 320508 12316
rect 318494 354 318606 480
rect 318076 326 318606 354
rect 318494 -960 318606 326
rect 319690 -960 319802 480
rect 320468 354 320496 12310
rect 322124 480 322152 16546
rect 320886 354 320998 480
rect 320468 326 320998 354
rect 320886 -960 320998 326
rect 322082 -960 322194 480
rect 322952 354 322980 72558
rect 324332 3398 324360 76599
rect 327092 16574 327120 76842
rect 328460 76832 328512 76838
rect 328460 76774 328512 76780
rect 328472 16574 328500 76774
rect 333980 58676 334032 58682
rect 333980 58618 334032 58624
rect 333992 16574 334020 58618
rect 327092 16546 328040 16574
rect 328472 16546 328776 16574
rect 333992 16546 334664 16574
rect 324410 12336 324466 12345
rect 324410 12271 324466 12280
rect 326344 12300 326396 12306
rect 324320 3392 324372 3398
rect 324320 3334 324372 3340
rect 324424 480 324452 12271
rect 326344 12242 326396 12248
rect 325608 3392 325660 3398
rect 325608 3334 325660 3340
rect 325620 480 325648 3334
rect 323278 354 323390 480
rect 322952 326 323390 354
rect 323278 -960 323390 326
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326356 354 326384 12242
rect 328012 480 328040 16546
rect 326774 354 326886 480
rect 326356 326 326886 354
rect 326774 -960 326886 326
rect 327970 -960 328082 480
rect 328748 354 328776 16546
rect 330392 12232 330444 12238
rect 330392 12174 330444 12180
rect 330404 480 330432 12174
rect 331220 12164 331272 12170
rect 331220 12106 331272 12112
rect 329166 354 329278 480
rect 328748 326 329278 354
rect 329166 -960 329278 326
rect 330362 -960 330474 480
rect 331232 354 331260 12106
rect 332600 12096 332652 12102
rect 332600 12038 332652 12044
rect 332612 3398 332640 12038
rect 332692 9512 332744 9518
rect 332692 9454 332744 9460
rect 332600 3392 332652 3398
rect 332600 3334 332652 3340
rect 332704 480 332732 9454
rect 333888 3392 333940 3398
rect 333888 3334 333940 3340
rect 333900 480 333928 3334
rect 331558 354 331670 480
rect 331232 326 331670 354
rect 331558 -960 331670 326
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 354 334664 16546
rect 337016 12028 337068 12034
rect 337016 11970 337068 11976
rect 336280 9444 336332 9450
rect 336280 9386 336332 9392
rect 336292 480 336320 9386
rect 335054 354 335166 480
rect 334636 326 335166 354
rect 335054 -960 335166 326
rect 336250 -960 336362 480
rect 337028 354 337056 11970
rect 337396 7886 337424 78134
rect 343640 73840 343692 73846
rect 343640 73782 343692 73788
rect 339500 31204 339552 31210
rect 339500 31146 339552 31152
rect 337384 7880 337436 7886
rect 337384 7822 337436 7828
rect 338670 5128 338726 5137
rect 338670 5063 338726 5072
rect 338684 480 338712 5063
rect 337446 354 337558 480
rect 337028 326 337558 354
rect 337446 -960 337558 326
rect 338642 -960 338754 480
rect 339512 354 339540 31146
rect 343652 16574 343680 73782
rect 346400 55888 346452 55894
rect 346400 55830 346452 55836
rect 346412 16574 346440 55830
rect 347056 20670 347084 81398
rect 374000 80164 374052 80170
rect 374000 80106 374052 80112
rect 362960 79824 363012 79830
rect 362960 79766 363012 79772
rect 349804 78124 349856 78130
rect 349804 78066 349856 78072
rect 347780 72548 347832 72554
rect 347780 72490 347832 72496
rect 347044 20664 347096 20670
rect 347044 20606 347096 20612
rect 347792 16574 347820 72490
rect 343652 16546 344600 16574
rect 346412 16546 346992 16574
rect 347792 16546 348096 16574
rect 340878 13152 340934 13161
rect 340878 13087 340934 13096
rect 340892 3398 340920 13087
rect 340970 12200 341026 12209
rect 340970 12135 341026 12144
rect 340880 3392 340932 3398
rect 340880 3334 340932 3340
rect 340984 480 341012 12135
rect 343362 9072 343418 9081
rect 343362 9007 343418 9016
rect 342168 3392 342220 3398
rect 342168 3334 342220 3340
rect 342180 480 342208 3334
rect 343376 480 343404 9007
rect 344572 480 344600 16546
rect 345296 13456 345348 13462
rect 345296 13398 345348 13404
rect 339838 354 339950 480
rect 339512 326 339950 354
rect 339838 -960 339950 326
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345308 354 345336 13398
rect 346964 480 346992 16546
rect 348068 480 348096 16546
rect 349816 10470 349844 78066
rect 354680 72480 354732 72486
rect 354680 72422 354732 72428
rect 350540 33856 350592 33862
rect 350540 33798 350592 33804
rect 349896 25764 349948 25770
rect 349896 25706 349948 25712
rect 349252 10464 349304 10470
rect 349252 10406 349304 10412
rect 349804 10464 349856 10470
rect 349804 10406 349856 10412
rect 349160 3936 349212 3942
rect 349160 3878 349212 3884
rect 349172 1986 349200 3878
rect 349264 3398 349292 10406
rect 349908 3942 349936 25706
rect 350552 16574 350580 33798
rect 354692 16574 354720 72422
rect 360200 71120 360252 71126
rect 360200 71062 360252 71068
rect 357438 20088 357494 20097
rect 357438 20023 357494 20032
rect 350552 16546 351224 16574
rect 354692 16546 355272 16574
rect 349896 3936 349948 3942
rect 349896 3878 349948 3884
rect 349252 3392 349304 3398
rect 349252 3334 349304 3340
rect 350448 3392 350500 3398
rect 350448 3334 350500 3340
rect 349172 1958 349292 1986
rect 349264 480 349292 1958
rect 350460 480 350488 3334
rect 345726 354 345838 480
rect 345308 326 345838 354
rect 345726 -960 345838 326
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351196 354 351224 16546
rect 352840 13388 352892 13394
rect 352840 13330 352892 13336
rect 352852 480 352880 13330
rect 353576 10532 353628 10538
rect 353576 10474 353628 10480
rect 351614 354 351726 480
rect 351196 326 351726 354
rect 351614 -960 351726 326
rect 352810 -960 352922 480
rect 353588 354 353616 10474
rect 355244 480 355272 16546
rect 356334 14920 356390 14929
rect 356334 14855 356390 14864
rect 356348 480 356376 14855
rect 357452 3398 357480 20023
rect 360212 16574 360240 71062
rect 361580 62892 361632 62898
rect 361580 62834 361632 62840
rect 361592 16574 361620 62834
rect 362972 16574 363000 79766
rect 368480 76764 368532 76770
rect 368480 76706 368532 76712
rect 367100 76696 367152 76702
rect 367100 76638 367152 76644
rect 365720 67108 365772 67114
rect 365720 67050 365772 67056
rect 364340 28416 364392 28422
rect 364340 28358 364392 28364
rect 364352 16574 364380 28358
rect 360212 16546 361160 16574
rect 361592 16546 361896 16574
rect 362972 16546 363552 16574
rect 364352 16546 364656 16574
rect 359462 14784 359518 14793
rect 359462 14719 359518 14728
rect 357530 12064 357586 12073
rect 357530 11999 357586 12008
rect 357440 3392 357492 3398
rect 357440 3334 357492 3340
rect 357544 480 357572 11999
rect 358728 3392 358780 3398
rect 358728 3334 358780 3340
rect 358740 480 358768 3334
rect 354006 354 354118 480
rect 353588 326 354118 354
rect 354006 -960 354118 326
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359476 354 359504 14719
rect 361132 480 361160 16546
rect 359894 354 360006 480
rect 359476 326 360006 354
rect 359894 -960 360006 326
rect 361090 -960 361202 480
rect 361868 354 361896 16546
rect 363524 480 363552 16546
rect 364628 480 364656 16546
rect 365732 1290 365760 67050
rect 367112 16574 367140 76638
rect 368492 16574 368520 76706
rect 372620 28348 372672 28354
rect 372620 28290 372672 28296
rect 371240 26988 371292 26994
rect 371240 26930 371292 26936
rect 367112 16546 367784 16574
rect 368492 16546 369440 16574
rect 365812 11960 365864 11966
rect 365812 11902 365864 11908
rect 365720 1284 365772 1290
rect 365720 1226 365772 1232
rect 365824 480 365852 11902
rect 367008 1284 367060 1290
rect 367008 1226 367060 1232
rect 367020 480 367048 1226
rect 362286 354 362398 480
rect 361868 326 362398 354
rect 362286 -960 362398 326
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 367756 354 367784 16546
rect 369412 480 369440 16546
rect 370136 14952 370188 14958
rect 370136 14894 370188 14900
rect 368174 354 368286 480
rect 367756 326 368286 354
rect 368174 -960 368286 326
rect 369370 -960 369482 480
rect 370148 354 370176 14894
rect 370566 354 370678 480
rect 370148 326 370678 354
rect 371252 354 371280 26930
rect 372632 16574 372660 28290
rect 372632 16546 372936 16574
rect 372908 480 372936 16546
rect 374012 1170 374040 80106
rect 397472 78985 397500 703520
rect 413664 700466 413692 703520
rect 413652 700460 413704 700466
rect 413652 700402 413704 700408
rect 429212 141438 429240 703582
rect 429672 703474 429700 703582
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494072 703582 494652 703610
rect 429856 703474 429884 703520
rect 429672 703446 429884 703474
rect 429200 141432 429252 141438
rect 429200 141374 429252 141380
rect 397458 78976 397514 78985
rect 397458 78911 397514 78920
rect 462332 78849 462360 703520
rect 478524 700398 478552 703520
rect 478512 700392 478564 700398
rect 478512 700334 478564 700340
rect 494072 140146 494100 703582
rect 494624 703474 494652 703582
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 494808 703474 494836 703520
rect 494624 703446 494836 703474
rect 494060 140140 494112 140146
rect 494060 140082 494112 140088
rect 523132 79688 523184 79694
rect 523132 79630 523184 79636
rect 462318 78840 462374 78849
rect 462318 78775 462374 78784
rect 431224 78056 431276 78062
rect 431224 77998 431276 78004
rect 396078 76528 396134 76537
rect 396078 76463 396134 76472
rect 376758 68232 376814 68241
rect 376758 68167 376814 68176
rect 375380 35420 375432 35426
rect 375380 35362 375432 35368
rect 374092 31136 374144 31142
rect 374092 31078 374144 31084
rect 374104 3398 374132 31078
rect 375392 16574 375420 35362
rect 376772 16574 376800 68167
rect 382280 64388 382332 64394
rect 382280 64330 382332 64336
rect 380900 61464 380952 61470
rect 380900 61406 380952 61412
rect 379520 27056 379572 27062
rect 379520 26998 379572 27004
rect 378138 23080 378194 23089
rect 378138 23015 378194 23024
rect 378152 16574 378180 23015
rect 375392 16546 376064 16574
rect 376772 16546 377720 16574
rect 378152 16546 378456 16574
rect 374092 3392 374144 3398
rect 374092 3334 374144 3340
rect 375288 3392 375340 3398
rect 375288 3334 375340 3340
rect 374012 1142 374132 1170
rect 374104 480 374132 1142
rect 375300 480 375328 3334
rect 371670 354 371782 480
rect 371252 326 371782 354
rect 370566 -960 370678 326
rect 371670 -960 371782 326
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376036 354 376064 16546
rect 377692 480 377720 16546
rect 376454 354 376566 480
rect 376036 326 376566 354
rect 376454 -960 376566 326
rect 377650 -960 377762 480
rect 378428 354 378456 16546
rect 378846 354 378958 480
rect 378428 326 378958 354
rect 379532 354 379560 26998
rect 380912 16574 380940 61406
rect 380912 16546 381216 16574
rect 381188 480 381216 16546
rect 382292 3398 382320 64330
rect 390560 51740 390612 51746
rect 390560 51682 390612 51688
rect 384304 16176 384356 16182
rect 384304 16118 384356 16124
rect 382372 9376 382424 9382
rect 382372 9318 382424 9324
rect 382280 3392 382332 3398
rect 382280 3334 382332 3340
rect 382384 480 382412 9318
rect 383568 3392 383620 3398
rect 383568 3334 383620 3340
rect 383580 480 383608 3334
rect 379950 354 380062 480
rect 379532 326 380062 354
rect 378846 -960 378958 326
rect 379950 -960 380062 326
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384316 354 384344 16118
rect 387800 16108 387852 16114
rect 387800 16050 387852 16056
rect 386696 11892 386748 11898
rect 386696 11834 386748 11840
rect 385960 9308 386012 9314
rect 385960 9250 386012 9256
rect 385972 480 386000 9250
rect 384734 354 384846 480
rect 384316 326 384846 354
rect 384734 -960 384846 326
rect 385930 -960 386042 480
rect 386708 354 386736 11834
rect 387126 354 387238 480
rect 386708 326 387238 354
rect 387812 354 387840 16050
rect 389456 9240 389508 9246
rect 389456 9182 389508 9188
rect 389468 480 389496 9182
rect 390572 3398 390600 51682
rect 395342 16008 395398 16017
rect 395342 15943 395398 15952
rect 390652 14884 390704 14890
rect 390652 14826 390704 14832
rect 390560 3392 390612 3398
rect 390560 3334 390612 3340
rect 390664 480 390692 14826
rect 394238 14648 394294 14657
rect 394238 14583 394294 14592
rect 392582 11928 392638 11937
rect 392582 11863 392638 11872
rect 391848 3392 391900 3398
rect 391848 3334 391900 3340
rect 391860 480 391888 3334
rect 388230 354 388342 480
rect 387812 326 388342 354
rect 387126 -960 387238 326
rect 388230 -960 388342 326
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392596 354 392624 11863
rect 394252 480 394280 14583
rect 395356 480 395384 15943
rect 393014 354 393126 480
rect 392596 326 393126 354
rect 393014 -960 393126 326
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396092 354 396120 76463
rect 415400 69896 415452 69902
rect 415400 69838 415452 69844
rect 397460 35352 397512 35358
rect 397460 35294 397512 35300
rect 397472 16574 397500 35294
rect 404360 35284 404412 35290
rect 404360 35226 404412 35232
rect 400220 32632 400272 32638
rect 400220 32574 400272 32580
rect 400232 16574 400260 32574
rect 397472 16546 397776 16574
rect 400232 16546 400904 16574
rect 397748 480 397776 16546
rect 398840 14816 398892 14822
rect 398840 14758 398892 14764
rect 398852 3210 398880 14758
rect 398932 11824 398984 11830
rect 398932 11766 398984 11772
rect 398944 3398 398972 11766
rect 398932 3392 398984 3398
rect 398932 3334 398984 3340
rect 400128 3392 400180 3398
rect 400128 3334 400180 3340
rect 398852 3182 398972 3210
rect 398944 480 398972 3182
rect 400140 480 400168 3334
rect 396510 354 396622 480
rect 396092 326 396622 354
rect 396510 -960 396622 326
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 400876 354 400904 16546
rect 402520 14612 402572 14618
rect 402520 14554 402572 14560
rect 402532 480 402560 14554
rect 403624 13320 403676 13326
rect 403624 13262 403676 13268
rect 403636 480 403664 13262
rect 401294 354 401406 480
rect 400876 326 401406 354
rect 401294 -960 401406 326
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404372 354 404400 35226
rect 411260 25696 411312 25702
rect 411260 25638 411312 25644
rect 407120 19032 407172 19038
rect 407120 18974 407172 18980
rect 405740 17400 405792 17406
rect 405740 17342 405792 17348
rect 405752 16574 405780 17342
rect 405752 16546 406056 16574
rect 406028 480 406056 16546
rect 407132 3398 407160 18974
rect 408498 17776 408554 17785
rect 408498 17711 408554 17720
rect 408512 16574 408540 17711
rect 411272 16574 411300 25638
rect 414018 22944 414074 22953
rect 414018 22879 414074 22888
rect 412638 17640 412694 17649
rect 412638 17575 412694 17584
rect 408512 16546 409184 16574
rect 411272 16546 411944 16574
rect 407212 13252 407264 13258
rect 407212 13194 407264 13200
rect 407120 3392 407172 3398
rect 407120 3334 407172 3340
rect 407224 480 407252 13194
rect 408408 3392 408460 3398
rect 408408 3334 408460 3340
rect 408420 480 408448 3334
rect 404790 354 404902 480
rect 404372 326 404902 354
rect 404790 -960 404902 326
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409156 354 409184 16546
rect 410798 15872 410854 15881
rect 410798 15807 410854 15816
rect 410812 480 410840 15807
rect 411916 480 411944 16546
rect 409574 354 409686 480
rect 409156 326 409686 354
rect 409574 -960 409686 326
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 412652 354 412680 17575
rect 414032 16574 414060 22879
rect 414032 16546 414336 16574
rect 414308 480 414336 16546
rect 415412 3398 415440 69838
rect 419540 64320 419592 64326
rect 419540 64262 419592 64268
rect 416780 29708 416832 29714
rect 416780 29650 416832 29656
rect 415492 21684 415544 21690
rect 415492 21626 415544 21632
rect 415400 3392 415452 3398
rect 415400 3334 415452 3340
rect 415504 480 415532 21626
rect 416792 16574 416820 29650
rect 418160 24268 418212 24274
rect 418160 24210 418212 24216
rect 418172 16574 418200 24210
rect 419552 16574 419580 64262
rect 423680 64252 423732 64258
rect 423680 64194 423732 64200
rect 422300 35216 422352 35222
rect 422300 35158 422352 35164
rect 422312 16574 422340 35158
rect 416792 16546 417464 16574
rect 418172 16546 418568 16574
rect 419552 16546 420224 16574
rect 422312 16546 422616 16574
rect 416688 3392 416740 3398
rect 416688 3334 416740 3340
rect 416700 480 416728 3334
rect 413070 354 413182 480
rect 412652 326 413182 354
rect 413070 -960 413182 326
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417436 354 417464 16546
rect 417854 354 417966 480
rect 417436 326 417966 354
rect 418540 354 418568 16546
rect 420196 480 420224 16546
rect 420920 14748 420972 14754
rect 420920 14690 420972 14696
rect 418958 354 419070 480
rect 418540 326 419070 354
rect 417854 -960 417966 326
rect 418958 -960 419070 326
rect 420154 -960 420266 480
rect 420932 354 420960 14690
rect 422588 480 422616 16546
rect 423692 3210 423720 64194
rect 429198 36544 429254 36553
rect 429198 36479 429254 36488
rect 423772 32564 423824 32570
rect 423772 32506 423824 32512
rect 423784 3398 423812 32506
rect 426440 18964 426492 18970
rect 426440 18906 426492 18912
rect 426452 16574 426480 18906
rect 426452 16546 426848 16574
rect 426164 7812 426216 7818
rect 426164 7754 426216 7760
rect 423772 3392 423824 3398
rect 423772 3334 423824 3340
rect 424968 3392 425020 3398
rect 424968 3334 425020 3340
rect 423692 3182 423812 3210
rect 423784 480 423812 3182
rect 424980 480 425008 3334
rect 426176 480 426204 7754
rect 421350 354 421462 480
rect 420932 326 421462 354
rect 421350 -960 421462 326
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 426820 354 426848 16546
rect 428464 14680 428516 14686
rect 428464 14622 428516 14628
rect 428476 480 428504 14622
rect 427238 354 427350 480
rect 426820 326 427350 354
rect 427238 -960 427350 326
rect 428434 -960 428546 480
rect 429212 354 429240 36479
rect 430578 18592 430634 18601
rect 430578 18527 430634 18536
rect 430592 16574 430620 18527
rect 430592 16546 430896 16574
rect 430868 480 430896 16546
rect 431236 5166 431264 77998
rect 489920 77988 489972 77994
rect 489920 77930 489972 77936
rect 480258 77888 480314 77897
rect 480258 77823 480314 77832
rect 431958 75440 432014 75449
rect 431958 75375 432014 75384
rect 431224 5160 431276 5166
rect 431224 5102 431276 5108
rect 431972 1170 432000 75375
rect 451280 69828 451332 69834
rect 451280 69770 451332 69776
rect 433340 68468 433392 68474
rect 433340 68410 433392 68416
rect 432052 44872 432104 44878
rect 432052 44814 432104 44820
rect 432064 3398 432092 44814
rect 433352 16574 433380 68410
rect 437480 65748 437532 65754
rect 437480 65690 437532 65696
rect 434720 32496 434772 32502
rect 434720 32438 434772 32444
rect 434732 16574 434760 32438
rect 433352 16546 434024 16574
rect 434732 16546 435128 16574
rect 432052 3392 432104 3398
rect 432052 3334 432104 3340
rect 433248 3392 433300 3398
rect 433248 3334 433300 3340
rect 431972 1142 432092 1170
rect 432064 480 432092 1142
rect 433260 480 433288 3334
rect 429630 354 429742 480
rect 429212 326 429742 354
rect 429630 -960 429742 326
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 433996 354 434024 16546
rect 434414 354 434526 480
rect 433996 326 434526 354
rect 435100 354 435128 16546
rect 436744 9172 436796 9178
rect 436744 9114 436796 9120
rect 436756 480 436784 9114
rect 435518 354 435630 480
rect 435100 326 435630 354
rect 434414 -960 434526 326
rect 435518 -960 435630 326
rect 436714 -960 436826 480
rect 437492 354 437520 65690
rect 441620 33788 441672 33794
rect 441620 33730 441672 33736
rect 438860 32428 438912 32434
rect 438860 32370 438912 32376
rect 438872 16574 438900 32370
rect 440240 18896 440292 18902
rect 440240 18838 440292 18844
rect 438872 16546 439176 16574
rect 439148 480 439176 16546
rect 440252 610 440280 18838
rect 441632 16574 441660 33730
rect 444378 19952 444434 19961
rect 444378 19887 444434 19896
rect 444392 16574 444420 19887
rect 451292 16574 451320 69770
rect 456800 68400 456852 68406
rect 456800 68342 456852 68348
rect 441632 16546 442672 16574
rect 444392 16546 445064 16574
rect 451292 16546 451688 16574
rect 440332 10396 440384 10402
rect 440332 10338 440384 10344
rect 440240 604 440292 610
rect 440240 546 440292 552
rect 440344 480 440372 10338
rect 441528 604 441580 610
rect 441528 546 441580 552
rect 441540 480 441568 546
rect 442644 480 442672 16546
rect 443828 5092 443880 5098
rect 443828 5034 443880 5040
rect 443840 480 443868 5034
rect 445036 480 445064 16546
rect 447416 13184 447468 13190
rect 447416 13126 447468 13132
rect 446218 4992 446274 5001
rect 446218 4927 446274 4936
rect 446232 480 446260 4927
rect 447428 480 447456 13126
rect 448518 11792 448574 11801
rect 448518 11727 448574 11736
rect 448532 3330 448560 11727
rect 448610 6488 448666 6497
rect 448610 6423 448666 6432
rect 448520 3324 448572 3330
rect 448520 3266 448572 3272
rect 448624 480 448652 6423
rect 450912 6316 450964 6322
rect 450912 6258 450964 6264
rect 449808 3324 449860 3330
rect 449808 3266 449860 3272
rect 449820 480 449848 3266
rect 450924 480 450952 6258
rect 437910 354 438022 480
rect 437492 326 438022 354
rect 437910 -960 438022 326
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 451660 354 451688 16546
rect 454040 14544 454092 14550
rect 454040 14486 454092 14492
rect 453304 9104 453356 9110
rect 453304 9046 453356 9052
rect 453316 480 453344 9046
rect 452078 354 452190 480
rect 451660 326 452190 354
rect 452078 -960 452190 326
rect 453274 -960 453386 480
rect 454052 354 454080 14486
rect 455696 7744 455748 7750
rect 455696 7686 455748 7692
rect 455708 480 455736 7686
rect 456812 3398 456840 68342
rect 473360 67040 473412 67046
rect 473360 66982 473412 66988
rect 467840 20188 467892 20194
rect 467840 20130 467892 20136
rect 460940 20120 460992 20126
rect 460940 20062 460992 20068
rect 460952 16574 460980 20062
rect 462320 20052 462372 20058
rect 462320 19994 462372 20000
rect 460952 16546 461624 16574
rect 456892 10328 456944 10334
rect 456892 10270 456944 10276
rect 456800 3392 456852 3398
rect 456800 3334 456852 3340
rect 456904 480 456932 10270
rect 459192 9036 459244 9042
rect 459192 8978 459244 8984
rect 458088 3392 458140 3398
rect 458088 3334 458140 3340
rect 458100 480 458128 3334
rect 459204 480 459232 8978
rect 460388 6248 460440 6254
rect 460388 6190 460440 6196
rect 460400 480 460428 6190
rect 461596 480 461624 16546
rect 454470 354 454582 480
rect 454052 326 454582 354
rect 454470 -960 454582 326
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462332 354 462360 19994
rect 466458 17504 466514 17513
rect 466458 17439 466514 17448
rect 466472 16574 466500 17439
rect 467852 16574 467880 20130
rect 466472 16546 467512 16574
rect 467852 16546 468248 16574
rect 463974 14512 464030 14521
rect 463974 14447 464030 14456
rect 465724 14476 465776 14482
rect 463988 480 464016 14447
rect 465724 14418 465776 14424
rect 465736 3738 465764 14418
rect 466274 8936 466330 8945
rect 466274 8871 466330 8880
rect 465172 3732 465224 3738
rect 465172 3674 465224 3680
rect 465724 3732 465776 3738
rect 465724 3674 465776 3680
rect 465184 480 465212 3674
rect 466288 480 466316 8871
rect 467484 480 467512 16546
rect 462750 354 462862 480
rect 462332 326 462862 354
rect 462750 -960 462862 326
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468220 354 468248 16546
rect 469956 7676 470008 7682
rect 469956 7618 470008 7624
rect 469968 3874 469996 7618
rect 471060 7608 471112 7614
rect 471060 7550 471112 7556
rect 469864 3868 469916 3874
rect 469864 3810 469916 3816
rect 469956 3868 470008 3874
rect 469956 3810 470008 3816
rect 469876 480 469904 3810
rect 471072 480 471100 7550
rect 473372 6914 473400 66982
rect 473452 25628 473504 25634
rect 473452 25570 473504 25576
rect 473464 16574 473492 25570
rect 476120 21616 476172 21622
rect 476120 21558 476172 21564
rect 476132 16574 476160 21558
rect 480272 16574 480300 77823
rect 485780 76628 485832 76634
rect 485780 76570 485832 76576
rect 481638 75304 481694 75313
rect 481638 75239 481694 75248
rect 473464 16546 474136 16574
rect 476132 16546 476528 16574
rect 480272 16546 480576 16574
rect 473372 6886 473492 6914
rect 472256 3800 472308 3806
rect 472256 3742 472308 3748
rect 472268 480 472296 3742
rect 473464 480 473492 6886
rect 468638 354 468750 480
rect 468220 326 468750 354
rect 468638 -960 468750 326
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474108 354 474136 16546
rect 475752 5160 475804 5166
rect 475752 5102 475804 5108
rect 475764 480 475792 5102
rect 474526 354 474638 480
rect 474108 326 474638 354
rect 474526 -960 474638 326
rect 475722 -960 475834 480
rect 476500 354 476528 16546
rect 478144 16040 478196 16046
rect 478144 15982 478196 15988
rect 478156 480 478184 15982
rect 478880 15972 478932 15978
rect 478880 15914 478932 15920
rect 476918 354 477030 480
rect 476500 326 477030 354
rect 476918 -960 477030 326
rect 478114 -960 478226 480
rect 478892 354 478920 15914
rect 480548 480 480576 16546
rect 481652 3398 481680 75239
rect 483018 64288 483074 64297
rect 483018 64223 483074 64232
rect 483032 16574 483060 64223
rect 485792 16574 485820 76570
rect 487160 71052 487212 71058
rect 487160 70994 487212 71000
rect 483032 16546 484072 16574
rect 485792 16546 486464 16574
rect 481730 10296 481786 10305
rect 481730 10231 481786 10240
rect 481640 3392 481692 3398
rect 481640 3334 481692 3340
rect 481744 480 481772 10231
rect 482468 3392 482520 3398
rect 482468 3334 482520 3340
rect 479310 354 479422 480
rect 478892 326 479422 354
rect 479310 -960 479422 326
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482480 354 482508 3334
rect 484044 480 484072 16546
rect 484766 13016 484822 13025
rect 484766 12951 484822 12960
rect 482806 354 482918 480
rect 482480 326 482918 354
rect 482806 -960 482918 326
rect 484002 -960 484114 480
rect 484780 354 484808 12951
rect 486436 480 486464 16546
rect 485198 354 485310 480
rect 484780 326 485310 354
rect 485198 -960 485310 326
rect 486394 -960 486506 480
rect 487172 354 487200 70994
rect 488540 62824 488592 62830
rect 488540 62766 488592 62772
rect 488552 16574 488580 62766
rect 488552 16546 488856 16574
rect 488828 480 488856 16546
rect 489932 3398 489960 77930
rect 499580 75472 499632 75478
rect 499580 75414 499632 75420
rect 498200 69760 498252 69766
rect 498200 69702 498252 69708
rect 496820 31068 496872 31074
rect 496820 31010 496872 31016
rect 495440 21548 495492 21554
rect 495440 21490 495492 21496
rect 492680 17332 492732 17338
rect 492680 17274 492732 17280
rect 492692 16574 492720 17274
rect 492692 16546 493088 16574
rect 490012 13116 490064 13122
rect 490012 13058 490064 13064
rect 489920 3392 489972 3398
rect 489920 3334 489972 3340
rect 490024 3210 490052 13058
rect 492312 11756 492364 11762
rect 492312 11698 492364 11704
rect 490748 3392 490800 3398
rect 490748 3334 490800 3340
rect 489932 3182 490052 3210
rect 489932 480 489960 3182
rect 487590 354 487702 480
rect 487172 326 487702 354
rect 487590 -960 487702 326
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 490760 354 490788 3334
rect 492324 480 492352 11698
rect 491086 354 491198 480
rect 490760 326 491198 354
rect 491086 -960 491198 326
rect 492282 -960 492394 480
rect 493060 354 493088 16546
rect 494704 3664 494756 3670
rect 494704 3606 494756 3612
rect 494716 480 494744 3606
rect 493478 354 493590 480
rect 493060 326 493590 354
rect 493478 -960 493590 326
rect 494674 -960 494786 480
rect 495452 354 495480 21490
rect 496832 16574 496860 31010
rect 496832 16546 497136 16574
rect 497108 480 497136 16546
rect 498212 480 498240 69702
rect 498292 21480 498344 21486
rect 498292 21422 498344 21428
rect 498304 16574 498332 21422
rect 499592 16574 499620 75414
rect 506480 75404 506532 75410
rect 506480 75346 506532 75352
rect 502338 22808 502394 22817
rect 502338 22743 502394 22752
rect 502352 16574 502380 22743
rect 498304 16546 498976 16574
rect 499592 16546 500632 16574
rect 502352 16546 503024 16574
rect 495870 354 495982 480
rect 495452 326 495982 354
rect 495870 -960 495982 326
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 498948 354 498976 16546
rect 500604 480 500632 16546
rect 501788 3528 501840 3534
rect 501788 3470 501840 3476
rect 501800 480 501828 3470
rect 502996 480 503024 16546
rect 504180 3868 504232 3874
rect 504180 3810 504232 3816
rect 504192 480 504220 3810
rect 505376 3596 505428 3602
rect 505376 3538 505428 3544
rect 505388 480 505416 3538
rect 506492 3534 506520 75346
rect 514760 75336 514812 75342
rect 514760 75278 514812 75284
rect 512000 66972 512052 66978
rect 512000 66914 512052 66920
rect 510620 65680 510672 65686
rect 510620 65622 510672 65628
rect 506572 60104 506624 60110
rect 506572 60046 506624 60052
rect 506480 3528 506532 3534
rect 506480 3470 506532 3476
rect 506584 3346 506612 60046
rect 509240 19984 509292 19990
rect 509240 19926 509292 19932
rect 509252 16574 509280 19926
rect 510632 16574 510660 65622
rect 509252 16546 509648 16574
rect 510632 16546 511304 16574
rect 508872 5024 508924 5030
rect 508872 4966 508924 4972
rect 507308 3528 507360 3534
rect 507308 3470 507360 3476
rect 506492 3318 506612 3346
rect 506492 480 506520 3318
rect 499366 354 499478 480
rect 498948 326 499478 354
rect 499366 -960 499478 326
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507320 354 507348 3470
rect 508884 480 508912 4966
rect 507646 354 507758 480
rect 507320 326 507758 354
rect 507646 -960 507758 326
rect 508842 -960 508954 480
rect 509620 354 509648 16546
rect 511276 480 511304 16546
rect 510038 354 510150 480
rect 509620 326 510150 354
rect 510038 -960 510150 326
rect 511234 -960 511346 480
rect 512012 354 512040 66914
rect 513380 22976 513432 22982
rect 513380 22918 513432 22924
rect 512430 354 512542 480
rect 512012 326 512542 354
rect 513392 354 513420 22918
rect 514772 480 514800 75278
rect 521660 75268 521712 75274
rect 521660 75210 521712 75216
rect 514852 68332 514904 68338
rect 514852 68274 514904 68280
rect 514864 16574 514892 68274
rect 518898 61432 518954 61441
rect 518898 61367 518954 61376
rect 517518 17368 517574 17377
rect 517518 17303 517574 17312
rect 517532 16574 517560 17303
rect 518912 16574 518940 61367
rect 520278 22672 520334 22681
rect 520278 22607 520334 22616
rect 514864 16546 515536 16574
rect 517532 16546 517928 16574
rect 518912 16546 519584 16574
rect 513534 354 513646 480
rect 513392 326 513646 354
rect 512430 -960 512542 326
rect 513534 -960 513646 326
rect 514730 -960 514842 480
rect 515508 354 515536 16546
rect 517150 11656 517206 11665
rect 517150 11591 517206 11600
rect 517164 480 517192 11591
rect 515926 354 516038 480
rect 515508 326 516038 354
rect 515926 -960 516038 326
rect 517122 -960 517234 480
rect 517900 354 517928 16546
rect 519556 480 519584 16546
rect 518318 354 518430 480
rect 517900 326 518430 354
rect 518318 -960 518430 326
rect 519514 -960 519626 480
rect 520292 354 520320 22607
rect 520710 354 520822 480
rect 520292 326 520822 354
rect 521672 354 521700 75210
rect 523144 16574 523172 79630
rect 527192 79354 527220 703520
rect 543476 700330 543504 703520
rect 559668 702434 559696 703520
rect 558932 702406 559696 702434
rect 543464 700324 543516 700330
rect 543464 700266 543516 700272
rect 531964 258120 532016 258126
rect 531964 258062 532016 258068
rect 531976 92478 532004 258062
rect 532056 218068 532108 218074
rect 532056 218010 532108 218016
rect 531964 92472 532016 92478
rect 531964 92414 532016 92420
rect 532068 89690 532096 218010
rect 558932 140078 558960 702406
rect 580262 697232 580318 697241
rect 580262 697167 580318 697176
rect 579618 683904 579674 683913
rect 579618 683839 579674 683848
rect 579632 683194 579660 683839
rect 579620 683188 579672 683194
rect 579620 683130 579672 683136
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 579986 630864 580042 630873
rect 579986 630799 580042 630808
rect 580000 630698 580028 630799
rect 579988 630692 580040 630698
rect 579988 630634 580040 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 580170 591016 580226 591025
rect 580170 590951 580226 590960
rect 580184 590714 580212 590951
rect 580172 590708 580224 590714
rect 580172 590650 580224 590656
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 580170 564360 580226 564369
rect 580170 564295 580226 564304
rect 580184 563106 580212 564295
rect 580172 563100 580224 563106
rect 580172 563042 580224 563048
rect 579894 537840 579950 537849
rect 579894 537775 579950 537784
rect 579908 536858 579936 537775
rect 579896 536852 579948 536858
rect 579896 536794 579948 536800
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 579618 458144 579674 458153
rect 579618 458079 579674 458088
rect 579632 456822 579660 458079
rect 579620 456816 579672 456822
rect 579620 456758 579672 456764
rect 579710 418296 579766 418305
rect 579710 418231 579766 418240
rect 579724 418198 579752 418231
rect 579712 418192 579764 418198
rect 579712 418134 579764 418140
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580184 404394 580212 404903
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580184 378214 580212 378383
rect 580172 378208 580224 378214
rect 580172 378150 580224 378156
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 580184 364410 580212 365055
rect 580172 364404 580224 364410
rect 580172 364346 580224 364352
rect 580172 351960 580224 351966
rect 580170 351928 580172 351937
rect 580224 351928 580226 351937
rect 580170 351863 580226 351872
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 580184 311914 580212 312015
rect 580172 311908 580224 311914
rect 580172 311850 580224 311856
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 580184 298178 580212 298687
rect 580172 298172 580224 298178
rect 580172 298114 580224 298120
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 580184 271930 580212 272167
rect 580172 271924 580224 271930
rect 580172 271866 580224 271872
rect 579618 258904 579674 258913
rect 579618 258839 579674 258848
rect 579632 258126 579660 258839
rect 579620 258120 579672 258126
rect 579620 258062 579672 258068
rect 580170 245576 580226 245585
rect 580170 245511 580226 245520
rect 580184 244322 580212 245511
rect 580172 244316 580224 244322
rect 580172 244258 580224 244264
rect 580170 219056 580226 219065
rect 580170 218991 580226 219000
rect 580184 218074 580212 218991
rect 580172 218068 580224 218074
rect 580172 218010 580224 218016
rect 580170 205728 580226 205737
rect 580170 205663 580172 205672
rect 580224 205663 580226 205672
rect 580172 205634 580224 205640
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 580184 191894 580212 192471
rect 580172 191888 580224 191894
rect 580172 191830 580224 191836
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580184 178090 580212 179143
rect 580172 178084 580224 178090
rect 580172 178026 580224 178032
rect 579618 165880 579674 165889
rect 579618 165815 579674 165824
rect 579632 165646 579660 165815
rect 579620 165640 579672 165646
rect 579620 165582 579672 165588
rect 579986 152688 580042 152697
rect 579986 152623 580042 152632
rect 580000 151842 580028 152623
rect 579988 151836 580040 151842
rect 579988 151778 580040 151784
rect 558920 140072 558972 140078
rect 558920 140014 558972 140020
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 580078 112840 580134 112849
rect 580078 112775 580134 112784
rect 580092 111858 580120 112775
rect 580080 111852 580132 111858
rect 580080 111794 580132 111800
rect 532056 89684 532108 89690
rect 532056 89626 532108 89632
rect 579986 86184 580042 86193
rect 579986 86119 580042 86128
rect 580000 80986 580028 86119
rect 580184 81161 580212 125967
rect 580170 81152 580226 81161
rect 580170 81087 580226 81096
rect 579988 80980 580040 80986
rect 579988 80922 580040 80928
rect 547972 80096 548024 80102
rect 547972 80038 548024 80044
rect 527180 79348 527232 79354
rect 527180 79290 527232 79296
rect 542360 76560 542412 76566
rect 542360 76502 542412 76508
rect 535458 75168 535514 75177
rect 535458 75103 535514 75112
rect 529940 66904 529992 66910
rect 529940 66846 529992 66852
rect 525800 61396 525852 61402
rect 525800 61338 525852 61344
rect 525812 16574 525840 61338
rect 528560 22908 528612 22914
rect 528560 22850 528612 22856
rect 523144 16546 523816 16574
rect 525812 16546 526208 16574
rect 523040 3460 523092 3466
rect 523040 3402 523092 3408
rect 523052 480 523080 3402
rect 521814 354 521926 480
rect 521672 326 521926 354
rect 520710 -960 520822 326
rect 521814 -960 521926 326
rect 523010 -960 523122 480
rect 523788 354 523816 16546
rect 525432 8968 525484 8974
rect 525432 8910 525484 8916
rect 525444 480 525472 8910
rect 524206 354 524318 480
rect 523788 326 524318 354
rect 524206 -960 524318 326
rect 525402 -960 525514 480
rect 526180 354 526208 16546
rect 527824 15904 527876 15910
rect 527824 15846 527876 15852
rect 527836 480 527864 15846
rect 526598 354 526710 480
rect 526180 326 526710 354
rect 526598 -960 526710 326
rect 527794 -960 527906 480
rect 528572 354 528600 22850
rect 528990 354 529102 480
rect 528572 326 529102 354
rect 529952 354 529980 66846
rect 534078 24304 534134 24313
rect 534078 24239 534134 24248
rect 531320 22840 531372 22846
rect 531320 22782 531372 22788
rect 531332 3534 531360 22782
rect 531412 17264 531464 17270
rect 531412 17206 531464 17212
rect 531320 3528 531372 3534
rect 531320 3470 531372 3476
rect 531424 3346 531452 17206
rect 534092 16574 534120 24239
rect 535472 16574 535500 75103
rect 536838 65512 536894 65521
rect 536838 65447 536894 65456
rect 536852 16574 536880 65447
rect 539600 60036 539652 60042
rect 539600 59978 539652 59984
rect 538218 24168 538274 24177
rect 538218 24103 538274 24112
rect 534092 16546 534488 16574
rect 535472 16546 536144 16574
rect 536852 16546 537248 16574
rect 533712 4956 533764 4962
rect 533712 4898 533764 4904
rect 532148 3528 532200 3534
rect 532148 3470 532200 3476
rect 531332 3318 531452 3346
rect 531332 480 531360 3318
rect 530094 354 530206 480
rect 529952 326 530206 354
rect 528990 -960 529102 326
rect 530094 -960 530206 326
rect 531290 -960 531402 480
rect 532160 354 532188 3470
rect 533724 480 533752 4898
rect 532486 354 532598 480
rect 532160 326 532598 354
rect 532486 -960 532598 326
rect 533682 -960 533794 480
rect 534460 354 534488 16546
rect 536116 480 536144 16546
rect 537220 480 537248 16546
rect 534878 354 534990 480
rect 534460 326 534990 354
rect 534878 -960 534990 326
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538232 354 538260 24103
rect 539612 3534 539640 59978
rect 539692 28280 539744 28286
rect 539692 28222 539744 28228
rect 539600 3528 539652 3534
rect 539600 3470 539652 3476
rect 539704 3346 539732 28222
rect 540980 24200 541032 24206
rect 540980 24142 541032 24148
rect 540992 16574 541020 24142
rect 542372 16574 542400 76502
rect 546500 25560 546552 25566
rect 546500 25502 546552 25508
rect 540992 16546 542032 16574
rect 542372 16546 542768 16574
rect 540428 3528 540480 3534
rect 540428 3470 540480 3476
rect 539612 3318 539732 3346
rect 539612 480 539640 3318
rect 538374 354 538486 480
rect 538232 326 538486 354
rect 538374 -960 538486 326
rect 539570 -960 539682 480
rect 540440 354 540468 3470
rect 542004 480 542032 16546
rect 540766 354 540878 480
rect 540440 326 540878 354
rect 540766 -960 540878 326
rect 541962 -960 542074 480
rect 542740 354 542768 16546
rect 545488 3936 545540 3942
rect 545488 3878 545540 3884
rect 544382 3496 544438 3505
rect 544382 3431 544438 3440
rect 544396 480 544424 3431
rect 545500 480 545528 3878
rect 543158 354 543270 480
rect 542740 326 543270 354
rect 543158 -960 543270 326
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546512 354 546540 25502
rect 547984 6914 548012 80038
rect 580276 79393 580304 697167
rect 580354 484664 580410 484673
rect 580354 484599 580410 484608
rect 580262 79384 580318 79393
rect 580262 79319 580318 79328
rect 580368 77858 580396 484599
rect 580446 471472 580502 471481
rect 580446 471407 580502 471416
rect 580460 97986 580488 471407
rect 580538 431624 580594 431633
rect 580538 431559 580594 431568
rect 580448 97980 580500 97986
rect 580448 97922 580500 97928
rect 580552 78713 580580 431559
rect 580630 325272 580686 325281
rect 580630 325207 580686 325216
rect 580644 80753 580672 325207
rect 580814 232384 580870 232393
rect 580814 232319 580870 232328
rect 580722 139360 580778 139369
rect 580722 139295 580778 139304
rect 580736 86970 580764 139295
rect 580724 86964 580776 86970
rect 580724 86906 580776 86912
rect 580828 80889 580856 232319
rect 580906 99512 580962 99521
rect 580906 99447 580962 99456
rect 580920 85542 580948 99447
rect 580908 85536 580960 85542
rect 580908 85478 580960 85484
rect 580814 80880 580870 80889
rect 580814 80815 580870 80824
rect 580630 80744 580686 80753
rect 580630 80679 580686 80688
rect 580538 78704 580594 78713
rect 580538 78639 580594 78648
rect 580356 77852 580408 77858
rect 580356 77794 580408 77800
rect 549260 75200 549312 75206
rect 549260 75142 549312 75148
rect 549272 16574 549300 75142
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 571338 71088 571394 71097
rect 571338 71023 571394 71032
rect 561680 69692 561732 69698
rect 561680 69634 561732 69640
rect 552020 64184 552072 64190
rect 552020 64126 552072 64132
rect 554778 64152 554834 64161
rect 552032 16574 552060 64126
rect 554778 64087 554834 64096
rect 553400 18828 553452 18834
rect 553400 18770 553452 18776
rect 553412 16574 553440 18770
rect 549272 16546 550312 16574
rect 552032 16546 552704 16574
rect 553412 16546 553808 16574
rect 547892 6886 548012 6914
rect 547892 480 547920 6886
rect 549076 3732 549128 3738
rect 549076 3674 549128 3680
rect 549088 480 549116 3674
rect 550284 480 550312 16546
rect 551468 4888 551520 4894
rect 551468 4830 551520 4836
rect 551480 480 551508 4830
rect 552676 480 552704 16546
rect 553780 480 553808 16546
rect 546654 354 546766 480
rect 546512 326 546766 354
rect 546654 -960 546766 326
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554792 354 554820 64087
rect 556158 46200 556214 46209
rect 556158 46135 556214 46144
rect 556172 480 556200 46135
rect 556252 18760 556304 18766
rect 556252 18702 556304 18708
rect 556264 16574 556292 18702
rect 558920 18692 558972 18698
rect 558920 18634 558972 18640
rect 558932 16574 558960 18634
rect 560300 18624 560352 18630
rect 560300 18566 560352 18572
rect 560312 16574 560340 18566
rect 561692 16574 561720 69634
rect 564440 65612 564492 65618
rect 564440 65554 564492 65560
rect 563060 21412 563112 21418
rect 563060 21354 563112 21360
rect 556264 16546 556936 16574
rect 558932 16546 559328 16574
rect 560312 16546 560432 16574
rect 561692 16546 562088 16574
rect 554934 354 555046 480
rect 554792 326 555046 354
rect 554934 -960 555046 326
rect 556130 -960 556242 480
rect 556908 354 556936 16546
rect 558550 3360 558606 3369
rect 558550 3295 558606 3304
rect 558564 480 558592 3295
rect 557326 354 557438 480
rect 556908 326 557438 354
rect 557326 -960 557438 326
rect 558522 -960 558634 480
rect 559300 354 559328 16546
rect 559718 354 559830 480
rect 559300 326 559830 354
rect 560404 354 560432 16546
rect 562060 480 562088 16546
rect 560822 354 560934 480
rect 560404 326 560934 354
rect 559718 -960 559830 326
rect 560822 -960 560934 326
rect 562018 -960 562130 480
rect 563072 354 563100 21354
rect 564452 3534 564480 65554
rect 568580 65544 568632 65550
rect 568580 65486 568632 65492
rect 564532 29640 564584 29646
rect 564532 29582 564584 29588
rect 564440 3528 564492 3534
rect 564440 3470 564492 3476
rect 564544 3346 564572 29582
rect 567200 24132 567252 24138
rect 567200 24074 567252 24080
rect 567212 16574 567240 24074
rect 568592 16574 568620 65486
rect 567212 16546 567608 16574
rect 568592 16546 568712 16574
rect 566832 4820 566884 4826
rect 566832 4762 566884 4768
rect 565268 3528 565320 3534
rect 565268 3470 565320 3476
rect 564452 3318 564572 3346
rect 564452 480 564480 3318
rect 563214 354 563326 480
rect 563072 326 563326 354
rect 563214 -960 563326 326
rect 564410 -960 564522 480
rect 565280 354 565308 3470
rect 566844 480 566872 4762
rect 565606 354 565718 480
rect 565280 326 565718 354
rect 565606 -960 565718 326
rect 566802 -960 566914 480
rect 567580 354 567608 16546
rect 567998 354 568110 480
rect 567580 326 568110 354
rect 568684 354 568712 16546
rect 570326 4856 570382 4865
rect 570326 4791 570382 4800
rect 570340 480 570368 4791
rect 569102 354 569214 480
rect 568684 326 569214 354
rect 567998 -960 568110 326
rect 569102 -960 569214 326
rect 570298 -960 570410 480
rect 571352 354 571380 71023
rect 575478 66872 575534 66881
rect 575478 66807 575534 66816
rect 574100 26920 574152 26926
rect 574100 26862 574152 26868
rect 574112 16574 574140 26862
rect 575492 16574 575520 66807
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 580170 33144 580226 33153
rect 580170 33079 580172 33088
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 576858 25528 576914 25537
rect 576858 25463 576914 25472
rect 576872 16574 576900 25463
rect 580264 22772 580316 22778
rect 580264 22714 580316 22720
rect 579988 20664 580040 20670
rect 579988 20606 580040 20612
rect 580000 19825 580028 20606
rect 579986 19816 580042 19825
rect 579986 19751 580042 19760
rect 574112 16546 575152 16574
rect 575492 16546 575888 16574
rect 576872 16546 576992 16574
rect 572718 6352 572774 6361
rect 572718 6287 572774 6296
rect 572732 480 572760 6287
rect 573914 6216 573970 6225
rect 573914 6151 573970 6160
rect 573928 480 573956 6151
rect 575124 480 575152 16546
rect 571494 354 571606 480
rect 571352 326 571606 354
rect 571494 -960 571606 326
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 575860 354 575888 16546
rect 576278 354 576390 480
rect 575860 326 576390 354
rect 576964 354 576992 16546
rect 580276 6633 580304 22714
rect 580998 17232 581054 17241
rect 580998 17167 581054 17176
rect 581012 16574 581040 17167
rect 581012 16546 581776 16574
rect 581000 7880 581052 7886
rect 581000 7822 581052 7828
rect 580262 6624 580318 6633
rect 580262 6559 580318 6568
rect 578608 6180 578660 6186
rect 578608 6122 578660 6128
rect 578620 480 578648 6122
rect 581012 480 581040 7822
rect 577382 354 577494 480
rect 576964 326 577494 354
rect 576278 -960 576390 326
rect 577382 -960 577494 326
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 581748 354 581776 16546
rect 583392 10464 583444 10470
rect 583392 10406 583444 10412
rect 583404 480 583432 10406
rect 582166 354 582278 480
rect 581748 326 582278 354
rect 582166 -960 582278 326
rect 583362 -960 583474 480
<< via2 >>
rect 2778 684256 2834 684312
rect 3422 671200 3478 671256
rect 3422 658144 3478 658200
rect 2778 632068 2780 632088
rect 2780 632068 2832 632088
rect 2832 632068 2834 632088
rect 2778 632032 2834 632068
rect 3146 579944 3202 580000
rect 3054 566888 3110 566944
rect 3330 553832 3386 553888
rect 2962 527856 3018 527912
rect 3330 475632 3386 475688
rect 2962 423544 3018 423600
rect 3330 410488 3386 410544
rect 3330 371320 3386 371376
rect 3330 358400 3386 358456
rect 3330 345344 3386 345400
rect 2778 319232 2834 319288
rect 2870 306176 2926 306232
rect 3330 293120 3386 293176
rect 3238 267144 3294 267200
rect 2870 254088 2926 254144
rect 3238 241032 3294 241088
rect 3330 214920 3386 214976
rect 3330 201864 3386 201920
rect 3330 162868 3332 162888
rect 3332 162868 3384 162888
rect 3384 162868 3386 162888
rect 3330 162832 3386 162868
rect 3330 149776 3386 149832
rect 2778 136740 2834 136776
rect 2778 136720 2780 136740
rect 2780 136720 2832 136740
rect 2832 136720 2834 136740
rect 3330 110608 3386 110664
rect 3514 619112 3570 619168
rect 3606 606056 3662 606112
rect 3514 501744 3570 501800
rect 3422 79056 3478 79112
rect 3698 514800 3754 514856
rect 3974 462576 4030 462632
rect 3790 449520 3846 449576
rect 3698 97552 3754 97608
rect 3698 84632 3754 84688
rect 3606 79192 3662 79248
rect 3882 397432 3938 397488
rect 4066 188808 4122 188864
rect 6918 79328 6974 79384
rect 6918 75112 6974 75168
rect 3422 71576 3478 71632
rect 3514 58520 3570 58576
rect 3422 45500 3424 45520
rect 3424 45500 3476 45520
rect 3476 45500 3478 45520
rect 3422 45464 3478 45500
rect 3238 19352 3294 19408
rect 3514 32408 3570 32464
rect 3422 6432 3478 6488
rect 9954 8880 10010 8936
rect 8758 4800 8814 4856
rect 13082 77832 13138 77888
rect 11058 76472 11114 76528
rect 117318 137536 117374 137592
rect 117318 136040 117374 136096
rect 117318 134544 117374 134600
rect 117410 133048 117466 133104
rect 117318 131552 117374 131608
rect 117318 130056 117374 130112
rect 117318 128560 117374 128616
rect 117318 127064 117374 127120
rect 117318 125568 117374 125624
rect 117318 124108 117320 124128
rect 117320 124108 117372 124128
rect 117372 124108 117374 124128
rect 117318 124072 117374 124108
rect 117318 122576 117374 122632
rect 117318 121080 117374 121136
rect 117318 119584 117374 119640
rect 117318 118088 117374 118144
rect 117318 116592 117374 116648
rect 117318 115096 117374 115152
rect 118054 113600 118110 113656
rect 118790 112104 118846 112160
rect 118882 110608 118938 110664
rect 119250 109112 119306 109168
rect 119158 107616 119214 107672
rect 119066 106120 119122 106176
rect 118974 104624 119030 104680
rect 118698 101632 118754 101688
rect 118606 95648 118662 95704
rect 118514 94152 118570 94208
rect 118422 92656 118478 92712
rect 118330 91160 118386 91216
rect 118238 89664 118294 89720
rect 118146 88168 118202 88224
rect 118422 86672 118478 86728
rect 118330 82184 118386 82240
rect 26238 73752 26294 73808
rect 25318 9016 25374 9072
rect 27710 7520 27766 7576
rect 60738 75384 60794 75440
rect 44178 75248 44234 75304
rect 48318 73888 48374 73944
rect 45466 9152 45522 9208
rect 63498 22616 63554 22672
rect 80058 76608 80114 76664
rect 60830 9288 60886 9344
rect 63222 6160 63278 6216
rect 78586 9424 78642 9480
rect 95238 21256 95294 21312
rect 115938 76880 115994 76936
rect 97998 76744 98054 76800
rect 118606 85176 118662 85232
rect 118514 83680 118570 83736
rect 118422 81096 118478 81152
rect 119342 78784 119398 78840
rect 120722 103400 120778 103456
rect 120814 100680 120870 100736
rect 120906 98640 120962 98696
rect 120998 97144 121054 97200
rect 179602 80688 179658 80744
rect 119434 78512 119490 78568
rect 101034 4936 101090 4992
rect 114006 10240 114062 10296
rect 119894 7656 119950 7712
rect 118790 3304 118846 3360
rect 129002 77152 129058 77208
rect 129554 77696 129610 77752
rect 130566 78920 130622 78976
rect 131256 79906 131312 79962
rect 131394 79736 131450 79792
rect 131716 79906 131772 79962
rect 131900 79872 131956 79928
rect 131210 77968 131266 78024
rect 131394 79600 131450 79656
rect 131302 77832 131358 77888
rect 132728 79872 132784 79928
rect 131854 79600 131910 79656
rect 132544 79736 132600 79792
rect 133096 79872 133152 79928
rect 133280 79838 133336 79894
rect 133464 79872 133520 79928
rect 132774 79464 132830 79520
rect 132498 78648 132554 78704
rect 133050 78376 133106 78432
rect 133418 79736 133474 79792
rect 134016 79906 134072 79962
rect 134108 79770 134164 79826
rect 134292 79872 134348 79928
rect 133970 78124 134026 78160
rect 133970 78104 133972 78124
rect 133972 78104 134024 78124
rect 134024 78104 134026 78124
rect 134844 79906 134900 79962
rect 134798 79736 134854 79792
rect 134890 79600 134946 79656
rect 134430 77968 134486 78024
rect 134798 79464 134854 79520
rect 134154 77152 134210 77208
rect 135166 79736 135222 79792
rect 135488 79906 135544 79962
rect 135672 79906 135728 79962
rect 136408 79906 136464 79962
rect 135902 79736 135958 79792
rect 136132 79770 136188 79826
rect 135442 79464 135498 79520
rect 135442 77968 135498 78024
rect 135626 77968 135682 78024
rect 135350 75384 135406 75440
rect 136178 79600 136234 79656
rect 136362 79464 136418 79520
rect 136684 79906 136740 79962
rect 137696 79872 137752 79928
rect 136822 78376 136878 78432
rect 136638 76608 136694 76664
rect 137880 79872 137936 79928
rect 138202 79736 138258 79792
rect 137742 79464 137798 79520
rect 137926 78648 137982 78704
rect 138616 79906 138672 79962
rect 138800 79906 138856 79962
rect 139076 79906 139132 79962
rect 138432 79772 138434 79792
rect 138434 79772 138486 79792
rect 138486 79772 138488 79792
rect 138432 79736 138488 79772
rect 138570 79736 138626 79792
rect 138754 79736 138810 79792
rect 139030 79464 139086 79520
rect 139398 79600 139454 79656
rect 139904 79906 139960 79962
rect 140272 79838 140328 79894
rect 139490 76880 139546 76936
rect 140134 79736 140190 79792
rect 140640 79906 140696 79962
rect 139858 79600 139914 79656
rect 139858 75248 139914 75304
rect 140824 79736 140880 79792
rect 140318 79600 140374 79656
rect 141376 79872 141432 79928
rect 141560 79872 141616 79928
rect 141744 79906 141800 79962
rect 141928 79838 141984 79894
rect 141698 79736 141754 79792
rect 140594 79600 140650 79656
rect 140870 79600 140926 79656
rect 140962 74976 141018 75032
rect 141330 79600 141386 79656
rect 141514 79464 141570 79520
rect 141790 79600 141846 79656
rect 141790 78920 141846 78976
rect 142296 79872 142352 79928
rect 142158 75248 142214 75304
rect 143032 79872 143088 79928
rect 142894 79736 142950 79792
rect 143308 79872 143364 79928
rect 143492 79906 143548 79962
rect 143170 76744 143226 76800
rect 142986 76472 143042 76528
rect 143446 76608 143502 76664
rect 143768 79872 143824 79928
rect 143814 79736 143870 79792
rect 143630 79600 143686 79656
rect 143630 79464 143686 79520
rect 142802 44240 142858 44296
rect 144044 79736 144100 79792
rect 144412 79906 144468 79962
rect 143906 78104 143962 78160
rect 144596 79736 144652 79792
rect 144458 79600 144514 79656
rect 144182 66136 144238 66192
rect 145148 79736 145204 79792
rect 145608 79838 145664 79894
rect 144918 79600 144974 79656
rect 145010 79464 145066 79520
rect 144826 78104 144882 78160
rect 144734 76608 144790 76664
rect 144642 75520 144698 75576
rect 145286 79464 145342 79520
rect 145746 79736 145802 79792
rect 146344 79838 146400 79894
rect 145562 79464 145618 79520
rect 145470 77288 145526 77344
rect 146114 79600 146170 79656
rect 146206 77424 146262 77480
rect 146942 77968 146998 78024
rect 147264 79872 147320 79928
rect 147310 77424 147366 77480
rect 147494 79600 147550 79656
rect 148000 79872 148056 79928
rect 148184 79906 148240 79962
rect 148644 79872 148700 79928
rect 147402 77288 147458 77344
rect 147586 76336 147642 76392
rect 148874 79736 148930 79792
rect 149288 79872 149344 79928
rect 149656 79872 149712 79928
rect 148322 78376 148378 78432
rect 148414 76608 148470 76664
rect 148322 75384 148378 75440
rect 148690 77152 148746 77208
rect 149058 79464 149114 79520
rect 148966 76608 149022 76664
rect 148874 75112 148930 75168
rect 150024 79906 150080 79962
rect 150208 79906 150264 79962
rect 150162 79736 150218 79792
rect 149702 79600 149758 79656
rect 149610 79464 149666 79520
rect 149610 78920 149666 78976
rect 150070 79600 150126 79656
rect 150576 79906 150632 79962
rect 150760 79906 150816 79962
rect 150944 79872 151000 79928
rect 151128 79906 151184 79962
rect 150806 79736 150862 79792
rect 150254 79464 150310 79520
rect 150162 78648 150218 78704
rect 150346 77016 150402 77072
rect 150806 79600 150862 79656
rect 151404 79906 151460 79962
rect 150622 76608 150678 76664
rect 151680 79906 151736 79962
rect 151818 79736 151874 79792
rect 151634 79600 151690 79656
rect 151818 79600 151874 79656
rect 151726 76608 151782 76664
rect 152508 79872 152564 79928
rect 153060 79872 153116 79928
rect 153014 77288 153070 77344
rect 153336 79906 153392 79962
rect 153520 79872 153576 79928
rect 153704 79906 153760 79962
rect 154164 79906 154220 79962
rect 153382 79736 153438 79792
rect 153290 77424 153346 77480
rect 153474 77288 153530 77344
rect 153106 76880 153162 76936
rect 153290 76608 153346 76664
rect 153842 79600 153898 79656
rect 154624 79872 154680 79928
rect 154532 79736 154588 79792
rect 154302 77288 154358 77344
rect 154210 76744 154266 76800
rect 154486 77424 154542 77480
rect 155084 79872 155140 79928
rect 154854 79464 154910 79520
rect 154854 78104 154910 78160
rect 155360 79736 155416 79792
rect 155038 79600 155094 79656
rect 155130 79464 155186 79520
rect 155820 79906 155876 79962
rect 155406 79464 155462 79520
rect 155222 77288 155278 77344
rect 155774 79464 155830 79520
rect 155774 78376 155830 78432
rect 156142 79736 156198 79792
rect 156556 79872 156612 79928
rect 155866 76608 155922 76664
rect 156234 79600 156290 79656
rect 156878 79736 156934 79792
rect 157108 79906 157164 79962
rect 156510 79600 156566 79656
rect 156326 77288 156382 77344
rect 156694 79500 156696 79520
rect 156696 79500 156748 79520
rect 156748 79500 156750 79520
rect 156694 79464 156750 79500
rect 157338 79464 157394 79520
rect 157246 77560 157302 77616
rect 157154 77424 157210 77480
rect 157844 79872 157900 79928
rect 158304 79906 158360 79962
rect 158580 79872 158636 79928
rect 158258 78920 158314 78976
rect 158350 78648 158406 78704
rect 158626 77288 158682 77344
rect 159316 79872 159372 79928
rect 159960 79838 160016 79894
rect 160236 79872 160292 79928
rect 159914 79464 159970 79520
rect 160006 77288 160062 77344
rect 159362 65456 159418 65512
rect 161156 79872 161212 79928
rect 161524 79872 161580 79928
rect 161202 79736 161258 79792
rect 161294 79464 161350 79520
rect 160834 76472 160890 76528
rect 161386 76472 161442 76528
rect 162168 79872 162224 79928
rect 162720 79906 162776 79962
rect 161846 79600 161902 79656
rect 161570 77832 161626 77888
rect 162030 78240 162086 78296
rect 162674 76200 162730 76256
rect 162490 76064 162546 76120
rect 163226 78376 163282 78432
rect 164192 79838 164248 79894
rect 163732 79736 163788 79792
rect 164054 78920 164110 78976
rect 163962 78648 164018 78704
rect 164330 79500 164332 79520
rect 164332 79500 164384 79520
rect 164384 79500 164386 79520
rect 164330 79464 164386 79500
rect 165020 79872 165076 79928
rect 165572 79872 165628 79928
rect 165940 79906 165996 79962
rect 164698 76200 164754 76256
rect 165526 79736 165582 79792
rect 165250 77968 165306 78024
rect 165434 78104 165490 78160
rect 165618 78920 165674 78976
rect 165526 77968 165582 78024
rect 165618 77560 165674 77616
rect 166676 79872 166732 79928
rect 166584 79736 166640 79792
rect 166354 79600 166410 79656
rect 166538 79600 166594 79656
rect 166446 77968 166502 78024
rect 167320 79872 167376 79928
rect 166722 77424 166778 77480
rect 166630 77288 166686 77344
rect 166998 77560 167054 77616
rect 168056 79872 168112 79928
rect 168240 79872 168296 79928
rect 168792 79872 168848 79928
rect 168976 79906 169032 79962
rect 169528 79838 169584 79894
rect 168838 79736 168894 79792
rect 168010 77832 168066 77888
rect 168102 77288 168158 77344
rect 168654 79600 168710 79656
rect 168286 79464 168342 79520
rect 168194 75248 168250 75304
rect 168838 79464 168894 79520
rect 168562 78648 168618 78704
rect 170264 79906 170320 79962
rect 169390 79500 169392 79520
rect 169392 79500 169444 79520
rect 169444 79500 169446 79520
rect 169390 79464 169446 79500
rect 169574 79600 169630 79656
rect 169666 79464 169722 79520
rect 169942 77696 169998 77752
rect 170540 79906 170596 79962
rect 170724 79872 170780 79928
rect 170908 79906 170964 79962
rect 171092 79872 171148 79928
rect 170494 79600 170550 79656
rect 170678 78648 170734 78704
rect 170862 79600 170918 79656
rect 171046 79464 171102 79520
rect 171322 79600 171378 79656
rect 171736 79872 171792 79928
rect 171644 79736 171700 79792
rect 170954 78240 171010 78296
rect 170954 77832 171010 77888
rect 170770 77560 170826 77616
rect 170402 63552 170458 63608
rect 162490 4936 162546 4992
rect 161294 3440 161350 3496
rect 166078 4800 166134 4856
rect 163686 3304 163742 3360
rect 171690 79600 171746 79656
rect 171598 78240 171654 78296
rect 172472 79872 172528 79928
rect 172656 79872 172712 79928
rect 172380 79736 172436 79792
rect 172932 79872 172988 79928
rect 172058 78648 172114 78704
rect 172058 78240 172114 78296
rect 172242 78104 172298 78160
rect 172150 77424 172206 77480
rect 172610 79464 172666 79520
rect 172702 78648 172758 78704
rect 172978 79736 173034 79792
rect 172978 79600 173034 79656
rect 173576 79906 173632 79962
rect 173530 79736 173586 79792
rect 173162 79636 173164 79656
rect 173164 79636 173216 79656
rect 173216 79636 173218 79656
rect 173162 79600 173218 79636
rect 173070 78104 173126 78160
rect 173254 78956 173256 78976
rect 173256 78956 173308 78976
rect 173308 78956 173310 78976
rect 173254 78920 173310 78956
rect 174036 79906 174092 79962
rect 173530 79600 173586 79656
rect 173714 79464 173770 79520
rect 173622 78920 173678 78976
rect 173806 78648 173862 78704
rect 174956 79736 175012 79792
rect 175232 79872 175288 79928
rect 175508 79872 175564 79928
rect 175186 79620 175242 79656
rect 175186 79600 175188 79620
rect 175188 79600 175240 79620
rect 175240 79600 175242 79620
rect 175278 79192 175334 79248
rect 175094 78920 175150 78976
rect 175002 78648 175058 78704
rect 175278 77832 175334 77888
rect 175784 79736 175840 79792
rect 176520 79906 176576 79962
rect 176796 79872 176852 79928
rect 176750 79772 176752 79792
rect 176752 79772 176804 79792
rect 176804 79772 176806 79792
rect 176750 79736 176806 79772
rect 177348 79872 177404 79928
rect 175646 79056 175702 79112
rect 175554 78920 175610 78976
rect 175462 78648 175518 78704
rect 175830 78104 175886 78160
rect 176474 79600 176530 79656
rect 176290 79348 176346 79384
rect 176290 79328 176292 79348
rect 176292 79328 176344 79348
rect 176344 79328 176346 79348
rect 176658 79328 176714 79384
rect 176106 75656 176162 75712
rect 177808 79872 177864 79928
rect 177210 78784 177266 78840
rect 176934 78376 176990 78432
rect 176934 78104 176990 78160
rect 177762 79736 177818 79792
rect 178360 79872 178416 79928
rect 177762 79636 177764 79656
rect 177764 79636 177816 79656
rect 177816 79636 177818 79656
rect 177578 79328 177634 79384
rect 177762 79600 177818 79636
rect 177670 78920 177726 78976
rect 177486 78784 177542 78840
rect 177578 78376 177634 78432
rect 176566 74432 176622 74488
rect 175738 3440 175794 3496
rect 178038 79192 178094 79248
rect 178222 79192 178278 79248
rect 179142 79056 179198 79112
rect 179878 80416 179934 80472
rect 180062 80280 180118 80336
rect 179786 79464 179842 79520
rect 180706 80144 180762 80200
rect 180246 80008 180302 80064
rect 180246 78648 180302 78704
rect 189538 136992 189594 137048
rect 189446 126112 189502 126168
rect 189446 118496 189502 118552
rect 189446 117136 189502 117192
rect 189446 114144 189502 114200
rect 179694 78240 179750 78296
rect 180062 76336 180118 76392
rect 180246 78104 180302 78160
rect 180798 75520 180854 75576
rect 182178 69536 182234 69592
rect 183558 25608 183614 25664
rect 189722 133592 189778 133648
rect 189630 123936 189686 123992
rect 190642 134544 190698 134600
rect 190550 127064 190606 127120
rect 190458 119584 190514 119640
rect 190734 131552 190790 131608
rect 191010 136040 191066 136096
rect 190918 122576 190974 122632
rect 190826 115096 190882 115152
rect 192022 130056 192078 130112
rect 191930 128560 191986 128616
rect 191838 121080 191894 121136
rect 192206 101632 192262 101688
rect 192206 100136 192262 100192
rect 192206 98640 192262 98696
rect 192666 95648 192722 95704
rect 192666 83680 192722 83736
rect 193126 112104 193182 112160
rect 193126 110608 193182 110664
rect 193034 109112 193090 109168
rect 193034 107616 193090 107672
rect 193126 106156 193128 106176
rect 193128 106156 193180 106176
rect 193180 106156 193182 106176
rect 193126 106120 193182 106156
rect 193126 104660 193128 104680
rect 193128 104660 193180 104680
rect 193180 104660 193182 104680
rect 193126 104624 193182 104660
rect 193126 103164 193128 103184
rect 193128 103164 193180 103184
rect 193180 103164 193182 103184
rect 193126 103128 193182 103164
rect 193126 97144 193182 97200
rect 193126 94152 193182 94208
rect 192850 82184 192906 82240
rect 193126 92656 193182 92712
rect 193126 91160 193182 91216
rect 193126 89684 193182 89720
rect 193126 89664 193128 89684
rect 193128 89664 193180 89684
rect 193180 89664 193182 89684
rect 193126 88168 193182 88224
rect 193126 86672 193182 86728
rect 193126 85176 193182 85232
rect 196898 80960 196954 81016
rect 196714 80552 196770 80608
rect 266358 79600 266414 79656
rect 260102 77968 260158 78024
rect 233238 77152 233294 77208
rect 200118 62736 200174 62792
rect 201590 24384 201646 24440
rect 215298 28192 215354 28248
rect 214470 3712 214526 3768
rect 216678 18672 216734 18728
rect 218058 3576 218114 3632
rect 235998 29552 236054 29608
rect 232226 6024 232282 6080
rect 235814 6840 235870 6896
rect 234618 5208 234674 5264
rect 253938 77016 253994 77072
rect 251178 73888 251234 73944
rect 251270 7520 251326 7576
rect 253478 6704 253534 6760
rect 271878 30912 271934 30968
rect 269118 20168 269174 20224
rect 271234 9152 271290 9208
rect 289818 76880 289874 76936
rect 287058 73752 287114 73808
rect 285678 26832 285734 26888
rect 288990 10376 289046 10432
rect 303618 76744 303674 76800
rect 306378 55800 306434 55856
rect 305550 16088 305606 16144
rect 307942 6568 307998 6624
rect 331218 79464 331274 79520
rect 324318 76608 324374 76664
rect 324410 12280 324466 12336
rect 338670 5072 338726 5128
rect 340878 13096 340934 13152
rect 340970 12144 341026 12200
rect 343362 9016 343418 9072
rect 357438 20032 357494 20088
rect 356334 14864 356390 14920
rect 359462 14728 359518 14784
rect 357530 12008 357586 12064
rect 397458 78920 397514 78976
rect 462318 78784 462374 78840
rect 396078 76472 396134 76528
rect 376758 68176 376814 68232
rect 378138 23024 378194 23080
rect 395342 15952 395398 16008
rect 394238 14592 394294 14648
rect 392582 11872 392638 11928
rect 408498 17720 408554 17776
rect 414018 22888 414074 22944
rect 412638 17584 412694 17640
rect 410798 15816 410854 15872
rect 429198 36488 429254 36544
rect 430578 18536 430634 18592
rect 480258 77832 480314 77888
rect 431958 75384 432014 75440
rect 444378 19896 444434 19952
rect 446218 4936 446274 4992
rect 448518 11736 448574 11792
rect 448610 6432 448666 6488
rect 466458 17448 466514 17504
rect 463974 14456 464030 14512
rect 466274 8880 466330 8936
rect 481638 75248 481694 75304
rect 483018 64232 483074 64288
rect 481730 10240 481786 10296
rect 484766 12960 484822 13016
rect 502338 22752 502394 22808
rect 518898 61376 518954 61432
rect 517518 17312 517574 17368
rect 520278 22616 520334 22672
rect 517150 11600 517206 11656
rect 580262 697176 580318 697232
rect 579618 683848 579674 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580170 644000 580226 644056
rect 579986 630808 580042 630864
rect 580170 617480 580226 617536
rect 580170 590960 580226 591016
rect 580170 577632 580226 577688
rect 580170 564304 580226 564360
rect 579894 537784 579950 537840
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 511264 580226 511320
rect 579618 458088 579674 458144
rect 579710 418240 579766 418296
rect 580170 404912 580226 404968
rect 580170 378392 580226 378448
rect 580170 365064 580226 365120
rect 580170 351908 580172 351928
rect 580172 351908 580224 351928
rect 580224 351908 580226 351928
rect 580170 351872 580226 351908
rect 580170 312024 580226 312080
rect 580170 298696 580226 298752
rect 580170 272176 580226 272232
rect 579618 258848 579674 258904
rect 580170 245520 580226 245576
rect 580170 219000 580226 219056
rect 580170 205692 580226 205728
rect 580170 205672 580172 205692
rect 580172 205672 580224 205692
rect 580224 205672 580226 205692
rect 580170 192480 580226 192536
rect 580170 179152 580226 179208
rect 579618 165824 579674 165880
rect 579986 152632 580042 152688
rect 580170 125976 580226 126032
rect 580078 112784 580134 112840
rect 579986 86128 580042 86184
rect 580170 81096 580226 81152
rect 535458 75112 535514 75168
rect 534078 24248 534134 24304
rect 536838 65456 536894 65512
rect 538218 24112 538274 24168
rect 544382 3440 544438 3496
rect 580354 484608 580410 484664
rect 580262 79328 580318 79384
rect 580446 471416 580502 471472
rect 580538 431568 580594 431624
rect 580630 325216 580686 325272
rect 580814 232328 580870 232384
rect 580722 139304 580778 139360
rect 580906 99456 580962 99512
rect 580814 80824 580870 80880
rect 580630 80688 580686 80744
rect 580538 78648 580594 78704
rect 580170 72936 580226 72992
rect 571338 71032 571394 71088
rect 554778 64096 554834 64152
rect 556158 46144 556214 46200
rect 558550 3304 558606 3360
rect 570326 4800 570382 4856
rect 575478 66816 575534 66872
rect 580170 59608 580226 59664
rect 580170 46280 580226 46336
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 576858 25472 576914 25528
rect 579986 19760 580042 19816
rect 572718 6296 572774 6352
rect 573914 6160 573970 6216
rect 580998 17176 581054 17232
rect 580262 6568 580318 6624
<< metal3 >>
rect -960 697220 480 697460
rect 580257 697234 580323 697237
rect 583520 697234 584960 697324
rect 580257 697232 584960 697234
rect 580257 697176 580262 697232
rect 580318 697176 584960 697232
rect 580257 697174 584960 697176
rect 580257 697171 580323 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 2773 684314 2839 684317
rect -960 684312 2839 684314
rect -960 684256 2778 684312
rect 2834 684256 2839 684312
rect -960 684254 2839 684256
rect -960 684164 480 684254
rect 2773 684251 2839 684254
rect 579613 683906 579679 683909
rect 583520 683906 584960 683996
rect 579613 683904 584960 683906
rect 579613 683848 579618 683904
rect 579674 683848 584960 683904
rect 579613 683846 584960 683848
rect 579613 683843 579679 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3417 671258 3483 671261
rect -960 671256 3483 671258
rect -960 671200 3422 671256
rect 3478 671200 3483 671256
rect -960 671198 3483 671200
rect -960 671108 480 671198
rect 3417 671195 3483 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 2773 632090 2839 632093
rect -960 632088 2839 632090
rect -960 632032 2778 632088
rect 2834 632032 2839 632088
rect -960 632030 2839 632032
rect -960 631940 480 632030
rect 2773 632027 2839 632030
rect 579981 630866 580047 630869
rect 583520 630866 584960 630956
rect 579981 630864 584960 630866
rect 579981 630808 579986 630864
rect 580042 630808 584960 630864
rect 579981 630806 584960 630808
rect 579981 630803 580047 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3509 619170 3575 619173
rect -960 619168 3575 619170
rect -960 619112 3514 619168
rect 3570 619112 3575 619168
rect -960 619110 3575 619112
rect -960 619020 480 619110
rect 3509 619107 3575 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3601 606114 3667 606117
rect -960 606112 3667 606114
rect -960 606056 3606 606112
rect 3662 606056 3667 606112
rect -960 606054 3667 606056
rect -960 605964 480 606054
rect 3601 606051 3667 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 580165 591018 580231 591021
rect 583520 591018 584960 591108
rect 580165 591016 584960 591018
rect 580165 590960 580170 591016
rect 580226 590960 584960 591016
rect 580165 590958 584960 590960
rect 580165 590955 580231 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3141 580002 3207 580005
rect -960 580000 3207 580002
rect -960 579944 3146 580000
rect 3202 579944 3207 580000
rect -960 579942 3207 579944
rect -960 579852 480 579942
rect 3141 579939 3207 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3049 566946 3115 566949
rect -960 566944 3115 566946
rect -960 566888 3054 566944
rect 3110 566888 3115 566944
rect -960 566886 3115 566888
rect -960 566796 480 566886
rect 3049 566883 3115 566886
rect 580165 564362 580231 564365
rect 583520 564362 584960 564452
rect 580165 564360 584960 564362
rect 580165 564304 580170 564360
rect 580226 564304 584960 564360
rect 580165 564302 584960 564304
rect 580165 564299 580231 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3325 553890 3391 553893
rect -960 553888 3391 553890
rect -960 553832 3330 553888
rect 3386 553832 3391 553888
rect -960 553830 3391 553832
rect -960 553740 480 553830
rect 3325 553827 3391 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 579889 537842 579955 537845
rect 583520 537842 584960 537932
rect 579889 537840 584960 537842
rect 579889 537784 579894 537840
rect 579950 537784 584960 537840
rect 579889 537782 584960 537784
rect 579889 537779 579955 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 2957 527914 3023 527917
rect -960 527912 3023 527914
rect -960 527856 2962 527912
rect 3018 527856 3023 527912
rect -960 527854 3023 527856
rect -960 527764 480 527854
rect 2957 527851 3023 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3693 514858 3759 514861
rect -960 514856 3759 514858
rect -960 514800 3698 514856
rect 3754 514800 3759 514856
rect -960 514798 3759 514800
rect -960 514708 480 514798
rect 3693 514795 3759 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3509 501802 3575 501805
rect -960 501800 3575 501802
rect -960 501744 3514 501800
rect 3570 501744 3575 501800
rect -960 501742 3575 501744
rect -960 501652 480 501742
rect 3509 501739 3575 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580349 484666 580415 484669
rect 583520 484666 584960 484756
rect 580349 484664 584960 484666
rect 580349 484608 580354 484664
rect 580410 484608 584960 484664
rect 580349 484606 584960 484608
rect 580349 484603 580415 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3325 475690 3391 475693
rect -960 475688 3391 475690
rect -960 475632 3330 475688
rect 3386 475632 3391 475688
rect -960 475630 3391 475632
rect -960 475540 480 475630
rect 3325 475627 3391 475630
rect 580441 471474 580507 471477
rect 583520 471474 584960 471564
rect 580441 471472 584960 471474
rect 580441 471416 580446 471472
rect 580502 471416 584960 471472
rect 580441 471414 584960 471416
rect 580441 471411 580507 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3969 462634 4035 462637
rect -960 462632 4035 462634
rect -960 462576 3974 462632
rect 4030 462576 4035 462632
rect -960 462574 4035 462576
rect -960 462484 480 462574
rect 3969 462571 4035 462574
rect 579613 458146 579679 458149
rect 583520 458146 584960 458236
rect 579613 458144 584960 458146
rect 579613 458088 579618 458144
rect 579674 458088 584960 458144
rect 579613 458086 584960 458088
rect 579613 458083 579679 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3785 449578 3851 449581
rect -960 449576 3851 449578
rect -960 449520 3790 449576
rect 3846 449520 3851 449576
rect -960 449518 3851 449520
rect -960 449428 480 449518
rect 3785 449515 3851 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 580533 431626 580599 431629
rect 583520 431626 584960 431716
rect 580533 431624 584960 431626
rect 580533 431568 580538 431624
rect 580594 431568 584960 431624
rect 580533 431566 584960 431568
rect 580533 431563 580599 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 2957 423602 3023 423605
rect -960 423600 3023 423602
rect -960 423544 2962 423600
rect 3018 423544 3023 423600
rect -960 423542 3023 423544
rect -960 423452 480 423542
rect 2957 423539 3023 423542
rect 579705 418298 579771 418301
rect 583520 418298 584960 418388
rect 579705 418296 584960 418298
rect 579705 418240 579710 418296
rect 579766 418240 584960 418296
rect 579705 418238 584960 418240
rect 579705 418235 579771 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3325 410546 3391 410549
rect -960 410544 3391 410546
rect -960 410488 3330 410544
rect 3386 410488 3391 410544
rect -960 410486 3391 410488
rect -960 410396 480 410486
rect 3325 410483 3391 410486
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3877 397490 3943 397493
rect -960 397488 3943 397490
rect -960 397432 3882 397488
rect 3938 397432 3943 397488
rect -960 397430 3943 397432
rect -960 397340 480 397430
rect 3877 397427 3943 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 3325 371378 3391 371381
rect -960 371376 3391 371378
rect -960 371320 3330 371376
rect 3386 371320 3391 371376
rect -960 371318 3391 371320
rect -960 371228 480 371318
rect 3325 371315 3391 371318
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 3325 358458 3391 358461
rect -960 358456 3391 358458
rect -960 358400 3330 358456
rect 3386 358400 3391 358456
rect -960 358398 3391 358400
rect -960 358308 480 358398
rect 3325 358395 3391 358398
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 3325 345402 3391 345405
rect -960 345400 3391 345402
rect -960 345344 3330 345400
rect 3386 345344 3391 345400
rect -960 345342 3391 345344
rect -960 345252 480 345342
rect 3325 345339 3391 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 580625 325274 580691 325277
rect 583520 325274 584960 325364
rect 580625 325272 584960 325274
rect 580625 325216 580630 325272
rect 580686 325216 584960 325272
rect 580625 325214 584960 325216
rect 580625 325211 580691 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 2773 319290 2839 319293
rect -960 319288 2839 319290
rect -960 319232 2778 319288
rect 2834 319232 2839 319288
rect -960 319230 2839 319232
rect -960 319140 480 319230
rect 2773 319227 2839 319230
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 2865 306234 2931 306237
rect -960 306232 2931 306234
rect -960 306176 2870 306232
rect 2926 306176 2931 306232
rect -960 306174 2931 306176
rect -960 306084 480 306174
rect 2865 306171 2931 306174
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 3325 293178 3391 293181
rect -960 293176 3391 293178
rect -960 293120 3330 293176
rect 3386 293120 3391 293176
rect -960 293118 3391 293120
rect -960 293028 480 293118
rect 3325 293115 3391 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 3233 267202 3299 267205
rect -960 267200 3299 267202
rect -960 267144 3238 267200
rect 3294 267144 3299 267200
rect -960 267142 3299 267144
rect -960 267052 480 267142
rect 3233 267139 3299 267142
rect 579613 258906 579679 258909
rect 583520 258906 584960 258996
rect 579613 258904 584960 258906
rect 579613 258848 579618 258904
rect 579674 258848 584960 258904
rect 579613 258846 584960 258848
rect 579613 258843 579679 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 2865 254146 2931 254149
rect -960 254144 2931 254146
rect -960 254088 2870 254144
rect 2926 254088 2931 254144
rect -960 254086 2931 254088
rect -960 253996 480 254086
rect 2865 254083 2931 254086
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 3233 241090 3299 241093
rect -960 241088 3299 241090
rect -960 241032 3238 241088
rect 3294 241032 3299 241088
rect -960 241030 3299 241032
rect -960 240940 480 241030
rect 3233 241027 3299 241030
rect 580809 232386 580875 232389
rect 583520 232386 584960 232476
rect 580809 232384 584960 232386
rect 580809 232328 580814 232384
rect 580870 232328 584960 232384
rect 580809 232326 584960 232328
rect 580809 232323 580875 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 580165 219058 580231 219061
rect 583520 219058 584960 219148
rect 580165 219056 584960 219058
rect 580165 219000 580170 219056
rect 580226 219000 584960 219056
rect 580165 218998 584960 219000
rect 580165 218995 580231 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 3325 214978 3391 214981
rect -960 214976 3391 214978
rect -960 214920 3330 214976
rect 3386 214920 3391 214976
rect -960 214918 3391 214920
rect -960 214828 480 214918
rect 3325 214915 3391 214918
rect 580165 205730 580231 205733
rect 583520 205730 584960 205820
rect 580165 205728 584960 205730
rect 580165 205672 580170 205728
rect 580226 205672 584960 205728
rect 580165 205670 584960 205672
rect 580165 205667 580231 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3325 201922 3391 201925
rect -960 201920 3391 201922
rect -960 201864 3330 201920
rect 3386 201864 3391 201920
rect -960 201862 3391 201864
rect -960 201772 480 201862
rect 3325 201859 3391 201862
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 4061 188866 4127 188869
rect -960 188864 4127 188866
rect -960 188808 4066 188864
rect 4122 188808 4127 188864
rect -960 188806 4127 188808
rect -960 188716 480 188806
rect 4061 188803 4127 188806
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 579613 165882 579679 165885
rect 583520 165882 584960 165972
rect 579613 165880 584960 165882
rect 579613 165824 579618 165880
rect 579674 165824 584960 165880
rect 579613 165822 584960 165824
rect 579613 165819 579679 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3325 162890 3391 162893
rect -960 162888 3391 162890
rect -960 162832 3330 162888
rect 3386 162832 3391 162888
rect -960 162830 3391 162832
rect -960 162740 480 162830
rect 3325 162827 3391 162830
rect 579981 152690 580047 152693
rect 583520 152690 584960 152780
rect 579981 152688 584960 152690
rect 579981 152632 579986 152688
rect 580042 152632 584960 152688
rect 579981 152630 584960 152632
rect 579981 152627 580047 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3325 149834 3391 149837
rect -960 149832 3391 149834
rect -960 149776 3330 149832
rect 3386 149776 3391 149832
rect -960 149774 3391 149776
rect -960 149684 480 149774
rect 3325 149771 3391 149774
rect 580717 139362 580783 139365
rect 583520 139362 584960 139452
rect 580717 139360 584960 139362
rect 580717 139304 580722 139360
rect 580778 139304 584960 139360
rect 580717 139302 584960 139304
rect 580717 139299 580783 139302
rect 583520 139212 584960 139302
rect 117313 137594 117379 137597
rect 117313 137592 120060 137594
rect 117313 137536 117318 137592
rect 117374 137536 120060 137592
rect 117313 137534 120060 137536
rect 117313 137531 117379 137534
rect 189582 137053 189642 137564
rect 189533 137048 189642 137053
rect 189533 136992 189538 137048
rect 189594 136992 189642 137048
rect 189533 136990 189642 136992
rect 189533 136987 189599 136990
rect -960 136778 480 136868
rect 2773 136778 2839 136781
rect -960 136776 2839 136778
rect -960 136720 2778 136776
rect 2834 136720 2839 136776
rect -960 136718 2839 136720
rect -960 136628 480 136718
rect 2773 136715 2839 136718
rect 117313 136098 117379 136101
rect 191005 136098 191071 136101
rect 117313 136096 120060 136098
rect 117313 136040 117318 136096
rect 117374 136040 120060 136096
rect 117313 136038 120060 136040
rect 189796 136096 191071 136098
rect 189796 136040 191010 136096
rect 191066 136040 191071 136096
rect 189796 136038 191071 136040
rect 117313 136035 117379 136038
rect 191005 136035 191071 136038
rect 117313 134602 117379 134605
rect 190637 134602 190703 134605
rect 117313 134600 120060 134602
rect 117313 134544 117318 134600
rect 117374 134544 120060 134600
rect 117313 134542 120060 134544
rect 189796 134600 190703 134602
rect 189796 134544 190642 134600
rect 190698 134544 190703 134600
rect 189796 134542 190703 134544
rect 117313 134539 117379 134542
rect 190637 134539 190703 134542
rect 189717 133650 189783 133653
rect 189717 133648 189826 133650
rect 189717 133592 189722 133648
rect 189778 133592 189826 133648
rect 189717 133587 189826 133592
rect 117405 133106 117471 133109
rect 117405 133104 120060 133106
rect 117405 133048 117410 133104
rect 117466 133048 120060 133104
rect 189766 133076 189826 133587
rect 117405 133046 120060 133048
rect 117405 133043 117471 133046
rect 117313 131610 117379 131613
rect 190729 131610 190795 131613
rect 117313 131608 120060 131610
rect 117313 131552 117318 131608
rect 117374 131552 120060 131608
rect 117313 131550 120060 131552
rect 189796 131608 190795 131610
rect 189796 131552 190734 131608
rect 190790 131552 190795 131608
rect 189796 131550 190795 131552
rect 117313 131547 117379 131550
rect 190729 131547 190795 131550
rect 117313 130114 117379 130117
rect 192017 130114 192083 130117
rect 117313 130112 120060 130114
rect 117313 130056 117318 130112
rect 117374 130056 120060 130112
rect 117313 130054 120060 130056
rect 189796 130112 192083 130114
rect 189796 130056 192022 130112
rect 192078 130056 192083 130112
rect 189796 130054 192083 130056
rect 117313 130051 117379 130054
rect 192017 130051 192083 130054
rect 117313 128618 117379 128621
rect 191925 128618 191991 128621
rect 117313 128616 120060 128618
rect 117313 128560 117318 128616
rect 117374 128560 120060 128616
rect 117313 128558 120060 128560
rect 189796 128616 191991 128618
rect 189796 128560 191930 128616
rect 191986 128560 191991 128616
rect 189796 128558 191991 128560
rect 117313 128555 117379 128558
rect 191925 128555 191991 128558
rect 117313 127122 117379 127125
rect 190545 127122 190611 127125
rect 117313 127120 120060 127122
rect 117313 127064 117318 127120
rect 117374 127064 120060 127120
rect 117313 127062 120060 127064
rect 189796 127120 190611 127122
rect 189796 127064 190550 127120
rect 190606 127064 190611 127120
rect 189796 127062 190611 127064
rect 117313 127059 117379 127062
rect 190545 127059 190611 127062
rect 189441 126170 189507 126173
rect 189398 126168 189507 126170
rect 189398 126112 189446 126168
rect 189502 126112 189507 126168
rect 189398 126107 189507 126112
rect 117313 125626 117379 125629
rect 117313 125624 120060 125626
rect 117313 125568 117318 125624
rect 117374 125568 120060 125624
rect 189398 125596 189458 126107
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect 117313 125566 120060 125568
rect 117313 125563 117379 125566
rect 117313 124130 117379 124133
rect 117313 124128 120060 124130
rect 117313 124072 117318 124128
rect 117374 124072 120060 124128
rect 117313 124070 120060 124072
rect 117313 124067 117379 124070
rect 189582 123997 189642 124100
rect 189582 123992 189691 123997
rect 189582 123936 189630 123992
rect 189686 123936 189691 123992
rect 189582 123934 189691 123936
rect 189625 123931 189691 123934
rect -960 123572 480 123812
rect 117313 122634 117379 122637
rect 190913 122634 190979 122637
rect 117313 122632 120060 122634
rect 117313 122576 117318 122632
rect 117374 122576 120060 122632
rect 117313 122574 120060 122576
rect 189796 122632 190979 122634
rect 189796 122576 190918 122632
rect 190974 122576 190979 122632
rect 189796 122574 190979 122576
rect 117313 122571 117379 122574
rect 190913 122571 190979 122574
rect 117313 121138 117379 121141
rect 191833 121138 191899 121141
rect 117313 121136 120060 121138
rect 117313 121080 117318 121136
rect 117374 121080 120060 121136
rect 117313 121078 120060 121080
rect 189796 121136 191899 121138
rect 189796 121080 191838 121136
rect 191894 121080 191899 121136
rect 189796 121078 191899 121080
rect 117313 121075 117379 121078
rect 191833 121075 191899 121078
rect 117313 119642 117379 119645
rect 190453 119642 190519 119645
rect 117313 119640 120060 119642
rect 117313 119584 117318 119640
rect 117374 119584 120060 119640
rect 117313 119582 120060 119584
rect 189796 119640 190519 119642
rect 189796 119584 190458 119640
rect 190514 119584 190519 119640
rect 189796 119582 190519 119584
rect 117313 119579 117379 119582
rect 190453 119579 190519 119582
rect 189441 118554 189507 118557
rect 189398 118552 189507 118554
rect 189398 118496 189446 118552
rect 189502 118496 189507 118552
rect 189398 118491 189507 118496
rect 117313 118146 117379 118149
rect 117313 118144 120060 118146
rect 117313 118088 117318 118144
rect 117374 118088 120060 118144
rect 189398 118116 189458 118491
rect 117313 118086 120060 118088
rect 117313 118083 117379 118086
rect 189441 117194 189507 117197
rect 189398 117192 189507 117194
rect 189398 117136 189446 117192
rect 189502 117136 189507 117192
rect 189398 117131 189507 117136
rect 117313 116650 117379 116653
rect 117313 116648 120060 116650
rect 117313 116592 117318 116648
rect 117374 116592 120060 116648
rect 189398 116620 189458 117131
rect 117313 116590 120060 116592
rect 117313 116587 117379 116590
rect 117313 115154 117379 115157
rect 190821 115154 190887 115157
rect 117313 115152 120060 115154
rect 117313 115096 117318 115152
rect 117374 115096 120060 115152
rect 117313 115094 120060 115096
rect 189796 115152 190887 115154
rect 189796 115096 190826 115152
rect 190882 115096 190887 115152
rect 189796 115094 190887 115096
rect 117313 115091 117379 115094
rect 190821 115091 190887 115094
rect 189441 114202 189507 114205
rect 189398 114200 189507 114202
rect 189398 114144 189446 114200
rect 189502 114144 189507 114200
rect 189398 114139 189507 114144
rect 118049 113658 118115 113661
rect 118049 113656 120060 113658
rect 118049 113600 118054 113656
rect 118110 113600 120060 113656
rect 189398 113628 189458 114139
rect 118049 113598 120060 113600
rect 118049 113595 118115 113598
rect 580073 112842 580139 112845
rect 583520 112842 584960 112932
rect 580073 112840 584960 112842
rect 580073 112784 580078 112840
rect 580134 112784 584960 112840
rect 580073 112782 584960 112784
rect 580073 112779 580139 112782
rect 583520 112692 584960 112782
rect 118785 112162 118851 112165
rect 193121 112162 193187 112165
rect 118785 112160 120060 112162
rect 118785 112104 118790 112160
rect 118846 112104 120060 112160
rect 118785 112102 120060 112104
rect 189796 112160 193187 112162
rect 189796 112104 193126 112160
rect 193182 112104 193187 112160
rect 189796 112102 193187 112104
rect 118785 112099 118851 112102
rect 193121 112099 193187 112102
rect -960 110666 480 110756
rect 3325 110666 3391 110669
rect -960 110664 3391 110666
rect -960 110608 3330 110664
rect 3386 110608 3391 110664
rect -960 110606 3391 110608
rect -960 110516 480 110606
rect 3325 110603 3391 110606
rect 118877 110666 118943 110669
rect 193121 110666 193187 110669
rect 118877 110664 120060 110666
rect 118877 110608 118882 110664
rect 118938 110608 120060 110664
rect 118877 110606 120060 110608
rect 189796 110664 193187 110666
rect 189796 110608 193126 110664
rect 193182 110608 193187 110664
rect 189796 110606 193187 110608
rect 118877 110603 118943 110606
rect 193121 110603 193187 110606
rect 119245 109170 119311 109173
rect 193029 109170 193095 109173
rect 119245 109168 120060 109170
rect 119245 109112 119250 109168
rect 119306 109112 120060 109168
rect 119245 109110 120060 109112
rect 189796 109168 193095 109170
rect 189796 109112 193034 109168
rect 193090 109112 193095 109168
rect 189796 109110 193095 109112
rect 119245 109107 119311 109110
rect 193029 109107 193095 109110
rect 119153 107674 119219 107677
rect 193029 107674 193095 107677
rect 119153 107672 120060 107674
rect 119153 107616 119158 107672
rect 119214 107616 120060 107672
rect 119153 107614 120060 107616
rect 189796 107672 193095 107674
rect 189796 107616 193034 107672
rect 193090 107616 193095 107672
rect 189796 107614 193095 107616
rect 119153 107611 119219 107614
rect 193029 107611 193095 107614
rect 119061 106178 119127 106181
rect 193121 106178 193187 106181
rect 119061 106176 120060 106178
rect 119061 106120 119066 106176
rect 119122 106120 120060 106176
rect 119061 106118 120060 106120
rect 189796 106176 193187 106178
rect 189796 106120 193126 106176
rect 193182 106120 193187 106176
rect 189796 106118 193187 106120
rect 119061 106115 119127 106118
rect 193121 106115 193187 106118
rect 118969 104682 119035 104685
rect 193121 104682 193187 104685
rect 118969 104680 120060 104682
rect 118969 104624 118974 104680
rect 119030 104624 120060 104680
rect 118969 104622 120060 104624
rect 189796 104680 193187 104682
rect 189796 104624 193126 104680
rect 193182 104624 193187 104680
rect 189796 104622 193187 104624
rect 118969 104619 119035 104622
rect 193121 104619 193187 104622
rect 120717 103458 120783 103461
rect 120582 103456 120783 103458
rect 120582 103400 120722 103456
rect 120778 103400 120783 103456
rect 120582 103398 120783 103400
rect 120582 103156 120642 103398
rect 120717 103395 120783 103398
rect 193121 103186 193187 103189
rect 189796 103184 193187 103186
rect 189796 103128 193126 103184
rect 193182 103128 193187 103184
rect 189796 103126 193187 103128
rect 193121 103123 193187 103126
rect 118693 101690 118759 101693
rect 192201 101690 192267 101693
rect 118693 101688 120060 101690
rect 118693 101632 118698 101688
rect 118754 101632 120060 101688
rect 118693 101630 120060 101632
rect 189796 101688 192267 101690
rect 189796 101632 192206 101688
rect 192262 101632 192267 101688
rect 189796 101630 192267 101632
rect 118693 101627 118759 101630
rect 192201 101627 192267 101630
rect 120809 100738 120875 100741
rect 120582 100736 120875 100738
rect 120582 100680 120814 100736
rect 120870 100680 120875 100736
rect 120582 100678 120875 100680
rect 120582 100164 120642 100678
rect 120809 100675 120875 100678
rect 192201 100194 192267 100197
rect 189796 100192 192267 100194
rect 189796 100136 192206 100192
rect 192262 100136 192267 100192
rect 189796 100134 192267 100136
rect 192201 100131 192267 100134
rect 580901 99514 580967 99517
rect 583520 99514 584960 99604
rect 580901 99512 584960 99514
rect 580901 99456 580906 99512
rect 580962 99456 584960 99512
rect 580901 99454 584960 99456
rect 580901 99451 580967 99454
rect 583520 99364 584960 99454
rect 120901 98698 120967 98701
rect 192201 98698 192267 98701
rect 120612 98696 120967 98698
rect 120612 98640 120906 98696
rect 120962 98640 120967 98696
rect 120612 98638 120967 98640
rect 189796 98696 192267 98698
rect 189796 98640 192206 98696
rect 192262 98640 192267 98696
rect 189796 98638 192267 98640
rect 120901 98635 120967 98638
rect 192201 98635 192267 98638
rect -960 97610 480 97700
rect 3693 97610 3759 97613
rect -960 97608 3759 97610
rect -960 97552 3698 97608
rect 3754 97552 3759 97608
rect -960 97550 3759 97552
rect -960 97460 480 97550
rect 3693 97547 3759 97550
rect 120993 97202 121059 97205
rect 193121 97202 193187 97205
rect 120612 97200 121059 97202
rect 120612 97144 120998 97200
rect 121054 97144 121059 97200
rect 120612 97142 121059 97144
rect 189796 97200 193187 97202
rect 189796 97144 193126 97200
rect 193182 97144 193187 97200
rect 189796 97142 193187 97144
rect 120993 97139 121059 97142
rect 193121 97139 193187 97142
rect 118601 95706 118667 95709
rect 192661 95706 192727 95709
rect 118601 95704 120060 95706
rect 118601 95648 118606 95704
rect 118662 95648 120060 95704
rect 118601 95646 120060 95648
rect 189796 95704 192727 95706
rect 189796 95648 192666 95704
rect 192722 95648 192727 95704
rect 189796 95646 192727 95648
rect 118601 95643 118667 95646
rect 192661 95643 192727 95646
rect 118509 94210 118575 94213
rect 193121 94210 193187 94213
rect 118509 94208 120060 94210
rect 118509 94152 118514 94208
rect 118570 94152 120060 94208
rect 118509 94150 120060 94152
rect 189796 94208 193187 94210
rect 189796 94152 193126 94208
rect 193182 94152 193187 94208
rect 189796 94150 193187 94152
rect 118509 94147 118575 94150
rect 193121 94147 193187 94150
rect 118417 92714 118483 92717
rect 193121 92714 193187 92717
rect 118417 92712 120060 92714
rect 118417 92656 118422 92712
rect 118478 92656 120060 92712
rect 118417 92654 120060 92656
rect 189796 92712 193187 92714
rect 189796 92656 193126 92712
rect 193182 92656 193187 92712
rect 189796 92654 193187 92656
rect 118417 92651 118483 92654
rect 193121 92651 193187 92654
rect 118325 91218 118391 91221
rect 193121 91218 193187 91221
rect 118325 91216 120060 91218
rect 118325 91160 118330 91216
rect 118386 91160 120060 91216
rect 118325 91158 120060 91160
rect 189796 91216 193187 91218
rect 189796 91160 193126 91216
rect 193182 91160 193187 91216
rect 189796 91158 193187 91160
rect 118325 91155 118391 91158
rect 193121 91155 193187 91158
rect 118233 89722 118299 89725
rect 193121 89722 193187 89725
rect 118233 89720 120060 89722
rect 118233 89664 118238 89720
rect 118294 89664 120060 89720
rect 118233 89662 120060 89664
rect 189796 89720 193187 89722
rect 189796 89664 193126 89720
rect 193182 89664 193187 89720
rect 189796 89662 193187 89664
rect 118233 89659 118299 89662
rect 193121 89659 193187 89662
rect 118141 88226 118207 88229
rect 193121 88226 193187 88229
rect 118141 88224 120060 88226
rect 118141 88168 118146 88224
rect 118202 88168 120060 88224
rect 118141 88166 120060 88168
rect 189796 88224 193187 88226
rect 189796 88168 193126 88224
rect 193182 88168 193187 88224
rect 189796 88166 193187 88168
rect 118141 88163 118207 88166
rect 193121 88163 193187 88166
rect 118417 86730 118483 86733
rect 193121 86730 193187 86733
rect 118417 86728 120060 86730
rect 118417 86672 118422 86728
rect 118478 86672 120060 86728
rect 118417 86670 120060 86672
rect 189796 86728 193187 86730
rect 189796 86672 193126 86728
rect 193182 86672 193187 86728
rect 189796 86670 193187 86672
rect 118417 86667 118483 86670
rect 193121 86667 193187 86670
rect 579981 86186 580047 86189
rect 583520 86186 584960 86276
rect 579981 86184 584960 86186
rect 579981 86128 579986 86184
rect 580042 86128 584960 86184
rect 579981 86126 584960 86128
rect 579981 86123 580047 86126
rect 583520 86036 584960 86126
rect 118601 85234 118667 85237
rect 193121 85234 193187 85237
rect 118601 85232 120060 85234
rect 118601 85176 118606 85232
rect 118662 85176 120060 85232
rect 118601 85174 120060 85176
rect 189796 85232 193187 85234
rect 189796 85176 193126 85232
rect 193182 85176 193187 85232
rect 189796 85174 193187 85176
rect 118601 85171 118667 85174
rect 193121 85171 193187 85174
rect -960 84690 480 84780
rect 3693 84690 3759 84693
rect -960 84688 3759 84690
rect -960 84632 3698 84688
rect 3754 84632 3759 84688
rect -960 84630 3759 84632
rect -960 84540 480 84630
rect 3693 84627 3759 84630
rect 118509 83738 118575 83741
rect 192661 83738 192727 83741
rect 118509 83736 120060 83738
rect 118509 83680 118514 83736
rect 118570 83680 120060 83736
rect 118509 83678 120060 83680
rect 189796 83736 192727 83738
rect 189796 83680 192666 83736
rect 192722 83680 192727 83736
rect 189796 83678 192727 83680
rect 118509 83675 118575 83678
rect 192661 83675 192727 83678
rect 118325 82242 118391 82245
rect 192845 82242 192911 82245
rect 118325 82240 120060 82242
rect 118325 82184 118330 82240
rect 118386 82184 120060 82240
rect 118325 82182 120060 82184
rect 189796 82240 192911 82242
rect 189796 82184 192850 82240
rect 192906 82184 192911 82240
rect 189796 82182 192911 82184
rect 118325 82179 118391 82182
rect 192845 82179 192911 82182
rect 118417 81154 118483 81157
rect 580165 81154 580231 81157
rect 118417 81152 580231 81154
rect 118417 81096 118422 81152
rect 118478 81096 580170 81152
rect 580226 81096 580231 81152
rect 118417 81094 580231 81096
rect 118417 81091 118483 81094
rect 580165 81091 580231 81094
rect 176694 80956 176700 81020
rect 176764 81018 176770 81020
rect 196893 81018 196959 81021
rect 176764 81016 196959 81018
rect 176764 80960 196898 81016
rect 196954 80960 196959 81016
rect 176764 80958 196959 80960
rect 176764 80956 176770 80958
rect 196893 80955 196959 80958
rect 176878 80820 176884 80884
rect 176948 80882 176954 80884
rect 580809 80882 580875 80885
rect 176948 80880 580875 80882
rect 176948 80824 580814 80880
rect 580870 80824 580875 80880
rect 176948 80822 580875 80824
rect 176948 80820 176954 80822
rect 580809 80819 580875 80822
rect 179597 80746 179663 80749
rect 580625 80746 580691 80749
rect 179597 80744 580691 80746
rect 179597 80688 179602 80744
rect 179658 80688 580630 80744
rect 580686 80688 580691 80744
rect 179597 80686 580691 80688
rect 179597 80683 179663 80686
rect 580625 80683 580691 80686
rect 177430 80548 177436 80612
rect 177500 80610 177506 80612
rect 196709 80610 196775 80613
rect 177500 80608 196775 80610
rect 177500 80552 196714 80608
rect 196770 80552 196775 80608
rect 177500 80550 196775 80552
rect 177500 80548 177506 80550
rect 196709 80547 196775 80550
rect 175222 80412 175228 80476
rect 175292 80474 175298 80476
rect 179873 80474 179939 80477
rect 175292 80472 179939 80474
rect 175292 80416 179878 80472
rect 179934 80416 179939 80472
rect 175292 80414 179939 80416
rect 175292 80412 175298 80414
rect 179873 80411 179939 80414
rect 180057 80338 180123 80341
rect 176518 80336 180123 80338
rect 176518 80280 180062 80336
rect 180118 80280 180123 80336
rect 176518 80278 180123 80280
rect 134006 80140 134012 80204
rect 134076 80140 134082 80204
rect 143206 80140 143212 80204
rect 143276 80202 143282 80204
rect 143276 80142 143550 80202
rect 143276 80140 143282 80142
rect 133270 80066 133276 80068
rect 132496 80006 133276 80066
rect 131251 79962 131317 79967
rect 131711 79964 131777 79967
rect 131251 79906 131256 79962
rect 131312 79930 131317 79962
rect 131576 79962 131777 79964
rect 131430 79930 131436 79932
rect 131312 79906 131436 79930
rect 131251 79901 131436 79906
rect 131254 79870 131436 79901
rect 131430 79868 131436 79870
rect 131500 79868 131506 79932
rect 131576 79906 131716 79962
rect 131772 79906 131777 79962
rect 131576 79904 131777 79906
rect 131389 79796 131455 79797
rect 131389 79794 131436 79796
rect 131344 79792 131436 79794
rect 131344 79736 131394 79792
rect 131344 79734 131436 79736
rect 131389 79732 131436 79734
rect 131500 79732 131506 79796
rect 131389 79731 131455 79732
rect 131389 79658 131455 79661
rect 131576 79658 131636 79904
rect 131711 79901 131777 79904
rect 131895 79930 131961 79933
rect 131895 79928 132188 79930
rect 131895 79872 131900 79928
rect 131956 79872 132188 79928
rect 131895 79870 132188 79872
rect 131895 79867 131961 79870
rect 131389 79656 131636 79658
rect 131389 79600 131394 79656
rect 131450 79600 131636 79656
rect 131389 79598 131636 79600
rect 131849 79658 131915 79661
rect 132128 79658 132188 79870
rect 132496 79797 132556 80006
rect 133270 80004 133276 80006
rect 133340 80004 133346 80068
rect 134014 79967 134074 80140
rect 143490 79967 143550 80142
rect 149646 80140 149652 80204
rect 149716 80202 149722 80204
rect 149716 80142 150266 80202
rect 149716 80140 149722 80142
rect 150206 79967 150266 80142
rect 170622 80140 170628 80204
rect 170692 80202 170698 80204
rect 170692 80142 171150 80202
rect 170692 80140 170698 80142
rect 161238 80004 161244 80068
rect 161308 80066 161314 80068
rect 161308 80004 161352 80066
rect 166758 80004 166764 80068
rect 166828 80066 166834 80068
rect 166828 80004 166872 80066
rect 134011 79962 134077 79967
rect 134839 79964 134905 79967
rect 132723 79932 132789 79933
rect 132718 79930 132724 79932
rect 132632 79870 132724 79930
rect 132718 79868 132724 79870
rect 132788 79868 132794 79932
rect 133091 79930 133157 79933
rect 132910 79928 133157 79930
rect 132910 79872 133096 79928
rect 133152 79872 133157 79928
rect 133459 79928 133525 79933
rect 132910 79870 133157 79872
rect 132723 79867 132789 79868
rect 132496 79792 132605 79797
rect 132496 79736 132544 79792
rect 132600 79736 132605 79792
rect 132496 79734 132605 79736
rect 132539 79731 132605 79734
rect 131849 79656 132188 79658
rect 131849 79600 131854 79656
rect 131910 79600 132188 79656
rect 131849 79598 132188 79600
rect 131389 79595 131455 79598
rect 131849 79595 131915 79598
rect 132769 79522 132835 79525
rect 132910 79522 132970 79870
rect 133091 79867 133157 79870
rect 133275 79894 133341 79899
rect 133275 79838 133280 79894
rect 133336 79838 133341 79894
rect 133459 79872 133464 79928
rect 133520 79872 133525 79928
rect 134011 79906 134016 79962
rect 134072 79906 134077 79962
rect 134750 79962 134905 79964
rect 134011 79901 134077 79906
rect 134287 79930 134353 79933
rect 134558 79930 134564 79932
rect 134287 79928 134564 79930
rect 133459 79867 133525 79872
rect 134287 79872 134292 79928
rect 134348 79872 134564 79928
rect 134287 79870 134564 79872
rect 134287 79867 134353 79870
rect 134558 79868 134564 79870
rect 134628 79868 134634 79932
rect 134750 79906 134844 79962
rect 134900 79930 134905 79962
rect 135483 79962 135549 79967
rect 134900 79906 134994 79930
rect 134750 79870 134994 79906
rect 133275 79833 133341 79838
rect 133278 79658 133338 79833
rect 133462 79797 133522 79867
rect 133413 79792 133522 79797
rect 133413 79736 133418 79792
rect 133474 79736 133522 79792
rect 134103 79828 134169 79831
rect 134103 79826 134212 79828
rect 134103 79770 134108 79826
rect 134164 79796 134212 79826
rect 134164 79770 134196 79796
rect 134103 79765 134196 79770
rect 133413 79734 133522 79736
rect 134152 79734 134196 79765
rect 133413 79731 133479 79734
rect 134190 79732 134196 79734
rect 134260 79732 134266 79796
rect 134793 79794 134859 79797
rect 134750 79792 134859 79794
rect 134750 79736 134798 79792
rect 134854 79736 134859 79792
rect 134750 79731 134859 79736
rect 133638 79658 133644 79660
rect 133278 79598 133644 79658
rect 133638 79596 133644 79598
rect 133708 79596 133714 79660
rect 132769 79520 132970 79522
rect 132769 79464 132774 79520
rect 132830 79464 132970 79520
rect 132769 79462 132970 79464
rect 134750 79525 134810 79731
rect 134934 79661 134994 79870
rect 135294 79868 135300 79932
rect 135364 79930 135370 79932
rect 135483 79930 135488 79962
rect 135364 79906 135488 79930
rect 135544 79906 135549 79962
rect 135364 79901 135549 79906
rect 135667 79962 135733 79967
rect 135667 79906 135672 79962
rect 135728 79906 135733 79962
rect 135667 79901 135733 79906
rect 136403 79962 136469 79967
rect 136403 79906 136408 79962
rect 136464 79906 136469 79962
rect 136403 79901 136469 79906
rect 136679 79962 136745 79967
rect 136679 79906 136684 79962
rect 136740 79930 136745 79962
rect 138611 79962 138677 79967
rect 137502 79930 137508 79932
rect 136740 79906 137508 79930
rect 136679 79901 137508 79906
rect 135364 79870 135546 79901
rect 135364 79868 135370 79870
rect 135161 79794 135227 79797
rect 135478 79794 135484 79796
rect 135161 79792 135484 79794
rect 135161 79736 135166 79792
rect 135222 79736 135484 79792
rect 135161 79734 135484 79736
rect 135161 79731 135227 79734
rect 135478 79732 135484 79734
rect 135548 79732 135554 79796
rect 134885 79656 134994 79661
rect 134885 79600 134890 79656
rect 134946 79600 134994 79656
rect 134885 79598 134994 79600
rect 135670 79658 135730 79901
rect 136127 79828 136193 79831
rect 136127 79826 136236 79828
rect 135897 79794 135963 79797
rect 136127 79794 136132 79826
rect 135897 79792 136132 79794
rect 135897 79736 135902 79792
rect 135958 79770 136132 79792
rect 136188 79770 136236 79826
rect 135958 79736 136236 79770
rect 135897 79734 136236 79736
rect 135897 79731 135963 79734
rect 136173 79658 136239 79661
rect 135670 79656 136239 79658
rect 135670 79600 136178 79656
rect 136234 79600 136239 79656
rect 135670 79598 136239 79600
rect 134885 79595 134951 79598
rect 136173 79595 136239 79598
rect 136406 79525 136466 79901
rect 136682 79870 137508 79901
rect 137502 79868 137508 79870
rect 137572 79868 137578 79932
rect 137691 79928 137757 79933
rect 137875 79932 137941 79933
rect 137691 79872 137696 79928
rect 137752 79872 137757 79928
rect 137691 79867 137757 79872
rect 137870 79868 137876 79932
rect 137940 79930 137946 79932
rect 137940 79870 138032 79930
rect 138611 79906 138616 79962
rect 138672 79906 138677 79962
rect 138611 79901 138677 79906
rect 138795 79962 138861 79967
rect 138795 79906 138800 79962
rect 138856 79906 138861 79962
rect 138795 79901 138861 79906
rect 139071 79964 139137 79967
rect 139071 79962 139272 79964
rect 139071 79906 139076 79962
rect 139132 79906 139272 79962
rect 139071 79904 139272 79906
rect 139071 79901 139137 79904
rect 137940 79868 137946 79870
rect 137875 79867 137941 79868
rect 134750 79520 134859 79525
rect 134750 79464 134798 79520
rect 134854 79464 134859 79520
rect 134750 79462 134859 79464
rect 132769 79459 132835 79462
rect 134793 79459 134859 79462
rect 135294 79460 135300 79524
rect 135364 79522 135370 79524
rect 135437 79522 135503 79525
rect 135364 79520 135503 79522
rect 135364 79464 135442 79520
rect 135498 79464 135503 79520
rect 135364 79462 135503 79464
rect 135364 79460 135370 79462
rect 135437 79459 135503 79462
rect 136357 79520 136466 79525
rect 136357 79464 136362 79520
rect 136418 79464 136466 79520
rect 136357 79462 136466 79464
rect 137694 79525 137754 79867
rect 138614 79797 138674 79901
rect 138798 79797 138858 79901
rect 138054 79732 138060 79796
rect 138124 79794 138130 79796
rect 138197 79794 138263 79797
rect 138427 79796 138493 79797
rect 138422 79794 138428 79796
rect 138124 79792 138263 79794
rect 138124 79736 138202 79792
rect 138258 79736 138263 79792
rect 138124 79734 138263 79736
rect 138336 79734 138428 79794
rect 138124 79732 138130 79734
rect 138197 79731 138263 79734
rect 138422 79732 138428 79734
rect 138492 79732 138498 79796
rect 138565 79792 138674 79797
rect 138565 79736 138570 79792
rect 138626 79736 138674 79792
rect 138565 79734 138674 79736
rect 138749 79792 138858 79797
rect 138749 79736 138754 79792
rect 138810 79736 138858 79792
rect 138749 79734 138858 79736
rect 138427 79731 138493 79732
rect 138565 79731 138631 79734
rect 138749 79731 138815 79734
rect 137694 79520 137803 79525
rect 137694 79464 137742 79520
rect 137798 79464 137803 79520
rect 137694 79462 137803 79464
rect 136357 79459 136423 79462
rect 137737 79459 137803 79462
rect 139025 79522 139091 79525
rect 139212 79522 139272 79904
rect 139899 79962 139965 79967
rect 139899 79906 139904 79962
rect 139960 79906 139965 79962
rect 139899 79901 139965 79906
rect 140635 79962 140701 79967
rect 140635 79906 140640 79962
rect 140696 79906 140701 79962
rect 141739 79962 141805 79967
rect 140635 79901 140701 79906
rect 141371 79928 141437 79933
rect 139902 79794 139962 79901
rect 140267 79894 140333 79899
rect 140267 79838 140272 79894
rect 140328 79838 140333 79894
rect 140267 79833 140333 79838
rect 140129 79794 140195 79797
rect 139902 79792 140195 79794
rect 139902 79736 140134 79792
rect 140190 79736 140195 79792
rect 139902 79734 140195 79736
rect 140129 79731 140195 79734
rect 140270 79661 140330 79833
rect 140638 79661 140698 79901
rect 141371 79872 141376 79928
rect 141432 79872 141437 79928
rect 141371 79867 141437 79872
rect 141555 79928 141621 79933
rect 141555 79872 141560 79928
rect 141616 79872 141621 79928
rect 141739 79906 141744 79962
rect 141800 79906 141805 79962
rect 143487 79962 143553 79967
rect 141739 79901 141805 79906
rect 141555 79867 141621 79872
rect 140819 79792 140885 79797
rect 140819 79736 140824 79792
rect 140880 79736 140885 79792
rect 140819 79731 140885 79736
rect 139393 79658 139459 79661
rect 139853 79660 139919 79661
rect 139710 79658 139716 79660
rect 139393 79656 139716 79658
rect 139393 79600 139398 79656
rect 139454 79600 139716 79656
rect 139393 79598 139716 79600
rect 139393 79595 139459 79598
rect 139710 79596 139716 79598
rect 139780 79596 139786 79660
rect 139853 79656 139900 79660
rect 139964 79658 139970 79660
rect 139853 79600 139858 79656
rect 139853 79596 139900 79600
rect 139964 79598 140010 79658
rect 140270 79656 140379 79661
rect 140270 79600 140318 79656
rect 140374 79600 140379 79656
rect 140270 79598 140379 79600
rect 139964 79596 139970 79598
rect 139853 79595 139919 79596
rect 140313 79595 140379 79598
rect 140589 79656 140698 79661
rect 140589 79600 140594 79656
rect 140650 79600 140698 79656
rect 140589 79598 140698 79600
rect 140822 79661 140882 79731
rect 141374 79661 141434 79867
rect 140822 79656 140931 79661
rect 140822 79600 140870 79656
rect 140926 79600 140931 79656
rect 140822 79598 140931 79600
rect 140589 79595 140655 79598
rect 140865 79595 140931 79598
rect 141325 79656 141434 79661
rect 141325 79600 141330 79656
rect 141386 79600 141434 79656
rect 141325 79598 141434 79600
rect 141325 79595 141391 79598
rect 141558 79525 141618 79867
rect 141742 79797 141802 79901
rect 141918 79868 141924 79932
rect 141988 79930 141994 79932
rect 142291 79930 142357 79933
rect 141988 79870 142046 79930
rect 142291 79928 142952 79930
rect 142291 79872 142296 79928
rect 142352 79872 142952 79928
rect 142291 79870 142952 79872
rect 141988 79868 141994 79870
rect 141923 79838 141928 79868
rect 141984 79838 141989 79868
rect 142291 79867 142357 79870
rect 141923 79833 141989 79838
rect 142892 79797 142952 79870
rect 143027 79928 143093 79933
rect 143027 79872 143032 79928
rect 143088 79872 143093 79928
rect 143027 79867 143093 79872
rect 143303 79930 143369 79933
rect 143303 79928 143412 79930
rect 143303 79872 143308 79928
rect 143364 79872 143412 79928
rect 143487 79906 143492 79962
rect 143548 79906 143553 79962
rect 144407 79964 144473 79967
rect 144407 79962 144516 79964
rect 143763 79932 143829 79933
rect 143758 79930 143764 79932
rect 143487 79901 143553 79906
rect 143303 79867 143412 79872
rect 143672 79870 143764 79930
rect 143758 79868 143764 79870
rect 143828 79868 143834 79932
rect 144407 79906 144412 79962
rect 144468 79932 144516 79962
rect 148179 79962 148245 79967
rect 144468 79906 144500 79932
rect 144407 79901 144500 79906
rect 144456 79870 144500 79901
rect 144494 79868 144500 79870
rect 144564 79868 144570 79932
rect 145603 79894 145669 79899
rect 143763 79867 143829 79868
rect 141693 79792 141802 79797
rect 141693 79736 141698 79792
rect 141754 79736 141802 79792
rect 141693 79734 141802 79736
rect 142889 79792 142955 79797
rect 142889 79736 142894 79792
rect 142950 79736 142955 79792
rect 141693 79731 141759 79734
rect 142889 79731 142955 79736
rect 141785 79658 141851 79661
rect 142102 79658 142108 79660
rect 141785 79656 142108 79658
rect 141785 79600 141790 79656
rect 141846 79600 142108 79656
rect 141785 79598 142108 79600
rect 141785 79595 141851 79598
rect 142102 79596 142108 79598
rect 142172 79596 142178 79660
rect 139025 79520 139272 79522
rect 139025 79464 139030 79520
rect 139086 79464 139272 79520
rect 139025 79462 139272 79464
rect 141509 79520 141618 79525
rect 141509 79464 141514 79520
rect 141570 79464 141618 79520
rect 141509 79462 141618 79464
rect 143030 79522 143090 79867
rect 143352 79796 143412 79867
rect 145603 79838 145608 79894
rect 145664 79838 145669 79894
rect 145603 79833 145669 79838
rect 146339 79894 146405 79899
rect 146339 79838 146344 79894
rect 146400 79838 146405 79894
rect 146886 79868 146892 79932
rect 146956 79930 146962 79932
rect 147259 79930 147325 79933
rect 147995 79932 148061 79933
rect 148179 79932 148184 79962
rect 148240 79932 148245 79962
rect 150019 79962 150085 79967
rect 147990 79930 147996 79932
rect 146956 79928 147325 79930
rect 146956 79872 147264 79928
rect 147320 79872 147325 79928
rect 146956 79870 147325 79872
rect 147904 79870 147996 79930
rect 146956 79868 146962 79870
rect 147259 79867 147325 79870
rect 147990 79868 147996 79870
rect 148060 79868 148066 79932
rect 148174 79868 148180 79932
rect 148244 79930 148250 79932
rect 148639 79930 148705 79933
rect 148910 79930 148916 79932
rect 148244 79870 148302 79930
rect 148639 79928 148916 79930
rect 148639 79872 148644 79928
rect 148700 79872 148916 79928
rect 148639 79870 148916 79872
rect 148244 79868 148250 79870
rect 147995 79867 148061 79868
rect 148639 79867 148705 79870
rect 148910 79868 148916 79870
rect 148980 79868 148986 79932
rect 149283 79928 149349 79933
rect 149283 79872 149288 79928
rect 149344 79872 149349 79928
rect 149283 79867 149349 79872
rect 149651 79930 149717 79933
rect 149651 79928 149944 79930
rect 149651 79872 149656 79928
rect 149712 79872 149944 79928
rect 150019 79906 150024 79962
rect 150080 79906 150085 79962
rect 150019 79901 150085 79906
rect 150203 79962 150269 79967
rect 150203 79906 150208 79962
rect 150264 79906 150269 79962
rect 150203 79901 150269 79906
rect 150571 79962 150637 79967
rect 150571 79906 150576 79962
rect 150632 79906 150637 79962
rect 150571 79901 150637 79906
rect 150755 79962 150821 79967
rect 150755 79906 150760 79962
rect 150816 79906 150821 79962
rect 151123 79962 151189 79967
rect 150755 79901 150821 79906
rect 150939 79928 151005 79933
rect 151123 79932 151128 79962
rect 151184 79932 151189 79962
rect 151399 79964 151465 79967
rect 151399 79962 151508 79964
rect 149651 79870 149944 79872
rect 149651 79867 149717 79870
rect 146339 79833 146405 79838
rect 143352 79734 143396 79796
rect 143390 79732 143396 79734
rect 143460 79732 143466 79796
rect 143809 79794 143875 79797
rect 144039 79794 144105 79797
rect 143809 79792 144105 79794
rect 143809 79736 143814 79792
rect 143870 79736 144044 79792
rect 144100 79736 144105 79792
rect 143809 79734 144105 79736
rect 143809 79731 143875 79734
rect 144039 79731 144105 79734
rect 144591 79794 144657 79797
rect 145143 79794 145209 79797
rect 144591 79792 144700 79794
rect 144591 79736 144596 79792
rect 144652 79736 144700 79792
rect 144591 79731 144700 79736
rect 145143 79792 145482 79794
rect 145143 79736 145148 79792
rect 145204 79736 145482 79792
rect 145143 79734 145482 79736
rect 145143 79731 145209 79734
rect 143625 79658 143691 79661
rect 144453 79658 144519 79661
rect 143625 79656 144519 79658
rect 143625 79600 143630 79656
rect 143686 79600 144458 79656
rect 144514 79600 144519 79656
rect 143625 79598 144519 79600
rect 144640 79660 144700 79731
rect 144640 79598 144684 79660
rect 143625 79595 143691 79598
rect 144453 79595 144519 79598
rect 144678 79596 144684 79598
rect 144748 79596 144754 79660
rect 144913 79658 144979 79661
rect 144913 79656 145114 79658
rect 144913 79600 144918 79656
rect 144974 79600 145114 79656
rect 144913 79598 145114 79600
rect 144913 79595 144979 79598
rect 145054 79525 145114 79598
rect 143625 79522 143691 79525
rect 143030 79520 143691 79522
rect 143030 79464 143630 79520
rect 143686 79464 143691 79520
rect 143030 79462 143691 79464
rect 139025 79459 139091 79462
rect 141509 79459 141575 79462
rect 143625 79459 143691 79462
rect 145005 79520 145114 79525
rect 145005 79464 145010 79520
rect 145066 79464 145114 79520
rect 145005 79462 145114 79464
rect 145281 79522 145347 79525
rect 145422 79522 145482 79734
rect 145606 79525 145666 79833
rect 145741 79794 145807 79797
rect 145741 79792 146172 79794
rect 145741 79736 145746 79792
rect 145802 79736 146172 79792
rect 145741 79734 146172 79736
rect 145741 79731 145807 79734
rect 146112 79661 146172 79734
rect 146109 79656 146175 79661
rect 146109 79600 146114 79656
rect 146170 79600 146175 79656
rect 146109 79595 146175 79600
rect 146342 79658 146402 79833
rect 148869 79796 148935 79797
rect 148869 79794 148916 79796
rect 148824 79792 148916 79794
rect 148824 79736 148874 79792
rect 148824 79734 148916 79736
rect 148869 79732 148916 79734
rect 148980 79732 148986 79796
rect 148869 79731 148935 79732
rect 147489 79658 147555 79661
rect 146342 79656 147555 79658
rect 146342 79600 147494 79656
rect 147550 79600 147555 79656
rect 146342 79598 147555 79600
rect 149286 79658 149346 79867
rect 149697 79658 149763 79661
rect 149286 79656 149763 79658
rect 149286 79600 149702 79656
rect 149758 79600 149763 79656
rect 149286 79598 149763 79600
rect 147489 79595 147555 79598
rect 149697 79595 149763 79598
rect 145281 79520 145482 79522
rect 145281 79464 145286 79520
rect 145342 79464 145482 79520
rect 145281 79462 145482 79464
rect 145557 79520 145666 79525
rect 145557 79464 145562 79520
rect 145618 79464 145666 79520
rect 145557 79462 145666 79464
rect 149053 79522 149119 79525
rect 149605 79522 149671 79525
rect 149053 79520 149671 79522
rect 149053 79464 149058 79520
rect 149114 79464 149610 79520
rect 149666 79464 149671 79520
rect 149053 79462 149671 79464
rect 149884 79522 149944 79870
rect 150022 79661 150082 79901
rect 150157 79796 150223 79797
rect 150157 79792 150204 79796
rect 150268 79794 150274 79796
rect 150157 79736 150162 79792
rect 150157 79732 150204 79736
rect 150268 79734 150314 79794
rect 150268 79732 150274 79734
rect 150157 79731 150223 79732
rect 150022 79656 150131 79661
rect 150022 79600 150070 79656
rect 150126 79600 150131 79656
rect 150022 79598 150131 79600
rect 150574 79658 150634 79901
rect 150758 79797 150818 79901
rect 150939 79872 150944 79928
rect 151000 79872 151005 79928
rect 150939 79867 151005 79872
rect 151118 79868 151124 79932
rect 151188 79930 151194 79932
rect 151188 79870 151246 79930
rect 151399 79906 151404 79962
rect 151460 79932 151508 79962
rect 151675 79962 151741 79967
rect 151675 79932 151680 79962
rect 151736 79932 151741 79962
rect 153331 79962 153397 79967
rect 151460 79906 151492 79932
rect 151399 79901 151492 79906
rect 151448 79870 151492 79901
rect 151188 79868 151194 79870
rect 151486 79868 151492 79870
rect 151556 79868 151562 79932
rect 151670 79868 151676 79932
rect 151740 79930 151746 79932
rect 152503 79930 152569 79933
rect 151740 79870 151798 79930
rect 152230 79928 152569 79930
rect 152230 79872 152508 79928
rect 152564 79872 152569 79928
rect 152230 79870 152569 79872
rect 151740 79868 151746 79870
rect 150758 79792 150867 79797
rect 150758 79736 150806 79792
rect 150862 79736 150867 79792
rect 150758 79734 150867 79736
rect 150801 79731 150867 79734
rect 150801 79658 150867 79661
rect 150574 79656 150867 79658
rect 150574 79600 150806 79656
rect 150862 79600 150867 79656
rect 150574 79598 150867 79600
rect 150942 79658 151002 79867
rect 151302 79732 151308 79796
rect 151372 79794 151378 79796
rect 151813 79794 151879 79797
rect 151372 79792 151879 79794
rect 151372 79736 151818 79792
rect 151874 79736 151879 79792
rect 151372 79734 151879 79736
rect 151372 79732 151378 79734
rect 151813 79731 151879 79734
rect 151629 79658 151695 79661
rect 150942 79656 151695 79658
rect 150942 79600 151634 79656
rect 151690 79600 151695 79656
rect 150942 79598 151695 79600
rect 150065 79595 150131 79598
rect 150801 79595 150867 79598
rect 151629 79595 151695 79598
rect 151813 79658 151879 79661
rect 152230 79658 152290 79870
rect 152503 79867 152569 79870
rect 152774 79868 152780 79932
rect 152844 79930 152850 79932
rect 153055 79930 153121 79933
rect 152844 79928 153121 79930
rect 152844 79872 153060 79928
rect 153116 79872 153121 79928
rect 153331 79906 153336 79962
rect 153392 79906 153397 79962
rect 153699 79962 153765 79967
rect 153331 79901 153397 79906
rect 153515 79928 153581 79933
rect 153699 79932 153704 79962
rect 153760 79932 153765 79962
rect 154159 79964 154225 79967
rect 154159 79962 154268 79964
rect 152844 79870 153121 79872
rect 152844 79868 152850 79870
rect 153055 79867 153121 79870
rect 153334 79797 153394 79901
rect 153515 79872 153520 79928
rect 153576 79872 153581 79928
rect 153515 79867 153581 79872
rect 153694 79868 153700 79932
rect 153764 79930 153770 79932
rect 153764 79870 153822 79930
rect 154159 79906 154164 79962
rect 154220 79930 154268 79962
rect 155815 79962 155881 79967
rect 154619 79932 154685 79933
rect 154430 79930 154436 79932
rect 154220 79906 154436 79930
rect 154159 79901 154436 79906
rect 154208 79870 154436 79901
rect 153764 79868 153770 79870
rect 154430 79868 154436 79870
rect 154500 79868 154506 79932
rect 154614 79868 154620 79932
rect 154684 79930 154690 79932
rect 155079 79930 155145 79933
rect 155350 79930 155356 79932
rect 154684 79870 154776 79930
rect 155079 79928 155356 79930
rect 155079 79872 155084 79928
rect 155140 79872 155356 79928
rect 155079 79870 155356 79872
rect 154684 79868 154690 79870
rect 154619 79867 154685 79868
rect 155079 79867 155145 79870
rect 155350 79868 155356 79870
rect 155420 79868 155426 79932
rect 155534 79868 155540 79932
rect 155604 79930 155610 79932
rect 155815 79930 155820 79962
rect 155604 79906 155820 79930
rect 155876 79906 155881 79962
rect 157103 79962 157169 79967
rect 155604 79901 155881 79906
rect 155604 79870 155878 79901
rect 155604 79868 155610 79870
rect 156270 79868 156276 79932
rect 156340 79930 156346 79932
rect 156551 79930 156617 79933
rect 156340 79928 156617 79930
rect 156340 79872 156556 79928
rect 156612 79872 156617 79928
rect 156340 79870 156617 79872
rect 156340 79868 156346 79870
rect 156551 79867 156617 79870
rect 156822 79868 156828 79932
rect 156892 79930 156898 79932
rect 157103 79930 157108 79962
rect 156892 79906 157108 79930
rect 157164 79906 157169 79962
rect 158299 79962 158365 79967
rect 157839 79930 157905 79933
rect 156892 79901 157169 79906
rect 157796 79928 157905 79930
rect 156892 79870 157166 79901
rect 157796 79872 157844 79928
rect 157900 79872 157905 79928
rect 156892 79868 156898 79870
rect 157796 79867 157905 79872
rect 158110 79868 158116 79932
rect 158180 79930 158186 79932
rect 158299 79930 158304 79962
rect 158180 79906 158304 79930
rect 158360 79906 158365 79962
rect 158180 79901 158365 79906
rect 158575 79930 158641 79933
rect 159311 79930 159377 79933
rect 159582 79930 159588 79932
rect 158575 79928 158684 79930
rect 158180 79870 158362 79901
rect 158575 79872 158580 79928
rect 158636 79872 158684 79928
rect 158180 79868 158186 79870
rect 158575 79867 158684 79872
rect 159311 79928 159588 79930
rect 159311 79872 159316 79928
rect 159372 79872 159588 79928
rect 159311 79870 159588 79872
rect 159311 79867 159377 79870
rect 159582 79868 159588 79870
rect 159652 79868 159658 79932
rect 160231 79930 160297 79933
rect 160686 79930 160692 79932
rect 160231 79928 160692 79930
rect 159955 79894 160021 79899
rect 153334 79792 153443 79797
rect 153334 79736 153382 79792
rect 153438 79736 153443 79792
rect 153334 79734 153443 79736
rect 153377 79731 153443 79734
rect 151813 79656 152290 79658
rect 151813 79600 151818 79656
rect 151874 79600 152290 79656
rect 151813 79598 152290 79600
rect 153518 79658 153578 79867
rect 154062 79732 154068 79796
rect 154132 79794 154138 79796
rect 154527 79794 154593 79797
rect 155355 79794 155421 79797
rect 154132 79792 154593 79794
rect 154132 79736 154532 79792
rect 154588 79736 154593 79792
rect 154132 79734 154593 79736
rect 154132 79732 154138 79734
rect 154527 79731 154593 79734
rect 155036 79792 155421 79794
rect 155036 79736 155360 79792
rect 155416 79736 155421 79792
rect 155036 79734 155421 79736
rect 155036 79661 155096 79734
rect 155355 79731 155421 79734
rect 156137 79794 156203 79797
rect 156873 79794 156939 79797
rect 156137 79792 156939 79794
rect 156137 79736 156142 79792
rect 156198 79736 156878 79792
rect 156934 79736 156939 79792
rect 156137 79734 156939 79736
rect 157796 79794 157856 79867
rect 157796 79734 157994 79794
rect 156137 79731 156203 79734
rect 156873 79731 156939 79734
rect 153837 79658 153903 79661
rect 153518 79656 153903 79658
rect 153518 79600 153842 79656
rect 153898 79600 153903 79656
rect 153518 79598 153903 79600
rect 151813 79595 151879 79598
rect 153837 79595 153903 79598
rect 155033 79656 155099 79661
rect 155033 79600 155038 79656
rect 155094 79600 155099 79656
rect 155033 79595 155099 79600
rect 156229 79658 156295 79661
rect 156505 79658 156571 79661
rect 156229 79656 156571 79658
rect 156229 79600 156234 79656
rect 156290 79600 156510 79656
rect 156566 79600 156571 79656
rect 156229 79598 156571 79600
rect 156229 79595 156295 79598
rect 156505 79595 156571 79598
rect 150249 79522 150315 79525
rect 149884 79520 150315 79522
rect 149884 79464 150254 79520
rect 150310 79464 150315 79520
rect 149884 79462 150315 79464
rect 145005 79459 145071 79462
rect 145281 79459 145347 79462
rect 145557 79459 145623 79462
rect 149053 79459 149119 79462
rect 149605 79459 149671 79462
rect 150249 79459 150315 79462
rect 154849 79522 154915 79525
rect 155125 79522 155191 79525
rect 154849 79520 155191 79522
rect 154849 79464 154854 79520
rect 154910 79464 155130 79520
rect 155186 79464 155191 79520
rect 154849 79462 155191 79464
rect 154849 79459 154915 79462
rect 155125 79459 155191 79462
rect 155401 79522 155467 79525
rect 155769 79522 155835 79525
rect 155401 79520 155835 79522
rect 155401 79464 155406 79520
rect 155462 79464 155774 79520
rect 155830 79464 155835 79520
rect 155401 79462 155835 79464
rect 155401 79459 155467 79462
rect 155769 79459 155835 79462
rect 156689 79522 156755 79525
rect 157190 79522 157196 79524
rect 156689 79520 157196 79522
rect 156689 79464 156694 79520
rect 156750 79464 157196 79520
rect 156689 79462 157196 79464
rect 156689 79459 156755 79462
rect 157190 79460 157196 79462
rect 157260 79460 157266 79524
rect 157333 79522 157399 79525
rect 157934 79522 157994 79734
rect 158294 79732 158300 79796
rect 158364 79794 158370 79796
rect 158624 79794 158684 79867
rect 159955 79838 159960 79894
rect 160016 79838 160021 79894
rect 160231 79872 160236 79928
rect 160292 79872 160692 79928
rect 160231 79870 160692 79872
rect 160231 79867 160297 79870
rect 160686 79868 160692 79870
rect 160756 79868 160762 79932
rect 161151 79930 161217 79933
rect 161292 79930 161352 80004
rect 162715 79962 162781 79967
rect 161151 79928 161352 79930
rect 161151 79872 161156 79928
rect 161212 79872 161352 79928
rect 161151 79870 161352 79872
rect 161519 79930 161585 79933
rect 161974 79930 161980 79932
rect 161519 79928 161980 79930
rect 161519 79872 161524 79928
rect 161580 79872 161980 79928
rect 161519 79870 161980 79872
rect 161151 79867 161217 79870
rect 161519 79867 161585 79870
rect 161974 79868 161980 79870
rect 162044 79868 162050 79932
rect 162163 79928 162229 79933
rect 162163 79872 162168 79928
rect 162224 79872 162229 79928
rect 162163 79867 162229 79872
rect 162342 79868 162348 79932
rect 162412 79930 162418 79932
rect 162715 79930 162720 79962
rect 162412 79906 162720 79930
rect 162776 79906 162781 79962
rect 165935 79962 166001 79967
rect 162412 79901 162781 79906
rect 162412 79870 162778 79901
rect 162412 79868 162418 79870
rect 163262 79868 163268 79932
rect 163332 79930 163338 79932
rect 163332 79899 164250 79930
rect 163332 79894 164253 79899
rect 163332 79870 164192 79894
rect 163332 79868 163338 79870
rect 159955 79833 160021 79838
rect 158364 79734 158684 79794
rect 158364 79732 158370 79734
rect 158846 79596 158852 79660
rect 158916 79658 158922 79660
rect 159958 79658 160018 79833
rect 161054 79732 161060 79796
rect 161124 79794 161130 79796
rect 161197 79794 161263 79797
rect 161124 79792 161263 79794
rect 161124 79736 161202 79792
rect 161258 79736 161263 79792
rect 161124 79734 161263 79736
rect 161124 79732 161130 79734
rect 161197 79731 161263 79734
rect 158916 79598 160018 79658
rect 161841 79658 161907 79661
rect 162166 79658 162226 79867
rect 164187 79838 164192 79870
rect 164248 79838 164253 79894
rect 164734 79868 164740 79932
rect 164804 79930 164810 79932
rect 165015 79930 165081 79933
rect 165567 79930 165633 79933
rect 164804 79928 165081 79930
rect 164804 79872 165020 79928
rect 165076 79872 165081 79928
rect 164804 79870 165081 79872
rect 164804 79868 164810 79870
rect 165015 79867 165081 79870
rect 165248 79928 165633 79930
rect 165248 79872 165572 79928
rect 165628 79872 165633 79928
rect 165935 79906 165940 79962
rect 165996 79906 166001 79962
rect 165935 79901 166001 79906
rect 166671 79930 166737 79933
rect 166812 79930 166872 80004
rect 168971 79962 169037 79967
rect 167315 79932 167381 79933
rect 168051 79932 168117 79933
rect 167310 79930 167316 79932
rect 166671 79928 166872 79930
rect 165248 79870 165633 79872
rect 164187 79833 164253 79838
rect 163727 79794 163793 79797
rect 163998 79794 164004 79796
rect 163727 79792 164004 79794
rect 163727 79736 163732 79792
rect 163788 79736 164004 79792
rect 163727 79734 164004 79736
rect 163727 79731 163793 79734
rect 163998 79732 164004 79734
rect 164068 79732 164074 79796
rect 165102 79732 165108 79796
rect 165172 79794 165178 79796
rect 165248 79794 165308 79870
rect 165567 79867 165633 79870
rect 165521 79796 165587 79797
rect 165470 79794 165476 79796
rect 165172 79734 165308 79794
rect 165430 79734 165476 79794
rect 165540 79792 165587 79796
rect 165582 79736 165587 79792
rect 165172 79732 165178 79734
rect 165470 79732 165476 79734
rect 165540 79732 165587 79736
rect 165521 79731 165587 79732
rect 161841 79656 162226 79658
rect 161841 79600 161846 79656
rect 161902 79600 162226 79656
rect 161841 79598 162226 79600
rect 165938 79658 165998 79901
rect 166671 79872 166676 79928
rect 166732 79872 166872 79928
rect 166671 79870 166872 79872
rect 167224 79870 167316 79930
rect 166671 79867 166737 79870
rect 167310 79868 167316 79870
rect 167380 79868 167386 79932
rect 168046 79930 168052 79932
rect 167960 79870 168052 79930
rect 168046 79868 168052 79870
rect 168116 79868 168122 79932
rect 168235 79928 168301 79933
rect 168787 79930 168853 79933
rect 168971 79932 168976 79962
rect 169032 79932 169037 79962
rect 170259 79962 170325 79967
rect 170535 79964 170601 79967
rect 170903 79964 170969 79967
rect 170259 79932 170264 79962
rect 170320 79932 170325 79962
rect 170492 79962 170601 79964
rect 168235 79872 168240 79928
rect 168296 79872 168301 79928
rect 167315 79867 167381 79868
rect 168051 79867 168117 79868
rect 168235 79867 168301 79872
rect 168606 79928 168853 79930
rect 168606 79872 168792 79928
rect 168848 79872 168853 79928
rect 168606 79870 168853 79872
rect 166579 79792 166645 79797
rect 166579 79736 166584 79792
rect 166640 79736 166645 79792
rect 166579 79731 166645 79736
rect 167678 79732 167684 79796
rect 167748 79794 167754 79796
rect 168238 79794 168298 79867
rect 167748 79734 168298 79794
rect 167748 79732 167754 79734
rect 166582 79661 166642 79731
rect 166349 79658 166415 79661
rect 165938 79656 166415 79658
rect 165938 79600 166354 79656
rect 166410 79600 166415 79656
rect 165938 79598 166415 79600
rect 158916 79596 158922 79598
rect 161841 79595 161907 79598
rect 166349 79595 166415 79598
rect 166533 79656 166642 79661
rect 166533 79600 166538 79656
rect 166594 79600 166642 79656
rect 166533 79598 166642 79600
rect 168606 79661 168666 79870
rect 168787 79867 168853 79870
rect 168966 79868 168972 79932
rect 169036 79930 169042 79932
rect 169036 79870 169094 79930
rect 169523 79894 169589 79899
rect 169036 79868 169042 79870
rect 169523 79838 169528 79894
rect 169584 79838 169589 79894
rect 170254 79868 170260 79932
rect 170324 79930 170330 79932
rect 170324 79870 170382 79930
rect 170492 79906 170540 79962
rect 170596 79906 170601 79962
rect 170860 79962 170969 79964
rect 170719 79930 170785 79933
rect 170492 79901 170601 79906
rect 170676 79928 170785 79930
rect 170324 79868 170330 79870
rect 169523 79833 169589 79838
rect 168833 79792 168899 79797
rect 168833 79736 168838 79792
rect 168894 79736 168899 79792
rect 168833 79731 168899 79736
rect 168606 79656 168715 79661
rect 168606 79600 168654 79656
rect 168710 79600 168715 79656
rect 168606 79598 168715 79600
rect 166533 79595 166599 79598
rect 168649 79595 168715 79598
rect 168836 79525 168896 79731
rect 169526 79661 169586 79833
rect 170492 79661 170552 79901
rect 170676 79872 170724 79928
rect 170780 79872 170785 79928
rect 170676 79867 170785 79872
rect 170860 79906 170908 79962
rect 170964 79906 170969 79962
rect 171090 79933 171150 80142
rect 171542 80004 171548 80068
rect 171612 80066 171618 80068
rect 171612 80006 171978 80066
rect 171612 80004 171618 80006
rect 170860 79901 170969 79906
rect 171087 79928 171153 79933
rect 171731 79932 171797 79933
rect 171726 79930 171732 79932
rect 169526 79656 169635 79661
rect 169526 79600 169574 79656
rect 169630 79600 169635 79656
rect 169526 79598 169635 79600
rect 169569 79595 169635 79598
rect 170489 79656 170555 79661
rect 170489 79600 170494 79656
rect 170550 79600 170555 79656
rect 170489 79595 170555 79600
rect 170676 79658 170736 79867
rect 170860 79796 170920 79901
rect 171087 79872 171092 79928
rect 171148 79872 171153 79928
rect 171087 79867 171153 79872
rect 171640 79870 171732 79930
rect 171726 79868 171732 79870
rect 171796 79868 171802 79932
rect 171918 79930 171978 80006
rect 176518 79967 176578 80278
rect 180057 80275 180123 80278
rect 177798 80140 177804 80204
rect 177868 80202 177874 80204
rect 180701 80202 180767 80205
rect 177868 80200 180767 80202
rect 177868 80144 180706 80200
rect 180762 80144 180767 80200
rect 177868 80142 180767 80144
rect 177868 80140 177874 80142
rect 180701 80139 180767 80142
rect 180241 80066 180307 80069
rect 177070 80064 180307 80066
rect 177070 80008 180246 80064
rect 180302 80008 180307 80064
rect 177070 80006 180307 80008
rect 173571 79962 173637 79967
rect 172467 79930 172533 79933
rect 172651 79932 172717 79933
rect 171918 79928 172533 79930
rect 171918 79872 172472 79928
rect 172528 79872 172533 79928
rect 171918 79870 172533 79872
rect 171731 79867 171797 79868
rect 172467 79867 172533 79870
rect 172646 79868 172652 79932
rect 172716 79930 172722 79932
rect 172927 79930 172993 79933
rect 173198 79930 173204 79932
rect 172716 79870 172808 79930
rect 172927 79928 173204 79930
rect 172927 79872 172932 79928
rect 172988 79872 173204 79928
rect 172927 79870 173204 79872
rect 172716 79868 172722 79870
rect 172651 79867 172717 79868
rect 172927 79867 172993 79870
rect 173198 79868 173204 79870
rect 173268 79868 173274 79932
rect 173571 79906 173576 79962
rect 173632 79930 173637 79962
rect 174031 79964 174097 79967
rect 174031 79962 174370 79964
rect 173632 79906 173772 79930
rect 173571 79901 173772 79906
rect 174031 79906 174036 79962
rect 174092 79906 174370 79962
rect 176515 79962 176581 79967
rect 174031 79904 174370 79906
rect 174031 79901 174097 79904
rect 173574 79870 173772 79901
rect 170806 79732 170812 79796
rect 170876 79734 170920 79796
rect 171639 79794 171705 79797
rect 172375 79794 172441 79797
rect 171639 79792 171748 79794
rect 171639 79736 171644 79792
rect 171700 79736 171748 79792
rect 170876 79732 170882 79734
rect 171639 79731 171748 79736
rect 171688 79661 171748 79731
rect 172240 79792 172441 79794
rect 172240 79736 172380 79792
rect 172436 79736 172441 79792
rect 172240 79734 172441 79736
rect 170857 79658 170923 79661
rect 170676 79656 170923 79658
rect 170676 79600 170862 79656
rect 170918 79600 170923 79656
rect 170676 79598 170923 79600
rect 170857 79595 170923 79598
rect 171317 79656 171383 79661
rect 171317 79600 171322 79656
rect 171378 79600 171383 79656
rect 171317 79595 171383 79600
rect 171685 79656 171751 79661
rect 171685 79600 171690 79656
rect 171746 79600 171751 79656
rect 171685 79595 171751 79600
rect 172094 79596 172100 79660
rect 172164 79658 172170 79660
rect 172240 79658 172300 79734
rect 172375 79731 172441 79734
rect 172973 79794 173039 79797
rect 172973 79792 173082 79794
rect 172973 79736 172978 79792
rect 173034 79736 173082 79792
rect 172973 79731 173082 79736
rect 173382 79732 173388 79796
rect 173452 79794 173458 79796
rect 173525 79794 173591 79797
rect 173452 79792 173591 79794
rect 173452 79736 173530 79792
rect 173586 79736 173591 79792
rect 173452 79734 173591 79736
rect 173452 79732 173458 79734
rect 173525 79731 173591 79734
rect 173022 79661 173082 79731
rect 172164 79598 172300 79658
rect 172973 79656 173082 79661
rect 172973 79600 172978 79656
rect 173034 79600 173082 79656
rect 172973 79598 173082 79600
rect 173157 79658 173223 79661
rect 173525 79658 173591 79661
rect 173157 79656 173591 79658
rect 173157 79600 173162 79656
rect 173218 79600 173530 79656
rect 173586 79600 173591 79656
rect 173157 79598 173591 79600
rect 172164 79596 172170 79598
rect 172973 79595 173039 79598
rect 173157 79595 173223 79598
rect 173525 79595 173591 79598
rect 157333 79520 157994 79522
rect 157333 79464 157338 79520
rect 157394 79464 157994 79520
rect 157333 79462 157994 79464
rect 157333 79459 157399 79462
rect 159582 79460 159588 79524
rect 159652 79522 159658 79524
rect 159909 79522 159975 79525
rect 159652 79520 159975 79522
rect 159652 79464 159914 79520
rect 159970 79464 159975 79520
rect 159652 79462 159975 79464
rect 159652 79460 159658 79462
rect 159909 79459 159975 79462
rect 160870 79460 160876 79524
rect 160940 79522 160946 79524
rect 161289 79522 161355 79525
rect 160940 79520 161355 79522
rect 160940 79464 161294 79520
rect 161350 79464 161355 79520
rect 160940 79462 161355 79464
rect 160940 79460 160946 79462
rect 161289 79459 161355 79462
rect 164325 79522 164391 79525
rect 164550 79522 164556 79524
rect 164325 79520 164556 79522
rect 164325 79464 164330 79520
rect 164386 79464 164556 79520
rect 164325 79462 164556 79464
rect 164325 79459 164391 79462
rect 164550 79460 164556 79462
rect 164620 79460 164626 79524
rect 167862 79460 167868 79524
rect 167932 79522 167938 79524
rect 168281 79522 168347 79525
rect 167932 79520 168347 79522
rect 167932 79464 168286 79520
rect 168342 79464 168347 79520
rect 167932 79462 168347 79464
rect 167932 79460 167938 79462
rect 168281 79459 168347 79462
rect 168833 79520 168899 79525
rect 169385 79524 169451 79525
rect 169334 79522 169340 79524
rect 168833 79464 168838 79520
rect 168894 79464 168899 79520
rect 168833 79459 168899 79464
rect 169294 79462 169340 79522
rect 169404 79520 169451 79524
rect 169446 79464 169451 79520
rect 169334 79460 169340 79462
rect 169404 79460 169451 79464
rect 169518 79460 169524 79524
rect 169588 79522 169594 79524
rect 169661 79522 169727 79525
rect 169588 79520 169727 79522
rect 169588 79464 169666 79520
rect 169722 79464 169727 79520
rect 169588 79462 169727 79464
rect 169588 79460 169594 79462
rect 169385 79459 169451 79460
rect 169661 79459 169727 79462
rect 170438 79460 170444 79524
rect 170508 79522 170514 79524
rect 171041 79522 171107 79525
rect 170508 79520 171107 79522
rect 170508 79464 171046 79520
rect 171102 79464 171107 79520
rect 170508 79462 171107 79464
rect 171320 79522 171380 79595
rect 173712 79525 173772 79870
rect 172605 79522 172671 79525
rect 171320 79520 172671 79522
rect 171320 79464 172610 79520
rect 172666 79464 172671 79520
rect 171320 79462 172671 79464
rect 170508 79460 170514 79462
rect 171041 79459 171107 79462
rect 172605 79459 172671 79462
rect 173709 79520 173775 79525
rect 173709 79464 173714 79520
rect 173770 79464 173775 79520
rect 173709 79459 173775 79464
rect 174310 79522 174370 79904
rect 174670 79868 174676 79932
rect 174740 79930 174746 79932
rect 175227 79930 175293 79933
rect 174740 79928 175293 79930
rect 174740 79872 175232 79928
rect 175288 79872 175293 79928
rect 174740 79870 175293 79872
rect 174740 79868 174746 79870
rect 175227 79867 175293 79870
rect 175503 79930 175569 79933
rect 176326 79930 176332 79932
rect 175503 79928 176332 79930
rect 175503 79872 175508 79928
rect 175564 79872 176332 79928
rect 175503 79870 176332 79872
rect 175503 79867 175569 79870
rect 176326 79868 176332 79870
rect 176396 79868 176402 79932
rect 176515 79906 176520 79962
rect 176576 79906 176581 79962
rect 176515 79901 176581 79906
rect 176791 79930 176857 79933
rect 177070 79930 177130 80006
rect 180241 80003 180307 80006
rect 176791 79928 177130 79930
rect 176791 79872 176796 79928
rect 176852 79872 177130 79928
rect 176791 79870 177130 79872
rect 177343 79930 177409 79933
rect 177803 79932 177869 79933
rect 178355 79932 178421 79933
rect 177343 79928 177682 79930
rect 177343 79872 177348 79928
rect 177404 79872 177682 79928
rect 177343 79870 177682 79872
rect 176791 79867 176857 79870
rect 177343 79867 177409 79870
rect 174951 79794 175017 79797
rect 175779 79794 175845 79797
rect 176142 79794 176148 79796
rect 174951 79792 175060 79794
rect 174951 79736 174956 79792
rect 175012 79736 175060 79792
rect 174951 79731 175060 79736
rect 175779 79792 176148 79794
rect 175779 79736 175784 79792
rect 175840 79736 176148 79792
rect 175779 79734 176148 79736
rect 175779 79731 175845 79734
rect 176142 79732 176148 79734
rect 176212 79732 176218 79796
rect 176745 79794 176811 79797
rect 176878 79794 176884 79796
rect 176745 79792 176884 79794
rect 176745 79736 176750 79792
rect 176806 79736 176884 79792
rect 176745 79734 176884 79736
rect 176745 79731 176811 79734
rect 176878 79732 176884 79734
rect 176948 79732 176954 79796
rect 175000 79660 175060 79731
rect 175181 79660 175247 79661
rect 175000 79598 175044 79660
rect 175038 79596 175044 79598
rect 175108 79596 175114 79660
rect 175181 79656 175228 79660
rect 175292 79658 175298 79660
rect 176469 79658 176535 79661
rect 177430 79658 177436 79660
rect 175181 79600 175186 79656
rect 175181 79596 175228 79600
rect 175292 79598 175338 79658
rect 176469 79656 177436 79658
rect 176469 79600 176474 79656
rect 176530 79600 177436 79656
rect 176469 79598 177436 79600
rect 175292 79596 175298 79598
rect 175181 79595 175247 79596
rect 176469 79595 176535 79598
rect 177430 79596 177436 79598
rect 177500 79596 177506 79660
rect 177062 79522 177068 79524
rect 174310 79462 177068 79522
rect 177062 79460 177068 79462
rect 177132 79460 177138 79524
rect 177622 79522 177682 79870
rect 177798 79868 177804 79932
rect 177868 79930 177874 79932
rect 178350 79930 178356 79932
rect 177868 79870 177960 79930
rect 178264 79870 178356 79930
rect 177868 79868 177874 79870
rect 178350 79868 178356 79870
rect 178420 79868 178426 79932
rect 177803 79867 177869 79868
rect 178355 79867 178421 79868
rect 177757 79794 177823 79797
rect 177757 79792 186330 79794
rect 177757 79736 177762 79792
rect 177818 79736 186330 79792
rect 177757 79734 186330 79736
rect 177757 79731 177823 79734
rect 177757 79658 177823 79661
rect 186270 79658 186330 79734
rect 266353 79658 266419 79661
rect 177757 79656 183570 79658
rect 177757 79600 177762 79656
rect 177818 79600 183570 79656
rect 177757 79598 183570 79600
rect 186270 79656 266419 79658
rect 186270 79600 266358 79656
rect 266414 79600 266419 79656
rect 186270 79598 266419 79600
rect 177757 79595 177823 79598
rect 179781 79522 179847 79525
rect 177622 79520 179847 79522
rect 177622 79464 179786 79520
rect 179842 79464 179847 79520
rect 177622 79462 179847 79464
rect 183510 79522 183570 79598
rect 266353 79595 266419 79598
rect 331213 79522 331279 79525
rect 183510 79520 331279 79522
rect 183510 79464 331218 79520
rect 331274 79464 331279 79520
rect 183510 79462 331279 79464
rect 179781 79459 179847 79462
rect 331213 79459 331279 79462
rect 6913 79386 6979 79389
rect 176285 79386 176351 79389
rect 176653 79388 176719 79389
rect 176653 79386 176700 79388
rect 6913 79384 176351 79386
rect 6913 79328 6918 79384
rect 6974 79328 176290 79384
rect 176346 79328 176351 79384
rect 6913 79326 176351 79328
rect 176608 79384 176700 79386
rect 176608 79328 176658 79384
rect 176608 79326 176700 79328
rect 6913 79323 6979 79326
rect 176285 79323 176351 79326
rect 176653 79324 176700 79326
rect 176764 79324 176770 79388
rect 177573 79386 177639 79389
rect 580257 79386 580323 79389
rect 177573 79384 580323 79386
rect 177573 79328 177578 79384
rect 177634 79328 580262 79384
rect 580318 79328 580323 79384
rect 177573 79326 580323 79328
rect 176653 79323 176719 79324
rect 177573 79323 177639 79326
rect 580257 79323 580323 79326
rect 3601 79250 3667 79253
rect 175273 79250 175339 79253
rect 178033 79250 178099 79253
rect 3601 79248 175339 79250
rect 3601 79192 3606 79248
rect 3662 79192 175278 79248
rect 175334 79192 175339 79248
rect 3601 79190 175339 79192
rect 3601 79187 3667 79190
rect 175273 79187 175339 79190
rect 175506 79248 178099 79250
rect 175506 79192 178038 79248
rect 178094 79192 178099 79248
rect 175506 79190 178099 79192
rect 3417 79114 3483 79117
rect 175506 79114 175566 79190
rect 178033 79187 178099 79190
rect 178217 79250 178283 79253
rect 178350 79250 178356 79252
rect 178217 79248 178356 79250
rect 178217 79192 178222 79248
rect 178278 79192 178356 79248
rect 178217 79190 178356 79192
rect 178217 79187 178283 79190
rect 178350 79188 178356 79190
rect 178420 79188 178426 79252
rect 3417 79112 175566 79114
rect 3417 79056 3422 79112
rect 3478 79056 175566 79112
rect 3417 79054 175566 79056
rect 175641 79114 175707 79117
rect 179137 79114 179203 79117
rect 175641 79112 179203 79114
rect 175641 79056 175646 79112
rect 175702 79056 179142 79112
rect 179198 79056 179203 79112
rect 175641 79054 179203 79056
rect 3417 79051 3483 79054
rect 175641 79051 175707 79054
rect 179137 79051 179203 79054
rect 130561 78978 130627 78981
rect 131246 78978 131252 78980
rect 130561 78976 131252 78978
rect 130561 78920 130566 78976
rect 130622 78920 131252 78976
rect 130561 78918 131252 78920
rect 130561 78915 130627 78918
rect 131246 78916 131252 78918
rect 131316 78916 131322 78980
rect 141785 78978 141851 78981
rect 141918 78978 141924 78980
rect 141785 78976 141924 78978
rect 141785 78920 141790 78976
rect 141846 78920 141924 78976
rect 141785 78918 141924 78920
rect 141785 78915 141851 78918
rect 141918 78916 141924 78918
rect 141988 78916 141994 78980
rect 149605 78978 149671 78981
rect 158253 78978 158319 78981
rect 149605 78976 158319 78978
rect 149605 78920 149610 78976
rect 149666 78920 158258 78976
rect 158314 78920 158319 78976
rect 149605 78918 158319 78920
rect 149605 78915 149671 78918
rect 158253 78915 158319 78918
rect 163630 78916 163636 78980
rect 163700 78978 163706 78980
rect 164049 78978 164115 78981
rect 163700 78976 164115 78978
rect 163700 78920 164054 78976
rect 164110 78920 164115 78976
rect 163700 78918 164115 78920
rect 163700 78916 163706 78918
rect 164049 78915 164115 78918
rect 165613 78978 165679 78981
rect 173249 78978 173315 78981
rect 173617 78980 173683 78981
rect 173566 78978 173572 78980
rect 165613 78976 173315 78978
rect 165613 78920 165618 78976
rect 165674 78920 173254 78976
rect 173310 78920 173315 78976
rect 165613 78918 173315 78920
rect 173526 78918 173572 78978
rect 173636 78976 173683 78980
rect 173678 78920 173683 78976
rect 165613 78915 165679 78918
rect 173249 78915 173315 78918
rect 173566 78916 173572 78918
rect 173636 78916 173683 78920
rect 173617 78915 173683 78916
rect 175089 78978 175155 78981
rect 175222 78978 175228 78980
rect 175089 78976 175228 78978
rect 175089 78920 175094 78976
rect 175150 78920 175228 78976
rect 175089 78918 175228 78920
rect 175089 78915 175155 78918
rect 175222 78916 175228 78918
rect 175292 78916 175298 78980
rect 175549 78978 175615 78981
rect 175774 78978 175780 78980
rect 175549 78976 175780 78978
rect 175549 78920 175554 78976
rect 175610 78920 175780 78976
rect 175549 78918 175780 78920
rect 175549 78915 175615 78918
rect 175774 78916 175780 78918
rect 175844 78916 175850 78980
rect 176142 78916 176148 78980
rect 176212 78978 176218 78980
rect 176510 78978 176516 78980
rect 176212 78918 176516 78978
rect 176212 78916 176218 78918
rect 176510 78916 176516 78918
rect 176580 78916 176586 78980
rect 177665 78978 177731 78981
rect 397453 78978 397519 78981
rect 177665 78976 397519 78978
rect 177665 78920 177670 78976
rect 177726 78920 397458 78976
rect 397514 78920 397519 78976
rect 177665 78918 397519 78920
rect 177665 78915 177731 78918
rect 397453 78915 397519 78918
rect 119337 78842 119403 78845
rect 177205 78842 177271 78845
rect 119337 78840 177271 78842
rect 119337 78784 119342 78840
rect 119398 78784 177210 78840
rect 177266 78784 177271 78840
rect 119337 78782 177271 78784
rect 119337 78779 119403 78782
rect 177205 78779 177271 78782
rect 177481 78842 177547 78845
rect 462313 78842 462379 78845
rect 177481 78840 462379 78842
rect 177481 78784 177486 78840
rect 177542 78784 462318 78840
rect 462374 78784 462379 78840
rect 177481 78782 462379 78784
rect 177481 78779 177547 78782
rect 462313 78779 462379 78782
rect 132493 78706 132559 78709
rect 133454 78706 133460 78708
rect 132493 78704 133460 78706
rect 132493 78648 132498 78704
rect 132554 78648 133460 78704
rect 132493 78646 133460 78648
rect 132493 78643 132559 78646
rect 133454 78644 133460 78646
rect 133524 78644 133530 78708
rect 137921 78706 137987 78709
rect 138238 78706 138244 78708
rect 137921 78704 138244 78706
rect 137921 78648 137926 78704
rect 137982 78648 138244 78704
rect 137921 78646 138244 78648
rect 137921 78643 137987 78646
rect 138238 78644 138244 78646
rect 138308 78644 138314 78708
rect 150014 78644 150020 78708
rect 150084 78706 150090 78708
rect 150157 78706 150223 78709
rect 150084 78704 150223 78706
rect 150084 78648 150162 78704
rect 150218 78648 150223 78704
rect 150084 78646 150223 78648
rect 150084 78644 150090 78646
rect 150157 78643 150223 78646
rect 157926 78644 157932 78708
rect 157996 78706 158002 78708
rect 158345 78706 158411 78709
rect 157996 78704 158411 78706
rect 157996 78648 158350 78704
rect 158406 78648 158411 78704
rect 157996 78646 158411 78648
rect 157996 78644 158002 78646
rect 158345 78643 158411 78646
rect 163446 78644 163452 78708
rect 163516 78706 163522 78708
rect 163957 78706 164023 78709
rect 163516 78704 164023 78706
rect 163516 78648 163962 78704
rect 164018 78648 164023 78704
rect 163516 78646 164023 78648
rect 163516 78644 163522 78646
rect 163957 78643 164023 78646
rect 168557 78706 168623 78709
rect 168966 78706 168972 78708
rect 168557 78704 168972 78706
rect 168557 78648 168562 78704
rect 168618 78648 168972 78704
rect 168557 78646 168972 78648
rect 168557 78643 168623 78646
rect 168966 78644 168972 78646
rect 169036 78644 169042 78708
rect 170673 78706 170739 78709
rect 170990 78706 170996 78708
rect 170673 78704 170996 78706
rect 170673 78648 170678 78704
rect 170734 78648 170996 78704
rect 170673 78646 170996 78648
rect 170673 78643 170739 78646
rect 170990 78644 170996 78646
rect 171060 78644 171066 78708
rect 172053 78706 172119 78709
rect 171550 78704 172119 78706
rect 171550 78648 172058 78704
rect 172114 78648 172119 78704
rect 171550 78646 172119 78648
rect 119429 78570 119495 78573
rect 171550 78570 171610 78646
rect 172053 78643 172119 78646
rect 172697 78706 172763 78709
rect 173801 78708 173867 78709
rect 173382 78706 173388 78708
rect 172697 78704 173388 78706
rect 172697 78648 172702 78704
rect 172758 78648 173388 78704
rect 172697 78646 173388 78648
rect 172697 78643 172763 78646
rect 173382 78644 173388 78646
rect 173452 78644 173458 78708
rect 173750 78706 173756 78708
rect 173710 78646 173756 78706
rect 173820 78704 173867 78708
rect 173862 78648 173867 78704
rect 173750 78644 173756 78646
rect 173820 78644 173867 78648
rect 174854 78644 174860 78708
rect 174924 78706 174930 78708
rect 174997 78706 175063 78709
rect 174924 78704 175063 78706
rect 174924 78648 175002 78704
rect 175058 78648 175063 78704
rect 174924 78646 175063 78648
rect 174924 78644 174930 78646
rect 173801 78643 173867 78644
rect 174997 78643 175063 78646
rect 175457 78706 175523 78709
rect 176142 78706 176148 78708
rect 175457 78704 176148 78706
rect 175457 78648 175462 78704
rect 175518 78648 176148 78704
rect 175457 78646 176148 78648
rect 175457 78643 175523 78646
rect 176142 78644 176148 78646
rect 176212 78644 176218 78708
rect 180241 78706 180307 78709
rect 580533 78706 580599 78709
rect 180241 78704 580599 78706
rect 180241 78648 180246 78704
rect 180302 78648 580538 78704
rect 580594 78648 580599 78704
rect 180241 78646 580599 78648
rect 180241 78643 180307 78646
rect 580533 78643 580599 78646
rect 119429 78568 171610 78570
rect 119429 78512 119434 78568
rect 119490 78512 171610 78568
rect 119429 78510 171610 78512
rect 171734 78510 177130 78570
rect 119429 78507 119495 78510
rect 133045 78434 133111 78437
rect 133638 78434 133644 78436
rect 133045 78432 133644 78434
rect 133045 78376 133050 78432
rect 133106 78376 133644 78432
rect 133045 78374 133644 78376
rect 133045 78371 133111 78374
rect 133638 78372 133644 78374
rect 133708 78372 133714 78436
rect 136817 78434 136883 78437
rect 137870 78434 137876 78436
rect 136817 78432 137876 78434
rect 136817 78376 136822 78432
rect 136878 78376 137876 78432
rect 136817 78374 137876 78376
rect 136817 78371 136883 78374
rect 137870 78372 137876 78374
rect 137940 78372 137946 78436
rect 144494 78372 144500 78436
rect 144564 78434 144570 78436
rect 148317 78434 148383 78437
rect 144564 78432 148383 78434
rect 144564 78376 148322 78432
rect 148378 78376 148383 78432
rect 144564 78374 148383 78376
rect 144564 78372 144570 78374
rect 148317 78371 148383 78374
rect 151486 78372 151492 78436
rect 151556 78434 151562 78436
rect 155769 78434 155835 78437
rect 151556 78432 155835 78434
rect 151556 78376 155774 78432
rect 155830 78376 155835 78432
rect 151556 78374 155835 78376
rect 151556 78372 151562 78374
rect 155769 78371 155835 78374
rect 163221 78434 163287 78437
rect 171734 78434 171794 78510
rect 176929 78434 176995 78437
rect 163221 78432 171794 78434
rect 163221 78376 163226 78432
rect 163282 78376 171794 78432
rect 163221 78374 171794 78376
rect 171918 78432 176995 78434
rect 171918 78376 176934 78432
rect 176990 78376 176995 78432
rect 171918 78374 176995 78376
rect 177070 78434 177130 78510
rect 177573 78434 177639 78437
rect 177070 78432 177639 78434
rect 177070 78376 177578 78432
rect 177634 78376 177639 78432
rect 177070 78374 177639 78376
rect 163221 78371 163287 78374
rect 162025 78298 162091 78301
rect 162526 78298 162532 78300
rect 162025 78296 162532 78298
rect 162025 78240 162030 78296
rect 162086 78240 162532 78296
rect 162025 78238 162532 78240
rect 162025 78235 162091 78238
rect 162526 78236 162532 78238
rect 162596 78236 162602 78300
rect 163998 78236 164004 78300
rect 164068 78298 164074 78300
rect 170949 78298 171015 78301
rect 164068 78296 171015 78298
rect 164068 78240 170954 78296
rect 171010 78240 171015 78296
rect 164068 78238 171015 78240
rect 164068 78236 164074 78238
rect 170949 78235 171015 78238
rect 171593 78298 171659 78301
rect 171726 78298 171732 78300
rect 171593 78296 171732 78298
rect 171593 78240 171598 78296
rect 171654 78240 171732 78296
rect 171593 78238 171732 78240
rect 171593 78235 171659 78238
rect 171726 78236 171732 78238
rect 171796 78236 171802 78300
rect 133965 78162 134031 78165
rect 134558 78162 134564 78164
rect 133965 78160 134564 78162
rect 133965 78104 133970 78160
rect 134026 78104 134564 78160
rect 133965 78102 134564 78104
rect 133965 78099 134031 78102
rect 134558 78100 134564 78102
rect 134628 78100 134634 78164
rect 143758 78100 143764 78164
rect 143828 78162 143834 78164
rect 143901 78162 143967 78165
rect 143828 78160 143967 78162
rect 143828 78104 143906 78160
rect 143962 78104 143967 78160
rect 143828 78102 143967 78104
rect 143828 78100 143834 78102
rect 143901 78099 143967 78102
rect 144678 78100 144684 78164
rect 144748 78162 144754 78164
rect 144821 78162 144887 78165
rect 144748 78160 144887 78162
rect 144748 78104 144826 78160
rect 144882 78104 144887 78160
rect 144748 78102 144887 78104
rect 144748 78100 144754 78102
rect 144821 78099 144887 78102
rect 154849 78162 154915 78165
rect 155350 78162 155356 78164
rect 154849 78160 155356 78162
rect 154849 78104 154854 78160
rect 154910 78104 155356 78160
rect 154849 78102 155356 78104
rect 154849 78099 154915 78102
rect 155350 78100 155356 78102
rect 155420 78100 155426 78164
rect 165429 78162 165495 78165
rect 171918 78162 171978 78374
rect 176929 78371 176995 78374
rect 177573 78371 177639 78374
rect 172053 78298 172119 78301
rect 179689 78298 179755 78301
rect 172053 78296 179755 78298
rect 172053 78240 172058 78296
rect 172114 78240 179694 78296
rect 179750 78240 179755 78296
rect 172053 78238 179755 78240
rect 172053 78235 172119 78238
rect 179689 78235 179755 78238
rect 165429 78160 171978 78162
rect 165429 78104 165434 78160
rect 165490 78104 171978 78160
rect 165429 78102 171978 78104
rect 172237 78164 172303 78165
rect 172237 78160 172284 78164
rect 172348 78162 172354 78164
rect 172237 78104 172242 78160
rect 165429 78099 165495 78102
rect 172237 78100 172284 78104
rect 172348 78102 172394 78162
rect 172348 78100 172354 78102
rect 172646 78100 172652 78164
rect 172716 78162 172722 78164
rect 173065 78162 173131 78165
rect 172716 78160 173131 78162
rect 172716 78104 173070 78160
rect 173126 78104 173131 78160
rect 172716 78102 173131 78104
rect 172716 78100 172722 78102
rect 172237 78099 172303 78100
rect 173065 78099 173131 78102
rect 173198 78100 173204 78164
rect 173268 78162 173274 78164
rect 175825 78162 175891 78165
rect 173268 78160 175891 78162
rect 173268 78104 175830 78160
rect 175886 78104 175891 78160
rect 173268 78102 175891 78104
rect 173268 78100 173274 78102
rect 175825 78099 175891 78102
rect 176929 78162 176995 78165
rect 180241 78162 180307 78165
rect 176929 78160 180307 78162
rect 176929 78104 176934 78160
rect 176990 78104 180246 78160
rect 180302 78104 180307 78160
rect 176929 78102 180307 78104
rect 176929 78099 176995 78102
rect 180241 78099 180307 78102
rect 131062 77964 131068 78028
rect 131132 78026 131138 78028
rect 131205 78026 131271 78029
rect 131132 78024 131271 78026
rect 131132 77968 131210 78024
rect 131266 77968 131271 78024
rect 131132 77966 131271 77968
rect 131132 77964 131138 77966
rect 131205 77963 131271 77966
rect 134190 77964 134196 78028
rect 134260 78026 134266 78028
rect 134425 78026 134491 78029
rect 134260 78024 134491 78026
rect 134260 77968 134430 78024
rect 134486 77968 134491 78024
rect 134260 77966 134491 77968
rect 134260 77964 134266 77966
rect 134425 77963 134491 77966
rect 135294 77964 135300 78028
rect 135364 78026 135370 78028
rect 135437 78026 135503 78029
rect 135364 78024 135503 78026
rect 135364 77968 135442 78024
rect 135498 77968 135503 78024
rect 135364 77966 135503 77968
rect 135364 77964 135370 77966
rect 135437 77963 135503 77966
rect 135621 78028 135687 78029
rect 135621 78024 135668 78028
rect 135732 78026 135738 78028
rect 135621 77968 135626 78024
rect 135621 77964 135668 77968
rect 135732 77966 135778 78026
rect 135732 77964 135738 77966
rect 139158 77964 139164 78028
rect 139228 78026 139234 78028
rect 146937 78026 147003 78029
rect 139228 78024 147003 78026
rect 139228 77968 146942 78024
rect 146998 77968 147003 78024
rect 139228 77966 147003 77968
rect 139228 77964 139234 77966
rect 135621 77963 135687 77964
rect 146937 77963 147003 77966
rect 164918 77964 164924 78028
rect 164988 78026 164994 78028
rect 165245 78026 165311 78029
rect 165521 78028 165587 78029
rect 165470 78026 165476 78028
rect 164988 78024 165311 78026
rect 164988 77968 165250 78024
rect 165306 77968 165311 78024
rect 164988 77966 165311 77968
rect 165430 77966 165476 78026
rect 165540 78024 165587 78028
rect 165582 77968 165587 78024
rect 164988 77964 164994 77966
rect 165245 77963 165311 77966
rect 165470 77964 165476 77966
rect 165540 77964 165587 77968
rect 165521 77963 165587 77964
rect 166441 78026 166507 78029
rect 260097 78026 260163 78029
rect 166441 78024 260163 78026
rect 166441 77968 166446 78024
rect 166502 77968 260102 78024
rect 260158 77968 260163 78024
rect 166441 77966 260163 77968
rect 166441 77963 166507 77966
rect 260097 77963 260163 77966
rect 13077 77890 13143 77893
rect 131297 77890 131363 77893
rect 161565 77890 161631 77893
rect 13077 77888 131363 77890
rect 13077 77832 13082 77888
rect 13138 77832 131302 77888
rect 131358 77832 131363 77888
rect 13077 77830 131363 77832
rect 13077 77827 13143 77830
rect 131297 77827 131363 77830
rect 131622 77888 161631 77890
rect 131622 77832 161570 77888
rect 161626 77832 161631 77888
rect 131622 77830 161631 77832
rect 129549 77754 129615 77757
rect 131622 77754 131682 77830
rect 161565 77827 161631 77830
rect 164550 77828 164556 77892
rect 164620 77890 164626 77892
rect 168005 77890 168071 77893
rect 164620 77888 168071 77890
rect 164620 77832 168010 77888
rect 168066 77832 168071 77888
rect 164620 77830 168071 77832
rect 164620 77828 164626 77830
rect 168005 77827 168071 77830
rect 170949 77890 171015 77893
rect 175273 77890 175339 77893
rect 480253 77890 480319 77893
rect 170949 77888 175339 77890
rect 170949 77832 170954 77888
rect 171010 77832 175278 77888
rect 175334 77832 175339 77888
rect 170949 77830 175339 77832
rect 170949 77827 171015 77830
rect 175273 77827 175339 77830
rect 176610 77888 480319 77890
rect 176610 77832 480258 77888
rect 480314 77832 480319 77888
rect 176610 77830 480319 77832
rect 129549 77752 131682 77754
rect 129549 77696 129554 77752
rect 129610 77696 131682 77752
rect 129549 77694 131682 77696
rect 169937 77754 170003 77757
rect 170254 77754 170260 77756
rect 169937 77752 170260 77754
rect 169937 77696 169942 77752
rect 169998 77696 170260 77752
rect 169937 77694 170260 77696
rect 129549 77691 129615 77694
rect 169937 77691 170003 77694
rect 170254 77692 170260 77694
rect 170324 77692 170330 77756
rect 156638 77556 156644 77620
rect 156708 77618 156714 77620
rect 157241 77618 157307 77621
rect 156708 77616 157307 77618
rect 156708 77560 157246 77616
rect 157302 77560 157307 77616
rect 156708 77558 157307 77560
rect 156708 77556 156714 77558
rect 157241 77555 157307 77558
rect 161974 77556 161980 77620
rect 162044 77618 162050 77620
rect 165613 77618 165679 77621
rect 162044 77616 165679 77618
rect 162044 77560 165618 77616
rect 165674 77560 165679 77616
rect 162044 77558 165679 77560
rect 162044 77556 162050 77558
rect 165613 77555 165679 77558
rect 166390 77556 166396 77620
rect 166460 77618 166466 77620
rect 166993 77618 167059 77621
rect 166460 77616 167059 77618
rect 166460 77560 166998 77616
rect 167054 77560 167059 77616
rect 166460 77558 167059 77560
rect 166460 77556 166466 77558
rect 166993 77555 167059 77558
rect 170765 77618 170831 77621
rect 176610 77618 176670 77830
rect 480253 77827 480319 77830
rect 170765 77616 176670 77618
rect 170765 77560 170770 77616
rect 170826 77560 176670 77616
rect 170765 77558 176670 77560
rect 170765 77555 170831 77558
rect 145414 77420 145420 77484
rect 145484 77482 145490 77484
rect 146201 77482 146267 77485
rect 145484 77480 146267 77482
rect 145484 77424 146206 77480
rect 146262 77424 146267 77480
rect 145484 77422 146267 77424
rect 145484 77420 145490 77422
rect 146201 77419 146267 77422
rect 147070 77420 147076 77484
rect 147140 77482 147146 77484
rect 147305 77482 147371 77485
rect 147140 77480 147371 77482
rect 147140 77424 147310 77480
rect 147366 77424 147371 77480
rect 147140 77422 147371 77424
rect 147140 77420 147146 77422
rect 147305 77419 147371 77422
rect 152406 77420 152412 77484
rect 152476 77482 152482 77484
rect 153285 77482 153351 77485
rect 152476 77480 153351 77482
rect 152476 77424 153290 77480
rect 153346 77424 153351 77480
rect 152476 77422 153351 77424
rect 152476 77420 152482 77422
rect 153285 77419 153351 77422
rect 154246 77420 154252 77484
rect 154316 77482 154322 77484
rect 154481 77482 154547 77485
rect 154316 77480 154547 77482
rect 154316 77424 154486 77480
rect 154542 77424 154547 77480
rect 154316 77422 154547 77424
rect 154316 77420 154322 77422
rect 154481 77419 154547 77422
rect 157006 77420 157012 77484
rect 157076 77482 157082 77484
rect 157149 77482 157215 77485
rect 157076 77480 157215 77482
rect 157076 77424 157154 77480
rect 157210 77424 157215 77480
rect 157076 77422 157215 77424
rect 157076 77420 157082 77422
rect 157149 77419 157215 77422
rect 166717 77484 166783 77485
rect 172145 77484 172211 77485
rect 166717 77480 166764 77484
rect 166828 77482 166834 77484
rect 172094 77482 172100 77484
rect 166717 77424 166722 77480
rect 166717 77420 166764 77424
rect 166828 77422 166874 77482
rect 172054 77422 172100 77482
rect 172164 77480 172211 77484
rect 172206 77424 172211 77480
rect 166828 77420 166834 77422
rect 172094 77420 172100 77422
rect 172164 77420 172211 77424
rect 166717 77419 166783 77420
rect 172145 77419 172211 77420
rect 145230 77284 145236 77348
rect 145300 77346 145306 77348
rect 145465 77346 145531 77349
rect 145300 77344 145531 77346
rect 145300 77288 145470 77344
rect 145526 77288 145531 77344
rect 145300 77286 145531 77288
rect 145300 77284 145306 77286
rect 145465 77283 145531 77286
rect 147254 77284 147260 77348
rect 147324 77346 147330 77348
rect 147397 77346 147463 77349
rect 147324 77344 147463 77346
rect 147324 77288 147402 77344
rect 147458 77288 147463 77344
rect 147324 77286 147463 77288
rect 147324 77284 147330 77286
rect 147397 77283 147463 77286
rect 152774 77284 152780 77348
rect 152844 77346 152850 77348
rect 153009 77346 153075 77349
rect 152844 77344 153075 77346
rect 152844 77288 153014 77344
rect 153070 77288 153075 77344
rect 152844 77286 153075 77288
rect 152844 77284 152850 77286
rect 153009 77283 153075 77286
rect 153469 77346 153535 77349
rect 153694 77346 153700 77348
rect 153469 77344 153700 77346
rect 153469 77288 153474 77344
rect 153530 77288 153700 77344
rect 153469 77286 153700 77288
rect 153469 77283 153535 77286
rect 153694 77284 153700 77286
rect 153764 77284 153770 77348
rect 154062 77284 154068 77348
rect 154132 77346 154138 77348
rect 154297 77346 154363 77349
rect 154132 77344 154363 77346
rect 154132 77288 154302 77344
rect 154358 77288 154363 77344
rect 154132 77286 154363 77288
rect 154132 77284 154138 77286
rect 154297 77283 154363 77286
rect 154614 77284 154620 77348
rect 154684 77346 154690 77348
rect 155217 77346 155283 77349
rect 156321 77348 156387 77349
rect 154684 77344 155283 77346
rect 154684 77288 155222 77344
rect 155278 77288 155283 77344
rect 154684 77286 155283 77288
rect 154684 77284 154690 77286
rect 155217 77283 155283 77286
rect 156270 77284 156276 77348
rect 156340 77346 156387 77348
rect 156340 77344 156432 77346
rect 156382 77288 156432 77344
rect 156340 77286 156432 77288
rect 156340 77284 156387 77286
rect 158478 77284 158484 77348
rect 158548 77346 158554 77348
rect 158621 77346 158687 77349
rect 158548 77344 158687 77346
rect 158548 77288 158626 77344
rect 158682 77288 158687 77344
rect 158548 77286 158687 77288
rect 158548 77284 158554 77286
rect 156321 77283 156387 77284
rect 158621 77283 158687 77286
rect 159030 77284 159036 77348
rect 159100 77346 159106 77348
rect 160001 77346 160067 77349
rect 159100 77344 160067 77346
rect 159100 77288 160006 77344
rect 160062 77288 160067 77344
rect 159100 77286 160067 77288
rect 159100 77284 159106 77286
rect 160001 77283 160067 77286
rect 166206 77284 166212 77348
rect 166276 77346 166282 77348
rect 166625 77346 166691 77349
rect 166276 77344 166691 77346
rect 166276 77288 166630 77344
rect 166686 77288 166691 77344
rect 166276 77286 166691 77288
rect 166276 77284 166282 77286
rect 166625 77283 166691 77286
rect 167310 77284 167316 77348
rect 167380 77346 167386 77348
rect 168097 77346 168163 77349
rect 167380 77344 168163 77346
rect 167380 77288 168102 77344
rect 168158 77288 168163 77344
rect 167380 77286 168163 77288
rect 167380 77284 167386 77286
rect 168097 77283 168163 77286
rect 128997 77210 129063 77213
rect 134149 77210 134215 77213
rect 128997 77208 134215 77210
rect 128997 77152 129002 77208
rect 129058 77152 134154 77208
rect 134210 77152 134215 77208
rect 128997 77150 134215 77152
rect 128997 77147 129063 77150
rect 134149 77147 134215 77150
rect 148685 77210 148751 77213
rect 233233 77210 233299 77213
rect 148685 77208 233299 77210
rect 148685 77152 148690 77208
rect 148746 77152 233238 77208
rect 233294 77152 233299 77208
rect 148685 77150 233299 77152
rect 148685 77147 148751 77150
rect 233233 77147 233299 77150
rect 150341 77074 150407 77077
rect 253933 77074 253999 77077
rect 150341 77072 253999 77074
rect 150341 77016 150346 77072
rect 150402 77016 253938 77072
rect 253994 77016 253999 77072
rect 150341 77014 253999 77016
rect 150341 77011 150407 77014
rect 253933 77011 253999 77014
rect 115933 76938 115999 76941
rect 139485 76938 139551 76941
rect 115933 76936 139551 76938
rect 115933 76880 115938 76936
rect 115994 76880 139490 76936
rect 139546 76880 139551 76936
rect 115933 76878 139551 76880
rect 115933 76875 115999 76878
rect 139485 76875 139551 76878
rect 153101 76938 153167 76941
rect 289813 76938 289879 76941
rect 153101 76936 289879 76938
rect 153101 76880 153106 76936
rect 153162 76880 289818 76936
rect 289874 76880 289879 76936
rect 153101 76878 289879 76880
rect 153101 76875 153167 76878
rect 289813 76875 289879 76878
rect 97993 76802 98059 76805
rect 138054 76802 138060 76804
rect 97993 76800 138060 76802
rect 97993 76744 97998 76800
rect 98054 76744 138060 76800
rect 97993 76742 138060 76744
rect 97993 76739 98059 76742
rect 138054 76740 138060 76742
rect 138124 76740 138130 76804
rect 143022 76740 143028 76804
rect 143092 76802 143098 76804
rect 143165 76802 143231 76805
rect 143092 76800 143231 76802
rect 143092 76744 143170 76800
rect 143226 76744 143231 76800
rect 143092 76742 143231 76744
rect 143092 76740 143098 76742
rect 143165 76739 143231 76742
rect 154205 76802 154271 76805
rect 303613 76802 303679 76805
rect 154205 76800 303679 76802
rect 154205 76744 154210 76800
rect 154266 76744 303618 76800
rect 303674 76744 303679 76800
rect 154205 76742 303679 76744
rect 154205 76739 154271 76742
rect 303613 76739 303679 76742
rect 80053 76666 80119 76669
rect 136633 76666 136699 76669
rect 80053 76664 136699 76666
rect 80053 76608 80058 76664
rect 80114 76608 136638 76664
rect 136694 76608 136699 76664
rect 80053 76606 136699 76608
rect 80053 76603 80119 76606
rect 136633 76603 136699 76606
rect 142838 76604 142844 76668
rect 142908 76666 142914 76668
rect 143441 76666 143507 76669
rect 142908 76664 143507 76666
rect 142908 76608 143446 76664
rect 143502 76608 143507 76664
rect 142908 76606 143507 76608
rect 142908 76604 142914 76606
rect 143441 76603 143507 76606
rect 144310 76604 144316 76668
rect 144380 76666 144386 76668
rect 144729 76666 144795 76669
rect 144380 76664 144795 76666
rect 144380 76608 144734 76664
rect 144790 76608 144795 76664
rect 144380 76606 144795 76608
rect 144380 76604 144386 76606
rect 144729 76603 144795 76606
rect 147990 76604 147996 76668
rect 148060 76666 148066 76668
rect 148409 76666 148475 76669
rect 148060 76664 148475 76666
rect 148060 76608 148414 76664
rect 148470 76608 148475 76664
rect 148060 76606 148475 76608
rect 148060 76604 148066 76606
rect 148409 76603 148475 76606
rect 148542 76604 148548 76668
rect 148612 76666 148618 76668
rect 148961 76666 149027 76669
rect 148612 76664 149027 76666
rect 148612 76608 148966 76664
rect 149022 76608 149027 76664
rect 148612 76606 149027 76608
rect 148612 76604 148618 76606
rect 148961 76603 149027 76606
rect 150617 76666 150683 76669
rect 151118 76666 151124 76668
rect 150617 76664 151124 76666
rect 150617 76608 150622 76664
rect 150678 76608 151124 76664
rect 150617 76606 151124 76608
rect 150617 76603 150683 76606
rect 151118 76604 151124 76606
rect 151188 76604 151194 76668
rect 151486 76604 151492 76668
rect 151556 76666 151562 76668
rect 151721 76666 151787 76669
rect 151556 76664 151787 76666
rect 151556 76608 151726 76664
rect 151782 76608 151787 76664
rect 151556 76606 151787 76608
rect 151556 76604 151562 76606
rect 151721 76603 151787 76606
rect 153285 76666 153351 76669
rect 154430 76666 154436 76668
rect 153285 76664 154436 76666
rect 153285 76608 153290 76664
rect 153346 76608 154436 76664
rect 153285 76606 154436 76608
rect 153285 76603 153351 76606
rect 154430 76604 154436 76606
rect 154500 76604 154506 76668
rect 155861 76666 155927 76669
rect 324313 76666 324379 76669
rect 155861 76664 324379 76666
rect 155861 76608 155866 76664
rect 155922 76608 324318 76664
rect 324374 76608 324379 76664
rect 155861 76606 324379 76608
rect 155861 76603 155927 76606
rect 324313 76603 324379 76606
rect 11053 76530 11119 76533
rect 131430 76530 131436 76532
rect 11053 76528 131436 76530
rect 11053 76472 11058 76528
rect 11114 76472 131436 76528
rect 11053 76470 131436 76472
rect 11053 76467 11119 76470
rect 131430 76468 131436 76470
rect 131500 76468 131506 76532
rect 140998 76468 141004 76532
rect 141068 76530 141074 76532
rect 142981 76530 143047 76533
rect 141068 76528 143047 76530
rect 141068 76472 142986 76528
rect 143042 76472 143047 76528
rect 141068 76470 143047 76472
rect 141068 76468 141074 76470
rect 142981 76467 143047 76470
rect 160686 76468 160692 76532
rect 160756 76530 160762 76532
rect 160829 76530 160895 76533
rect 160756 76528 160895 76530
rect 160756 76472 160834 76528
rect 160890 76472 160895 76528
rect 160756 76470 160895 76472
rect 160756 76468 160762 76470
rect 160829 76467 160895 76470
rect 161381 76530 161447 76533
rect 396073 76530 396139 76533
rect 161381 76528 396139 76530
rect 161381 76472 161386 76528
rect 161442 76472 396078 76528
rect 396134 76472 396139 76528
rect 161381 76470 396139 76472
rect 161381 76467 161447 76470
rect 396073 76467 396139 76470
rect 147581 76394 147647 76397
rect 180057 76394 180123 76397
rect 147581 76392 180123 76394
rect 147581 76336 147586 76392
rect 147642 76336 180062 76392
rect 180118 76336 180123 76392
rect 147581 76334 180123 76336
rect 147581 76331 147647 76334
rect 180057 76331 180123 76334
rect 162158 76196 162164 76260
rect 162228 76258 162234 76260
rect 162669 76258 162735 76261
rect 164693 76260 164759 76261
rect 164693 76258 164740 76260
rect 162228 76256 162735 76258
rect 162228 76200 162674 76256
rect 162730 76200 162735 76256
rect 162228 76198 162735 76200
rect 164648 76256 164740 76258
rect 164648 76200 164698 76256
rect 164648 76198 164740 76200
rect 162228 76196 162234 76198
rect 162669 76195 162735 76198
rect 164693 76196 164740 76198
rect 164804 76196 164810 76260
rect 164693 76195 164759 76196
rect 162485 76122 162551 76125
rect 162710 76122 162716 76124
rect 162485 76120 162716 76122
rect 162485 76064 162490 76120
rect 162546 76064 162716 76120
rect 162485 76062 162716 76064
rect 162485 76059 162551 76062
rect 162710 76060 162716 76062
rect 162780 76060 162786 76124
rect 166758 75652 166764 75716
rect 166828 75714 166834 75716
rect 176101 75714 176167 75717
rect 166828 75712 176167 75714
rect 166828 75656 176106 75712
rect 176162 75656 176167 75712
rect 166828 75654 176167 75656
rect 166828 75652 166834 75654
rect 176101 75651 176167 75654
rect 144637 75578 144703 75581
rect 180793 75578 180859 75581
rect 144637 75576 180859 75578
rect 144637 75520 144642 75576
rect 144698 75520 180798 75576
rect 180854 75520 180859 75576
rect 144637 75518 180859 75520
rect 144637 75515 144703 75518
rect 180793 75515 180859 75518
rect 60733 75442 60799 75445
rect 135345 75442 135411 75445
rect 60733 75440 135411 75442
rect 60733 75384 60738 75440
rect 60794 75384 135350 75440
rect 135406 75384 135411 75440
rect 60733 75382 135411 75384
rect 60733 75379 60799 75382
rect 135345 75379 135411 75382
rect 148174 75380 148180 75444
rect 148244 75442 148250 75444
rect 148317 75442 148383 75445
rect 148244 75440 148383 75442
rect 148244 75384 148322 75440
rect 148378 75384 148383 75440
rect 148244 75382 148383 75384
rect 148244 75380 148250 75382
rect 148317 75379 148383 75382
rect 163262 75380 163268 75444
rect 163332 75442 163338 75444
rect 431953 75442 432019 75445
rect 163332 75440 432019 75442
rect 163332 75384 431958 75440
rect 432014 75384 432019 75440
rect 163332 75382 432019 75384
rect 163332 75380 163338 75382
rect 431953 75379 432019 75382
rect 44173 75306 44239 75309
rect 133822 75306 133828 75308
rect 44173 75304 133828 75306
rect 44173 75248 44178 75304
rect 44234 75248 133828 75304
rect 44173 75246 133828 75248
rect 44173 75243 44239 75246
rect 133822 75244 133828 75246
rect 133892 75244 133898 75308
rect 139526 75244 139532 75308
rect 139596 75306 139602 75308
rect 139853 75306 139919 75309
rect 139596 75304 139919 75306
rect 139596 75248 139858 75304
rect 139914 75248 139919 75304
rect 139596 75246 139919 75248
rect 139596 75244 139602 75246
rect 139853 75243 139919 75246
rect 140814 75244 140820 75308
rect 140884 75306 140890 75308
rect 142153 75306 142219 75309
rect 140884 75304 142219 75306
rect 140884 75248 142158 75304
rect 142214 75248 142219 75304
rect 140884 75246 142219 75248
rect 140884 75244 140890 75246
rect 142153 75243 142219 75246
rect 168189 75306 168255 75309
rect 481633 75306 481699 75309
rect 168189 75304 481699 75306
rect 168189 75248 168194 75304
rect 168250 75248 481638 75304
rect 481694 75248 481699 75304
rect 168189 75246 481699 75248
rect 168189 75243 168255 75246
rect 481633 75243 481699 75246
rect 6913 75170 6979 75173
rect 131062 75170 131068 75172
rect 6913 75168 131068 75170
rect 6913 75112 6918 75168
rect 6974 75112 131068 75168
rect 6913 75110 131068 75112
rect 6913 75107 6979 75110
rect 131062 75108 131068 75110
rect 131132 75108 131138 75172
rect 145598 75108 145604 75172
rect 145668 75170 145674 75172
rect 148869 75170 148935 75173
rect 145668 75168 148935 75170
rect 145668 75112 148874 75168
rect 148930 75112 148935 75168
rect 145668 75110 148935 75112
rect 145668 75108 145674 75110
rect 148869 75107 148935 75110
rect 172278 75108 172284 75172
rect 172348 75170 172354 75172
rect 535453 75170 535519 75173
rect 172348 75168 535519 75170
rect 172348 75112 535458 75168
rect 535514 75112 535519 75168
rect 172348 75110 535519 75112
rect 172348 75108 172354 75110
rect 535453 75107 535519 75110
rect 140957 75034 141023 75037
rect 142102 75034 142108 75036
rect 140957 75032 142108 75034
rect 140957 74976 140962 75032
rect 141018 74976 142108 75032
rect 140957 74974 142108 74976
rect 140957 74971 141023 74974
rect 142102 74972 142108 74974
rect 142172 74972 142178 75036
rect 175774 74428 175780 74492
rect 175844 74490 175850 74492
rect 176561 74490 176627 74493
rect 175844 74488 176627 74490
rect 175844 74432 176566 74488
rect 176622 74432 176627 74488
rect 175844 74430 176627 74432
rect 175844 74428 175850 74430
rect 176561 74427 176627 74430
rect 48313 73946 48379 73949
rect 134190 73946 134196 73948
rect 48313 73944 134196 73946
rect 48313 73888 48318 73944
rect 48374 73888 134196 73944
rect 48313 73886 134196 73888
rect 48313 73883 48379 73886
rect 134190 73884 134196 73886
rect 134260 73884 134266 73948
rect 149646 73884 149652 73948
rect 149716 73946 149722 73948
rect 251173 73946 251239 73949
rect 149716 73944 251239 73946
rect 149716 73888 251178 73944
rect 251234 73888 251239 73944
rect 149716 73886 251239 73888
rect 149716 73884 149722 73886
rect 251173 73883 251239 73886
rect 26233 73810 26299 73813
rect 133454 73810 133460 73812
rect 26233 73808 133460 73810
rect 26233 73752 26238 73808
rect 26294 73752 133460 73808
rect 26233 73750 133460 73752
rect 26233 73747 26299 73750
rect 133454 73748 133460 73750
rect 133524 73748 133530 73812
rect 152406 73748 152412 73812
rect 152476 73810 152482 73812
rect 287053 73810 287119 73813
rect 152476 73808 287119 73810
rect 152476 73752 287058 73808
rect 287114 73752 287119 73808
rect 152476 73750 287119 73752
rect 152476 73748 152482 73750
rect 287053 73747 287119 73750
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3417 71634 3483 71637
rect -960 71632 3483 71634
rect -960 71576 3422 71632
rect 3478 71576 3483 71632
rect -960 71574 3483 71576
rect -960 71484 480 71574
rect 3417 71571 3483 71574
rect 175222 71028 175228 71092
rect 175292 71090 175298 71092
rect 571333 71090 571399 71093
rect 175292 71088 571399 71090
rect 175292 71032 571338 71088
rect 571394 71032 571399 71088
rect 175292 71030 571399 71032
rect 175292 71028 175298 71030
rect 571333 71027 571399 71030
rect 144310 69532 144316 69596
rect 144380 69594 144386 69596
rect 182173 69594 182239 69597
rect 144380 69592 182239 69594
rect 144380 69536 182178 69592
rect 182234 69536 182239 69592
rect 144380 69534 182239 69536
rect 144380 69532 144386 69534
rect 182173 69531 182239 69534
rect 158846 68172 158852 68236
rect 158916 68234 158922 68236
rect 376753 68234 376819 68237
rect 158916 68232 376819 68234
rect 158916 68176 376758 68232
rect 376814 68176 376819 68232
rect 158916 68174 376819 68176
rect 158916 68172 158922 68174
rect 376753 68171 376819 68174
rect 176142 66812 176148 66876
rect 176212 66874 176218 66876
rect 575473 66874 575539 66877
rect 176212 66872 575539 66874
rect 176212 66816 575478 66872
rect 575534 66816 575539 66872
rect 176212 66814 575539 66816
rect 176212 66812 176218 66814
rect 575473 66811 575539 66814
rect 142838 66132 142844 66196
rect 142908 66194 142914 66196
rect 144177 66194 144243 66197
rect 142908 66192 144243 66194
rect 142908 66136 144182 66192
rect 144238 66136 144243 66192
rect 142908 66134 144243 66136
rect 142908 66132 142914 66134
rect 144177 66131 144243 66134
rect 144494 65452 144500 65516
rect 144564 65514 144570 65516
rect 159357 65514 159423 65517
rect 144564 65512 159423 65514
rect 144564 65456 159362 65512
rect 159418 65456 159423 65512
rect 144564 65454 159423 65456
rect 144564 65452 144570 65454
rect 159357 65451 159423 65454
rect 171910 65452 171916 65516
rect 171980 65514 171986 65516
rect 536833 65514 536899 65517
rect 171980 65512 536899 65514
rect 171980 65456 536838 65512
rect 536894 65456 536899 65512
rect 171980 65454 536899 65456
rect 171980 65452 171986 65454
rect 536833 65451 536899 65454
rect 167678 64228 167684 64292
rect 167748 64290 167754 64292
rect 483013 64290 483079 64293
rect 167748 64288 483079 64290
rect 167748 64232 483018 64288
rect 483074 64232 483079 64288
rect 167748 64230 483079 64232
rect 167748 64228 167754 64230
rect 483013 64227 483079 64230
rect 173566 64092 173572 64156
rect 173636 64154 173642 64156
rect 554773 64154 554839 64157
rect 173636 64152 554839 64154
rect 173636 64096 554778 64152
rect 554834 64096 554839 64152
rect 173636 64094 554839 64096
rect 173636 64092 173642 64094
rect 554773 64091 554839 64094
rect 169334 63548 169340 63612
rect 169404 63610 169410 63612
rect 170397 63610 170463 63613
rect 169404 63608 170463 63610
rect 169404 63552 170402 63608
rect 170458 63552 170463 63608
rect 169404 63550 170463 63552
rect 169404 63548 169410 63550
rect 170397 63547 170463 63550
rect 145230 62732 145236 62796
rect 145300 62794 145306 62796
rect 200113 62794 200179 62797
rect 145300 62792 200179 62794
rect 145300 62736 200118 62792
rect 200174 62736 200179 62792
rect 145300 62734 200179 62736
rect 145300 62732 145306 62734
rect 200113 62731 200179 62734
rect 170438 61372 170444 61436
rect 170508 61434 170514 61436
rect 518893 61434 518959 61437
rect 170508 61432 518959 61434
rect 170508 61376 518898 61432
rect 518954 61376 518959 61432
rect 170508 61374 518959 61376
rect 170508 61372 170514 61374
rect 518893 61371 518959 61374
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3509 58578 3575 58581
rect -960 58576 3575 58578
rect -960 58520 3514 58576
rect 3570 58520 3575 58576
rect -960 58518 3575 58520
rect -960 58428 480 58518
rect 3509 58515 3575 58518
rect 154062 55796 154068 55860
rect 154132 55858 154138 55860
rect 306373 55858 306439 55861
rect 154132 55856 306439 55858
rect 154132 55800 306378 55856
rect 306434 55800 306439 55856
rect 154132 55798 306439 55800
rect 154132 55796 154138 55798
rect 306373 55795 306439 55798
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 173750 46140 173756 46204
rect 173820 46202 173826 46204
rect 556153 46202 556219 46205
rect 173820 46200 556219 46202
rect 173820 46144 556158 46200
rect 556214 46144 556219 46200
rect 583520 46188 584960 46278
rect 173820 46142 556219 46144
rect 173820 46140 173826 46142
rect 556153 46139 556219 46142
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 140814 44236 140820 44300
rect 140884 44298 140890 44300
rect 142797 44298 142863 44301
rect 140884 44296 142863 44298
rect 140884 44240 142802 44296
rect 142858 44240 142863 44296
rect 140884 44238 142863 44240
rect 140884 44236 140890 44238
rect 142797 44235 142863 44238
rect 163446 36484 163452 36548
rect 163516 36546 163522 36548
rect 429193 36546 429259 36549
rect 163516 36544 429259 36546
rect 163516 36488 429198 36544
rect 429254 36488 429259 36544
rect 163516 36486 429259 36488
rect 163516 36484 163522 36486
rect 429193 36483 429259 36486
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3509 32466 3575 32469
rect -960 32464 3575 32466
rect -960 32408 3514 32464
rect 3570 32408 3575 32464
rect -960 32406 3575 32408
rect -960 32316 480 32406
rect 3509 32403 3575 32406
rect 151302 30908 151308 30972
rect 151372 30970 151378 30972
rect 271873 30970 271939 30973
rect 151372 30968 271939 30970
rect 151372 30912 271878 30968
rect 271934 30912 271939 30968
rect 151372 30910 271939 30912
rect 151372 30908 151378 30910
rect 271873 30907 271939 30910
rect 148542 29548 148548 29612
rect 148612 29610 148618 29612
rect 235993 29610 236059 29613
rect 148612 29608 236059 29610
rect 148612 29552 235998 29608
rect 236054 29552 236059 29608
rect 148612 29550 236059 29552
rect 148612 29548 148618 29550
rect 235993 29547 236059 29550
rect 147070 28188 147076 28252
rect 147140 28250 147146 28252
rect 215293 28250 215359 28253
rect 147140 28248 215359 28250
rect 147140 28192 215298 28248
rect 215354 28192 215359 28248
rect 147140 28190 215359 28192
rect 147140 28188 147146 28190
rect 215293 28187 215359 28190
rect 152774 26828 152780 26892
rect 152844 26890 152850 26892
rect 285673 26890 285739 26893
rect 152844 26888 285739 26890
rect 152844 26832 285678 26888
rect 285734 26832 285739 26888
rect 152844 26830 285739 26832
rect 152844 26828 152850 26830
rect 285673 26827 285739 26830
rect 144678 25604 144684 25668
rect 144748 25666 144754 25668
rect 183553 25666 183619 25669
rect 144748 25664 183619 25666
rect 144748 25608 183558 25664
rect 183614 25608 183619 25664
rect 144748 25606 183619 25608
rect 144748 25604 144754 25606
rect 183553 25603 183619 25606
rect 176326 25468 176332 25532
rect 176396 25530 176402 25532
rect 576853 25530 576919 25533
rect 176396 25528 576919 25530
rect 176396 25472 576858 25528
rect 576914 25472 576919 25528
rect 176396 25470 576919 25472
rect 176396 25468 176402 25470
rect 576853 25467 576919 25470
rect 145414 24380 145420 24444
rect 145484 24442 145490 24444
rect 201585 24442 201651 24445
rect 145484 24440 201651 24442
rect 145484 24384 201590 24440
rect 201646 24384 201651 24440
rect 145484 24382 201651 24384
rect 145484 24380 145490 24382
rect 201585 24379 201651 24382
rect 172094 24244 172100 24308
rect 172164 24306 172170 24308
rect 534073 24306 534139 24309
rect 172164 24304 534139 24306
rect 172164 24248 534078 24304
rect 534134 24248 534139 24304
rect 172164 24246 534139 24248
rect 172164 24244 172170 24246
rect 534073 24243 534139 24246
rect 171726 24108 171732 24172
rect 171796 24170 171802 24172
rect 538213 24170 538279 24173
rect 171796 24168 538279 24170
rect 171796 24112 538218 24168
rect 538274 24112 538279 24168
rect 171796 24110 538279 24112
rect 171796 24108 171802 24110
rect 538213 24107 538279 24110
rect 159030 23020 159036 23084
rect 159100 23082 159106 23084
rect 378133 23082 378199 23085
rect 159100 23080 378199 23082
rect 159100 23024 378138 23080
rect 378194 23024 378199 23080
rect 159100 23022 378199 23024
rect 159100 23020 159106 23022
rect 378133 23019 378199 23022
rect 162158 22884 162164 22948
rect 162228 22946 162234 22948
rect 414013 22946 414079 22949
rect 162228 22944 414079 22946
rect 162228 22888 414018 22944
rect 414074 22888 414079 22944
rect 162228 22886 414079 22888
rect 162228 22884 162234 22886
rect 414013 22883 414079 22886
rect 169518 22748 169524 22812
rect 169588 22810 169594 22812
rect 502333 22810 502399 22813
rect 169588 22808 502399 22810
rect 169588 22752 502338 22808
rect 502394 22752 502399 22808
rect 169588 22750 502399 22752
rect 169588 22748 169594 22750
rect 502333 22747 502399 22750
rect 63493 22674 63559 22677
rect 135662 22674 135668 22676
rect 63493 22672 135668 22674
rect 63493 22616 63498 22672
rect 63554 22616 135668 22672
rect 63493 22614 135668 22616
rect 63493 22611 63559 22614
rect 135662 22612 135668 22614
rect 135732 22612 135738 22676
rect 170622 22612 170628 22676
rect 170692 22674 170698 22676
rect 520273 22674 520339 22677
rect 170692 22672 520339 22674
rect 170692 22616 520278 22672
rect 520334 22616 520339 22672
rect 170692 22614 520339 22616
rect 170692 22612 170698 22614
rect 520273 22611 520339 22614
rect 95233 21314 95299 21317
rect 138238 21314 138244 21316
rect 95233 21312 138244 21314
rect 95233 21256 95238 21312
rect 95294 21256 138244 21312
rect 95233 21254 138244 21256
rect 95233 21251 95299 21254
rect 138238 21252 138244 21254
rect 138308 21252 138314 21316
rect 151486 20164 151492 20228
rect 151556 20226 151562 20228
rect 269113 20226 269179 20229
rect 151556 20224 269179 20226
rect 151556 20168 269118 20224
rect 269174 20168 269179 20224
rect 151556 20166 269179 20168
rect 151556 20164 151562 20166
rect 269113 20163 269179 20166
rect 157926 20028 157932 20092
rect 157996 20090 158002 20092
rect 357433 20090 357499 20093
rect 157996 20088 357499 20090
rect 157996 20032 357438 20088
rect 357494 20032 357499 20088
rect 157996 20030 357499 20032
rect 157996 20028 158002 20030
rect 357433 20027 357499 20030
rect 164918 19892 164924 19956
rect 164988 19954 164994 19956
rect 444373 19954 444439 19957
rect 164988 19952 444439 19954
rect 164988 19896 444378 19952
rect 444434 19896 444439 19952
rect 164988 19894 444439 19896
rect 164988 19892 164994 19894
rect 444373 19891 444439 19894
rect 579981 19818 580047 19821
rect 583520 19818 584960 19908
rect 579981 19816 584960 19818
rect 579981 19760 579986 19816
rect 580042 19760 584960 19816
rect 579981 19758 584960 19760
rect 579981 19755 580047 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3233 19410 3299 19413
rect -960 19408 3299 19410
rect -960 19352 3238 19408
rect 3294 19352 3299 19408
rect -960 19350 3299 19352
rect -960 19260 480 19350
rect 3233 19347 3299 19350
rect 147254 18668 147260 18732
rect 147324 18730 147330 18732
rect 216673 18730 216739 18733
rect 147324 18728 216739 18730
rect 147324 18672 216678 18728
rect 216734 18672 216739 18728
rect 147324 18670 216739 18672
rect 147324 18668 147330 18670
rect 216673 18667 216739 18670
rect 163630 18532 163636 18596
rect 163700 18594 163706 18596
rect 430573 18594 430639 18597
rect 163700 18592 430639 18594
rect 163700 18536 430578 18592
rect 430634 18536 430639 18592
rect 163700 18534 430639 18536
rect 163700 18532 163706 18534
rect 430573 18531 430639 18534
rect 162526 17716 162532 17780
rect 162596 17778 162602 17780
rect 408493 17778 408559 17781
rect 162596 17776 408559 17778
rect 162596 17720 408498 17776
rect 408554 17720 408559 17776
rect 162596 17718 408559 17720
rect 162596 17716 162602 17718
rect 408493 17715 408559 17718
rect 162342 17580 162348 17644
rect 162412 17642 162418 17644
rect 412633 17642 412699 17645
rect 162412 17640 412699 17642
rect 162412 17584 412638 17640
rect 412694 17584 412699 17640
rect 162412 17582 412699 17584
rect 162412 17580 162418 17582
rect 412633 17579 412699 17582
rect 166390 17444 166396 17508
rect 166460 17506 166466 17508
rect 466453 17506 466519 17509
rect 166460 17504 466519 17506
rect 166460 17448 466458 17504
rect 466514 17448 466519 17504
rect 166460 17446 466519 17448
rect 166460 17444 166466 17446
rect 466453 17443 466519 17446
rect 170806 17308 170812 17372
rect 170876 17370 170882 17372
rect 517513 17370 517579 17373
rect 170876 17368 517579 17370
rect 170876 17312 517518 17368
rect 517574 17312 517579 17368
rect 170876 17310 517579 17312
rect 170876 17308 170882 17310
rect 517513 17307 517579 17310
rect 176510 17172 176516 17236
rect 176580 17234 176586 17236
rect 580993 17234 581059 17237
rect 176580 17232 581059 17234
rect 176580 17176 580998 17232
rect 581054 17176 581059 17232
rect 176580 17174 581059 17176
rect 176580 17172 176586 17174
rect 580993 17171 581059 17174
rect 154246 16084 154252 16148
rect 154316 16146 154322 16148
rect 305545 16146 305611 16149
rect 154316 16144 305611 16146
rect 154316 16088 305550 16144
rect 305606 16088 305611 16144
rect 154316 16086 305611 16088
rect 154316 16084 154322 16086
rect 305545 16083 305611 16086
rect 160870 15948 160876 16012
rect 160940 16010 160946 16012
rect 395337 16010 395403 16013
rect 160940 16008 395403 16010
rect 160940 15952 395342 16008
rect 395398 15952 395403 16008
rect 160940 15950 395403 15952
rect 160940 15948 160946 15950
rect 395337 15947 395403 15950
rect 162710 15812 162716 15876
rect 162780 15874 162786 15876
rect 410793 15874 410859 15877
rect 162780 15872 410859 15874
rect 162780 15816 410798 15872
rect 410854 15816 410859 15872
rect 162780 15814 410859 15816
rect 162780 15812 162786 15814
rect 410793 15811 410859 15814
rect 158110 14860 158116 14924
rect 158180 14922 158186 14924
rect 356329 14922 356395 14925
rect 158180 14920 356395 14922
rect 158180 14864 356334 14920
rect 356390 14864 356395 14920
rect 158180 14862 356395 14864
rect 158180 14860 158186 14862
rect 356329 14859 356395 14862
rect 158294 14724 158300 14788
rect 158364 14786 158370 14788
rect 359457 14786 359523 14789
rect 158364 14784 359523 14786
rect 158364 14728 359462 14784
rect 359518 14728 359523 14784
rect 158364 14726 359523 14728
rect 158364 14724 158370 14726
rect 359457 14723 359523 14726
rect 161054 14588 161060 14652
rect 161124 14650 161130 14652
rect 394233 14650 394299 14653
rect 161124 14648 394299 14650
rect 161124 14592 394238 14648
rect 394294 14592 394299 14648
rect 161124 14590 394299 14592
rect 161124 14588 161130 14590
rect 394233 14587 394299 14590
rect 166574 14452 166580 14516
rect 166644 14514 166650 14516
rect 463969 14514 464035 14517
rect 166644 14512 464035 14514
rect 166644 14456 463974 14512
rect 464030 14456 464035 14512
rect 166644 14454 464035 14456
rect 166644 14452 166650 14454
rect 463969 14451 464035 14454
rect 156638 13092 156644 13156
rect 156708 13154 156714 13156
rect 340873 13154 340939 13157
rect 156708 13152 340939 13154
rect 156708 13096 340878 13152
rect 340934 13096 340939 13152
rect 156708 13094 340939 13096
rect 156708 13092 156714 13094
rect 340873 13091 340939 13094
rect 167862 12956 167868 13020
rect 167932 13018 167938 13020
rect 484761 13018 484827 13021
rect 167932 13016 484827 13018
rect 167932 12960 484766 13016
rect 484822 12960 484827 13016
rect 167932 12958 484827 12960
rect 167932 12956 167938 12958
rect 484761 12955 484827 12958
rect 155534 12276 155540 12340
rect 155604 12338 155610 12340
rect 324405 12338 324471 12341
rect 155604 12336 324471 12338
rect 155604 12280 324410 12336
rect 324466 12280 324471 12336
rect 155604 12278 324471 12280
rect 155604 12276 155610 12278
rect 324405 12275 324471 12278
rect 156822 12140 156828 12204
rect 156892 12202 156898 12204
rect 340965 12202 341031 12205
rect 156892 12200 341031 12202
rect 156892 12144 340970 12200
rect 341026 12144 341031 12200
rect 156892 12142 341031 12144
rect 156892 12140 156898 12142
rect 340965 12139 341031 12142
rect 158478 12004 158484 12068
rect 158548 12066 158554 12068
rect 357525 12066 357591 12069
rect 158548 12064 357591 12066
rect 158548 12008 357530 12064
rect 357586 12008 357591 12064
rect 158548 12006 357591 12008
rect 158548 12004 158554 12006
rect 357525 12003 357591 12006
rect 161238 11868 161244 11932
rect 161308 11930 161314 11932
rect 392577 11930 392643 11933
rect 161308 11928 392643 11930
rect 161308 11872 392582 11928
rect 392638 11872 392643 11928
rect 161308 11870 392643 11872
rect 161308 11868 161314 11870
rect 392577 11867 392643 11870
rect 165102 11732 165108 11796
rect 165172 11794 165178 11796
rect 448513 11794 448579 11797
rect 165172 11792 448579 11794
rect 165172 11736 448518 11792
rect 448574 11736 448579 11792
rect 165172 11734 448579 11736
rect 165172 11732 165178 11734
rect 448513 11731 448579 11734
rect 170990 11596 170996 11660
rect 171060 11658 171066 11660
rect 517145 11658 517211 11661
rect 171060 11656 517211 11658
rect 171060 11600 517150 11656
rect 517206 11600 517211 11656
rect 171060 11598 517211 11600
rect 171060 11596 171066 11598
rect 517145 11595 517211 11598
rect 152958 10372 152964 10436
rect 153028 10434 153034 10436
rect 288985 10434 289051 10437
rect 153028 10432 289051 10434
rect 153028 10376 288990 10432
rect 289046 10376 289051 10432
rect 153028 10374 289051 10376
rect 153028 10372 153034 10374
rect 288985 10371 289051 10374
rect 114001 10298 114067 10301
rect 139710 10298 139716 10300
rect 114001 10296 139716 10298
rect 114001 10240 114006 10296
rect 114062 10240 139716 10296
rect 114001 10238 139716 10240
rect 114001 10235 114067 10238
rect 139710 10236 139716 10238
rect 139780 10236 139786 10300
rect 168046 10236 168052 10300
rect 168116 10298 168122 10300
rect 481725 10298 481791 10301
rect 168116 10296 481791 10298
rect 168116 10240 481730 10296
rect 481786 10240 481791 10296
rect 168116 10238 481791 10240
rect 168116 10236 168122 10238
rect 481725 10235 481791 10238
rect 78581 9482 78647 9485
rect 137502 9482 137508 9484
rect 78581 9480 137508 9482
rect 78581 9424 78586 9480
rect 78642 9424 137508 9480
rect 78581 9422 137508 9424
rect 78581 9419 78647 9422
rect 137502 9420 137508 9422
rect 137572 9420 137578 9484
rect 60825 9346 60891 9349
rect 135478 9346 135484 9348
rect 60825 9344 135484 9346
rect 60825 9288 60830 9344
rect 60886 9288 135484 9344
rect 60825 9286 135484 9288
rect 60825 9283 60891 9286
rect 135478 9284 135484 9286
rect 135548 9284 135554 9348
rect 45461 9210 45527 9213
rect 134374 9210 134380 9212
rect 45461 9208 134380 9210
rect 45461 9152 45466 9208
rect 45522 9152 134380 9208
rect 45461 9150 134380 9152
rect 45461 9147 45527 9150
rect 134374 9148 134380 9150
rect 134444 9148 134450 9212
rect 151670 9148 151676 9212
rect 151740 9210 151746 9212
rect 271229 9210 271295 9213
rect 151740 9208 271295 9210
rect 151740 9152 271234 9208
rect 271290 9152 271295 9208
rect 151740 9150 271295 9152
rect 151740 9148 151746 9150
rect 271229 9147 271295 9150
rect 25313 9074 25379 9077
rect 133270 9074 133276 9076
rect 25313 9072 133276 9074
rect 25313 9016 25318 9072
rect 25374 9016 133276 9072
rect 25313 9014 133276 9016
rect 25313 9011 25379 9014
rect 133270 9012 133276 9014
rect 133340 9012 133346 9076
rect 157006 9012 157012 9076
rect 157076 9074 157082 9076
rect 343357 9074 343423 9077
rect 157076 9072 343423 9074
rect 157076 9016 343362 9072
rect 343418 9016 343423 9072
rect 157076 9014 343423 9016
rect 157076 9012 157082 9014
rect 343357 9011 343423 9014
rect 9949 8938 10015 8941
rect 131246 8938 131252 8940
rect 9949 8936 131252 8938
rect 9949 8880 9954 8936
rect 10010 8880 131252 8936
rect 9949 8878 131252 8880
rect 9949 8875 10015 8878
rect 131246 8876 131252 8878
rect 131316 8876 131322 8940
rect 166206 8876 166212 8940
rect 166276 8938 166282 8940
rect 466269 8938 466335 8941
rect 166276 8936 466335 8938
rect 166276 8880 466274 8936
rect 466330 8880 466335 8936
rect 166276 8878 466335 8880
rect 166276 8876 166282 8878
rect 466269 8875 466335 8878
rect 119889 7714 119955 7717
rect 139526 7714 139532 7716
rect 119889 7712 139532 7714
rect 119889 7656 119894 7712
rect 119950 7656 139532 7712
rect 119889 7654 139532 7656
rect 119889 7651 119955 7654
rect 139526 7652 139532 7654
rect 139596 7652 139602 7716
rect 27705 7578 27771 7581
rect 133086 7578 133092 7580
rect 27705 7576 133092 7578
rect 27705 7520 27710 7576
rect 27766 7520 133092 7576
rect 27705 7518 133092 7520
rect 27705 7515 27771 7518
rect 133086 7516 133092 7518
rect 133156 7516 133162 7580
rect 149830 7516 149836 7580
rect 149900 7578 149906 7580
rect 251265 7578 251331 7581
rect 149900 7576 251331 7578
rect 149900 7520 251270 7576
rect 251326 7520 251331 7576
rect 149900 7518 251331 7520
rect 149900 7516 149906 7518
rect 251265 7515 251331 7518
rect 145598 6836 145604 6900
rect 145668 6898 145674 6900
rect 235809 6898 235875 6901
rect 145668 6896 235875 6898
rect 145668 6840 235814 6896
rect 235870 6840 235875 6896
rect 145668 6838 235875 6840
rect 145668 6836 145674 6838
rect 235809 6835 235875 6838
rect 150014 6700 150020 6764
rect 150084 6762 150090 6764
rect 253473 6762 253539 6765
rect 150084 6760 253539 6762
rect 150084 6704 253478 6760
rect 253534 6704 253539 6760
rect 150084 6702 253539 6704
rect 150084 6700 150090 6702
rect 253473 6699 253539 6702
rect -960 6490 480 6580
rect 153878 6564 153884 6628
rect 153948 6626 153954 6628
rect 307937 6626 308003 6629
rect 153948 6624 308003 6626
rect 153948 6568 307942 6624
rect 307998 6568 308003 6624
rect 153948 6566 308003 6568
rect 153948 6564 153954 6566
rect 307937 6563 308003 6566
rect 580257 6626 580323 6629
rect 583520 6626 584960 6716
rect 580257 6624 584960 6626
rect 580257 6568 580262 6624
rect 580318 6568 584960 6624
rect 580257 6566 584960 6568
rect 580257 6563 580323 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 165286 6428 165292 6492
rect 165356 6490 165362 6492
rect 448605 6490 448671 6493
rect 165356 6488 448671 6490
rect 165356 6432 448610 6488
rect 448666 6432 448671 6488
rect 583520 6476 584960 6566
rect 165356 6430 448671 6432
rect 165356 6428 165362 6430
rect 448605 6427 448671 6430
rect 174854 6292 174860 6356
rect 174924 6354 174930 6356
rect 572713 6354 572779 6357
rect 174924 6352 572779 6354
rect 174924 6296 572718 6352
rect 572774 6296 572779 6352
rect 174924 6294 572779 6296
rect 174924 6292 174930 6294
rect 572713 6291 572779 6294
rect 63217 6218 63283 6221
rect 135294 6218 135300 6220
rect 63217 6216 135300 6218
rect 63217 6160 63222 6216
rect 63278 6160 135300 6216
rect 63217 6158 135300 6160
rect 63217 6155 63283 6158
rect 135294 6156 135300 6158
rect 135364 6156 135370 6220
rect 174670 6156 174676 6220
rect 174740 6218 174746 6220
rect 573909 6218 573975 6221
rect 174740 6216 573975 6218
rect 174740 6160 573914 6216
rect 573970 6160 573975 6216
rect 174740 6158 573975 6160
rect 174740 6156 174746 6158
rect 573909 6155 573975 6158
rect 148726 6020 148732 6084
rect 148796 6082 148802 6084
rect 232221 6082 232287 6085
rect 148796 6080 232287 6082
rect 148796 6024 232226 6080
rect 232282 6024 232287 6080
rect 148796 6022 232287 6024
rect 148796 6020 148802 6022
rect 232221 6019 232287 6022
rect 148910 5204 148916 5268
rect 148980 5266 148986 5268
rect 234613 5266 234679 5269
rect 148980 5264 234679 5266
rect 148980 5208 234618 5264
rect 234674 5208 234679 5264
rect 148980 5206 234679 5208
rect 148980 5204 148986 5206
rect 234613 5203 234679 5206
rect 157190 5068 157196 5132
rect 157260 5130 157266 5132
rect 338665 5130 338731 5133
rect 157260 5128 338731 5130
rect 157260 5072 338670 5128
rect 338726 5072 338731 5128
rect 157260 5070 338731 5072
rect 157260 5068 157266 5070
rect 338665 5067 338731 5070
rect 101029 4994 101095 4997
rect 138422 4994 138428 4996
rect 101029 4992 138428 4994
rect 101029 4936 101034 4992
rect 101090 4936 138428 4992
rect 101029 4934 138428 4936
rect 101029 4931 101095 4934
rect 138422 4932 138428 4934
rect 138492 4932 138498 4996
rect 143022 4932 143028 4996
rect 143092 4994 143098 4996
rect 162485 4994 162551 4997
rect 143092 4992 162551 4994
rect 143092 4936 162490 4992
rect 162546 4936 162551 4992
rect 143092 4934 162551 4936
rect 143092 4932 143098 4934
rect 162485 4931 162551 4934
rect 165470 4932 165476 4996
rect 165540 4994 165546 4996
rect 446213 4994 446279 4997
rect 165540 4992 446279 4994
rect 165540 4936 446218 4992
rect 446274 4936 446279 4992
rect 165540 4934 446279 4936
rect 165540 4932 165546 4934
rect 446213 4931 446279 4934
rect 8753 4858 8819 4861
rect 131614 4858 131620 4860
rect 8753 4856 131620 4858
rect 8753 4800 8758 4856
rect 8814 4800 131620 4856
rect 8753 4798 131620 4800
rect 8753 4795 8819 4798
rect 131614 4796 131620 4798
rect 131684 4796 131690 4860
rect 143206 4796 143212 4860
rect 143276 4858 143282 4860
rect 166073 4858 166139 4861
rect 143276 4856 166139 4858
rect 143276 4800 166078 4856
rect 166134 4800 166139 4856
rect 143276 4798 166139 4800
rect 143276 4796 143282 4798
rect 166073 4795 166139 4798
rect 175038 4796 175044 4860
rect 175108 4858 175114 4860
rect 570321 4858 570387 4861
rect 175108 4856 570387 4858
rect 175108 4800 570326 4856
rect 570382 4800 570387 4856
rect 175108 4798 570387 4800
rect 175108 4796 175114 4798
rect 570321 4795 570387 4798
rect 146886 3708 146892 3772
rect 146956 3770 146962 3772
rect 214465 3770 214531 3773
rect 146956 3768 214531 3770
rect 146956 3712 214470 3768
rect 214526 3712 214531 3768
rect 146956 3710 214531 3712
rect 146956 3708 146962 3710
rect 214465 3707 214531 3710
rect 139158 3572 139164 3636
rect 139228 3634 139234 3636
rect 218053 3634 218119 3637
rect 139228 3632 218119 3634
rect 139228 3576 218058 3632
rect 218114 3576 218119 3632
rect 139228 3574 218119 3576
rect 139228 3572 139234 3574
rect 218053 3571 218119 3574
rect 140998 3436 141004 3500
rect 141068 3498 141074 3500
rect 161289 3498 161355 3501
rect 141068 3496 161355 3498
rect 141068 3440 161294 3496
rect 161350 3440 161355 3496
rect 141068 3438 161355 3440
rect 141068 3436 141074 3438
rect 161289 3435 161355 3438
rect 175733 3498 175799 3501
rect 544377 3498 544443 3501
rect 175733 3496 544443 3498
rect 175733 3440 175738 3496
rect 175794 3440 544382 3496
rect 544438 3440 544443 3496
rect 175733 3438 544443 3440
rect 175733 3435 175799 3438
rect 544377 3435 544443 3438
rect 118785 3362 118851 3365
rect 139894 3362 139900 3364
rect 118785 3360 139900 3362
rect 118785 3304 118790 3360
rect 118846 3304 139900 3360
rect 118785 3302 139900 3304
rect 118785 3299 118851 3302
rect 139894 3300 139900 3302
rect 139964 3300 139970 3364
rect 143390 3300 143396 3364
rect 143460 3362 143466 3364
rect 163681 3362 163747 3365
rect 143460 3360 163747 3362
rect 143460 3304 163686 3360
rect 163742 3304 163747 3360
rect 143460 3302 163747 3304
rect 143460 3300 143466 3302
rect 163681 3299 163747 3302
rect 177062 3300 177068 3364
rect 177132 3362 177138 3364
rect 558545 3362 558611 3365
rect 177132 3360 558611 3362
rect 177132 3304 558550 3360
rect 558606 3304 558611 3360
rect 177132 3302 558611 3304
rect 177132 3300 177138 3302
rect 558545 3299 558611 3302
<< via3 >>
rect 176700 80956 176764 81020
rect 176884 80820 176948 80884
rect 177436 80548 177500 80612
rect 175228 80412 175292 80476
rect 134012 80140 134076 80204
rect 143212 80140 143276 80204
rect 131436 79868 131500 79932
rect 131436 79792 131500 79796
rect 131436 79736 131450 79792
rect 131450 79736 131500 79792
rect 131436 79732 131500 79736
rect 133276 80004 133340 80068
rect 149652 80140 149716 80204
rect 170628 80140 170692 80204
rect 161244 80004 161308 80068
rect 166764 80004 166828 80068
rect 132724 79928 132788 79932
rect 132724 79872 132728 79928
rect 132728 79872 132784 79928
rect 132784 79872 132788 79928
rect 132724 79868 132788 79872
rect 134564 79868 134628 79932
rect 134196 79732 134260 79796
rect 133644 79596 133708 79660
rect 135300 79868 135364 79932
rect 135484 79732 135548 79796
rect 137508 79868 137572 79932
rect 137876 79928 137940 79932
rect 137876 79872 137880 79928
rect 137880 79872 137936 79928
rect 137936 79872 137940 79928
rect 137876 79868 137940 79872
rect 135300 79460 135364 79524
rect 138060 79732 138124 79796
rect 138428 79792 138492 79796
rect 138428 79736 138432 79792
rect 138432 79736 138488 79792
rect 138488 79736 138492 79792
rect 138428 79732 138492 79736
rect 139716 79596 139780 79660
rect 139900 79656 139964 79660
rect 139900 79600 139914 79656
rect 139914 79600 139964 79656
rect 139900 79596 139964 79600
rect 141924 79894 141988 79932
rect 141924 79868 141928 79894
rect 141928 79868 141984 79894
rect 141984 79868 141988 79894
rect 143764 79928 143828 79932
rect 143764 79872 143768 79928
rect 143768 79872 143824 79928
rect 143824 79872 143828 79928
rect 143764 79868 143828 79872
rect 144500 79868 144564 79932
rect 142108 79596 142172 79660
rect 146892 79868 146956 79932
rect 147996 79928 148060 79932
rect 147996 79872 148000 79928
rect 148000 79872 148056 79928
rect 148056 79872 148060 79928
rect 147996 79868 148060 79872
rect 148180 79906 148184 79932
rect 148184 79906 148240 79932
rect 148240 79906 148244 79932
rect 148180 79868 148244 79906
rect 148916 79868 148980 79932
rect 143396 79732 143460 79796
rect 144684 79596 144748 79660
rect 148916 79792 148980 79796
rect 148916 79736 148930 79792
rect 148930 79736 148980 79792
rect 148916 79732 148980 79736
rect 150204 79792 150268 79796
rect 150204 79736 150218 79792
rect 150218 79736 150268 79792
rect 150204 79732 150268 79736
rect 151124 79906 151128 79932
rect 151128 79906 151184 79932
rect 151184 79906 151188 79932
rect 151124 79868 151188 79906
rect 151492 79868 151556 79932
rect 151676 79906 151680 79932
rect 151680 79906 151736 79932
rect 151736 79906 151740 79932
rect 151676 79868 151740 79906
rect 151308 79732 151372 79796
rect 152780 79868 152844 79932
rect 153700 79906 153704 79932
rect 153704 79906 153760 79932
rect 153760 79906 153764 79932
rect 153700 79868 153764 79906
rect 154436 79868 154500 79932
rect 154620 79928 154684 79932
rect 154620 79872 154624 79928
rect 154624 79872 154680 79928
rect 154680 79872 154684 79928
rect 154620 79868 154684 79872
rect 155356 79868 155420 79932
rect 155540 79868 155604 79932
rect 156276 79868 156340 79932
rect 156828 79868 156892 79932
rect 158116 79868 158180 79932
rect 159588 79868 159652 79932
rect 154068 79732 154132 79796
rect 157196 79460 157260 79524
rect 158300 79732 158364 79796
rect 160692 79868 160756 79932
rect 161980 79868 162044 79932
rect 162348 79868 162412 79932
rect 163268 79868 163332 79932
rect 158852 79596 158916 79660
rect 161060 79732 161124 79796
rect 164740 79868 164804 79932
rect 164004 79732 164068 79796
rect 165108 79732 165172 79796
rect 165476 79792 165540 79796
rect 165476 79736 165526 79792
rect 165526 79736 165540 79792
rect 165476 79732 165540 79736
rect 167316 79928 167380 79932
rect 167316 79872 167320 79928
rect 167320 79872 167376 79928
rect 167376 79872 167380 79928
rect 167316 79868 167380 79872
rect 168052 79928 168116 79932
rect 168052 79872 168056 79928
rect 168056 79872 168112 79928
rect 168112 79872 168116 79928
rect 168052 79868 168116 79872
rect 167684 79732 167748 79796
rect 168972 79906 168976 79932
rect 168976 79906 169032 79932
rect 169032 79906 169036 79932
rect 168972 79868 169036 79906
rect 170260 79906 170264 79932
rect 170264 79906 170320 79932
rect 170320 79906 170324 79932
rect 170260 79868 170324 79906
rect 171548 80004 171612 80068
rect 171732 79928 171796 79932
rect 171732 79872 171736 79928
rect 171736 79872 171792 79928
rect 171792 79872 171796 79928
rect 171732 79868 171796 79872
rect 177804 80140 177868 80204
rect 172652 79928 172716 79932
rect 172652 79872 172656 79928
rect 172656 79872 172712 79928
rect 172712 79872 172716 79928
rect 172652 79868 172716 79872
rect 173204 79868 173268 79932
rect 170812 79732 170876 79796
rect 172100 79596 172164 79660
rect 173388 79732 173452 79796
rect 159588 79460 159652 79524
rect 160876 79460 160940 79524
rect 164556 79460 164620 79524
rect 167868 79460 167932 79524
rect 169340 79520 169404 79524
rect 169340 79464 169390 79520
rect 169390 79464 169404 79520
rect 169340 79460 169404 79464
rect 169524 79460 169588 79524
rect 170444 79460 170508 79524
rect 174676 79868 174740 79932
rect 176332 79868 176396 79932
rect 176148 79732 176212 79796
rect 176884 79732 176948 79796
rect 175044 79596 175108 79660
rect 175228 79656 175292 79660
rect 175228 79600 175242 79656
rect 175242 79600 175292 79656
rect 175228 79596 175292 79600
rect 177436 79596 177500 79660
rect 177068 79460 177132 79524
rect 177804 79928 177868 79932
rect 177804 79872 177808 79928
rect 177808 79872 177864 79928
rect 177864 79872 177868 79928
rect 177804 79868 177868 79872
rect 178356 79928 178420 79932
rect 178356 79872 178360 79928
rect 178360 79872 178416 79928
rect 178416 79872 178420 79928
rect 178356 79868 178420 79872
rect 176700 79384 176764 79388
rect 176700 79328 176714 79384
rect 176714 79328 176764 79384
rect 176700 79324 176764 79328
rect 178356 79188 178420 79252
rect 131252 78916 131316 78980
rect 141924 78916 141988 78980
rect 163636 78916 163700 78980
rect 173572 78976 173636 78980
rect 173572 78920 173622 78976
rect 173622 78920 173636 78976
rect 173572 78916 173636 78920
rect 175228 78916 175292 78980
rect 175780 78916 175844 78980
rect 176148 78916 176212 78980
rect 176516 78916 176580 78980
rect 133460 78644 133524 78708
rect 138244 78644 138308 78708
rect 150020 78644 150084 78708
rect 157932 78644 157996 78708
rect 163452 78644 163516 78708
rect 168972 78644 169036 78708
rect 170996 78644 171060 78708
rect 173388 78644 173452 78708
rect 173756 78704 173820 78708
rect 173756 78648 173806 78704
rect 173806 78648 173820 78704
rect 173756 78644 173820 78648
rect 174860 78644 174924 78708
rect 176148 78644 176212 78708
rect 133644 78372 133708 78436
rect 137876 78372 137940 78436
rect 144500 78372 144564 78436
rect 151492 78372 151556 78436
rect 162532 78236 162596 78300
rect 164004 78236 164068 78300
rect 171732 78236 171796 78300
rect 134564 78100 134628 78164
rect 143764 78100 143828 78164
rect 144684 78100 144748 78164
rect 155356 78100 155420 78164
rect 172284 78160 172348 78164
rect 172284 78104 172298 78160
rect 172298 78104 172348 78160
rect 172284 78100 172348 78104
rect 172652 78100 172716 78164
rect 173204 78100 173268 78164
rect 131068 77964 131132 78028
rect 134196 77964 134260 78028
rect 135300 77964 135364 78028
rect 135668 78024 135732 78028
rect 135668 77968 135682 78024
rect 135682 77968 135732 78024
rect 135668 77964 135732 77968
rect 139164 77964 139228 78028
rect 164924 77964 164988 78028
rect 165476 78024 165540 78028
rect 165476 77968 165526 78024
rect 165526 77968 165540 78024
rect 165476 77964 165540 77968
rect 164556 77828 164620 77892
rect 170260 77692 170324 77756
rect 156644 77556 156708 77620
rect 161980 77556 162044 77620
rect 166396 77556 166460 77620
rect 145420 77420 145484 77484
rect 147076 77420 147140 77484
rect 152412 77420 152476 77484
rect 154252 77420 154316 77484
rect 157012 77420 157076 77484
rect 166764 77480 166828 77484
rect 166764 77424 166778 77480
rect 166778 77424 166828 77480
rect 166764 77420 166828 77424
rect 172100 77480 172164 77484
rect 172100 77424 172150 77480
rect 172150 77424 172164 77480
rect 172100 77420 172164 77424
rect 145236 77284 145300 77348
rect 147260 77284 147324 77348
rect 152780 77284 152844 77348
rect 153700 77284 153764 77348
rect 154068 77284 154132 77348
rect 154620 77284 154684 77348
rect 156276 77344 156340 77348
rect 156276 77288 156326 77344
rect 156326 77288 156340 77344
rect 156276 77284 156340 77288
rect 158484 77284 158548 77348
rect 159036 77284 159100 77348
rect 166212 77284 166276 77348
rect 167316 77284 167380 77348
rect 138060 76740 138124 76804
rect 143028 76740 143092 76804
rect 142844 76604 142908 76668
rect 144316 76604 144380 76668
rect 147996 76604 148060 76668
rect 148548 76604 148612 76668
rect 151124 76604 151188 76668
rect 151492 76604 151556 76668
rect 154436 76604 154500 76668
rect 131436 76468 131500 76532
rect 141004 76468 141068 76532
rect 160692 76468 160756 76532
rect 162164 76196 162228 76260
rect 164740 76256 164804 76260
rect 164740 76200 164754 76256
rect 164754 76200 164804 76256
rect 164740 76196 164804 76200
rect 162716 76060 162780 76124
rect 166764 75652 166828 75716
rect 148180 75380 148244 75444
rect 163268 75380 163332 75444
rect 133828 75244 133892 75308
rect 139532 75244 139596 75308
rect 140820 75244 140884 75308
rect 131068 75108 131132 75172
rect 145604 75108 145668 75172
rect 172284 75108 172348 75172
rect 142108 74972 142172 75036
rect 175780 74428 175844 74492
rect 134196 73884 134260 73948
rect 149652 73884 149716 73948
rect 133460 73748 133524 73812
rect 152412 73748 152476 73812
rect 175228 71028 175292 71092
rect 144316 69532 144380 69596
rect 158852 68172 158916 68236
rect 176148 66812 176212 66876
rect 142844 66132 142908 66196
rect 144500 65452 144564 65516
rect 171916 65452 171980 65516
rect 167684 64228 167748 64292
rect 173572 64092 173636 64156
rect 169340 63548 169404 63612
rect 145236 62732 145300 62796
rect 170444 61372 170508 61436
rect 154068 55796 154132 55860
rect 173756 46140 173820 46204
rect 140820 44236 140884 44300
rect 163452 36484 163516 36548
rect 151308 30908 151372 30972
rect 148548 29548 148612 29612
rect 147076 28188 147140 28252
rect 152780 26828 152844 26892
rect 144684 25604 144748 25668
rect 176332 25468 176396 25532
rect 145420 24380 145484 24444
rect 172100 24244 172164 24308
rect 171732 24108 171796 24172
rect 159036 23020 159100 23084
rect 162164 22884 162228 22948
rect 169524 22748 169588 22812
rect 135668 22612 135732 22676
rect 170628 22612 170692 22676
rect 138244 21252 138308 21316
rect 151492 20164 151556 20228
rect 157932 20028 157996 20092
rect 164924 19892 164988 19956
rect 147260 18668 147324 18732
rect 163636 18532 163700 18596
rect 162532 17716 162596 17780
rect 162348 17580 162412 17644
rect 166396 17444 166460 17508
rect 170812 17308 170876 17372
rect 176516 17172 176580 17236
rect 154252 16084 154316 16148
rect 160876 15948 160940 16012
rect 162716 15812 162780 15876
rect 158116 14860 158180 14924
rect 158300 14724 158364 14788
rect 161060 14588 161124 14652
rect 166580 14452 166644 14516
rect 156644 13092 156708 13156
rect 167868 12956 167932 13020
rect 155540 12276 155604 12340
rect 156828 12140 156892 12204
rect 158484 12004 158548 12068
rect 161244 11868 161308 11932
rect 165108 11732 165172 11796
rect 170996 11596 171060 11660
rect 152964 10372 153028 10436
rect 139716 10236 139780 10300
rect 168052 10236 168116 10300
rect 137508 9420 137572 9484
rect 135484 9284 135548 9348
rect 134380 9148 134444 9212
rect 151676 9148 151740 9212
rect 133276 9012 133340 9076
rect 157012 9012 157076 9076
rect 131252 8876 131316 8940
rect 166212 8876 166276 8940
rect 139532 7652 139596 7716
rect 133092 7516 133156 7580
rect 149836 7516 149900 7580
rect 145604 6836 145668 6900
rect 150020 6700 150084 6764
rect 153884 6564 153948 6628
rect 165292 6428 165356 6492
rect 174860 6292 174924 6356
rect 135300 6156 135364 6220
rect 174676 6156 174740 6220
rect 148732 6020 148796 6084
rect 148916 5204 148980 5268
rect 157196 5068 157260 5132
rect 138428 4932 138492 4996
rect 143028 4932 143092 4996
rect 165476 4932 165540 4996
rect 131620 4796 131684 4860
rect 143212 4796 143276 4860
rect 175044 4796 175108 4860
rect 146892 3708 146956 3772
rect 139164 3572 139228 3636
rect 141004 3436 141068 3500
rect 139900 3300 139964 3364
rect 143396 3300 143460 3364
rect 177068 3300 177132 3364
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 682954 -8106 711002
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 -8106 682954
rect -8726 682634 -8106 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 -8106 682634
rect -8726 646954 -8106 682398
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 -8106 646954
rect -8726 646634 -8106 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 -8106 646634
rect -8726 610954 -8106 646398
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 -8106 610954
rect -8726 610634 -8106 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 -8106 610634
rect -8726 574954 -8106 610398
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 -8106 574954
rect -8726 574634 -8106 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 -8106 574634
rect -8726 538954 -8106 574398
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 -8106 538954
rect -8726 538634 -8106 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 -8106 538634
rect -8726 502954 -8106 538398
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 -8106 502954
rect -8726 502634 -8106 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 -8106 502634
rect -8726 466954 -8106 502398
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 -8106 466954
rect -8726 466634 -8106 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 -8106 466634
rect -8726 430954 -8106 466398
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 -8106 430954
rect -8726 430634 -8106 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 -8106 430634
rect -8726 394954 -8106 430398
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 -8106 394954
rect -8726 394634 -8106 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 -8106 394634
rect -8726 358954 -8106 394398
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 -8106 358954
rect -8726 358634 -8106 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 -8106 358634
rect -8726 322954 -8106 358398
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 -8106 322954
rect -8726 322634 -8106 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 -8106 322634
rect -8726 286954 -8106 322398
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 -8106 286954
rect -8726 286634 -8106 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 -8106 286634
rect -8726 250954 -8106 286398
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 -8106 250954
rect -8726 250634 -8106 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 -8106 250634
rect -8726 214954 -8106 250398
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 -8106 214954
rect -8726 214634 -8106 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 -8106 214634
rect -8726 178954 -8106 214398
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 -8106 178954
rect -8726 178634 -8106 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 -8106 178634
rect -8726 142954 -8106 178398
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 -8106 142954
rect -8726 142634 -8106 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 -8106 142634
rect -8726 106954 -8106 142398
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 -8106 106954
rect -8726 106634 -8106 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 -8106 106634
rect -8726 70954 -8106 106398
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 -8106 70954
rect -8726 70634 -8106 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 -8106 70634
rect -8726 34954 -8106 70398
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 -8106 34954
rect -8726 34634 -8106 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 -8106 34634
rect -8726 -7066 -8106 34398
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 678454 -7146 710042
rect -7766 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 -7146 678454
rect -7766 678134 -7146 678218
rect -7766 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 -7146 678134
rect -7766 642454 -7146 677898
rect -7766 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 -7146 642454
rect -7766 642134 -7146 642218
rect -7766 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 -7146 642134
rect -7766 606454 -7146 641898
rect -7766 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 -7146 606454
rect -7766 606134 -7146 606218
rect -7766 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 -7146 606134
rect -7766 570454 -7146 605898
rect -7766 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 -7146 570454
rect -7766 570134 -7146 570218
rect -7766 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 -7146 570134
rect -7766 534454 -7146 569898
rect -7766 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 -7146 534454
rect -7766 534134 -7146 534218
rect -7766 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 -7146 534134
rect -7766 498454 -7146 533898
rect -7766 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 -7146 498454
rect -7766 498134 -7146 498218
rect -7766 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 -7146 498134
rect -7766 462454 -7146 497898
rect -7766 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 -7146 462454
rect -7766 462134 -7146 462218
rect -7766 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 -7146 462134
rect -7766 426454 -7146 461898
rect -7766 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 -7146 426454
rect -7766 426134 -7146 426218
rect -7766 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 -7146 426134
rect -7766 390454 -7146 425898
rect -7766 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 -7146 390454
rect -7766 390134 -7146 390218
rect -7766 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 -7146 390134
rect -7766 354454 -7146 389898
rect -7766 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 -7146 354454
rect -7766 354134 -7146 354218
rect -7766 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 -7146 354134
rect -7766 318454 -7146 353898
rect -7766 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 -7146 318454
rect -7766 318134 -7146 318218
rect -7766 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 -7146 318134
rect -7766 282454 -7146 317898
rect -7766 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 -7146 282454
rect -7766 282134 -7146 282218
rect -7766 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 -7146 282134
rect -7766 246454 -7146 281898
rect -7766 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 -7146 246454
rect -7766 246134 -7146 246218
rect -7766 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 -7146 246134
rect -7766 210454 -7146 245898
rect -7766 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 -7146 210454
rect -7766 210134 -7146 210218
rect -7766 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 -7146 210134
rect -7766 174454 -7146 209898
rect -7766 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 -7146 174454
rect -7766 174134 -7146 174218
rect -7766 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 -7146 174134
rect -7766 138454 -7146 173898
rect -7766 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 -7146 138454
rect -7766 138134 -7146 138218
rect -7766 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 -7146 138134
rect -7766 102454 -7146 137898
rect -7766 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 -7146 102454
rect -7766 102134 -7146 102218
rect -7766 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 -7146 102134
rect -7766 66454 -7146 101898
rect -7766 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 -7146 66454
rect -7766 66134 -7146 66218
rect -7766 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 -7146 66134
rect -7766 30454 -7146 65898
rect -7766 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 -7146 30454
rect -7766 30134 -7146 30218
rect -7766 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 -7146 30134
rect -7766 -6106 -7146 29898
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 673954 -6186 709082
rect -6806 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 -6186 673954
rect -6806 673634 -6186 673718
rect -6806 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 -6186 673634
rect -6806 637954 -6186 673398
rect -6806 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 -6186 637954
rect -6806 637634 -6186 637718
rect -6806 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 -6186 637634
rect -6806 601954 -6186 637398
rect -6806 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 -6186 601954
rect -6806 601634 -6186 601718
rect -6806 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 -6186 601634
rect -6806 565954 -6186 601398
rect -6806 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 -6186 565954
rect -6806 565634 -6186 565718
rect -6806 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 -6186 565634
rect -6806 529954 -6186 565398
rect -6806 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 -6186 529954
rect -6806 529634 -6186 529718
rect -6806 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 -6186 529634
rect -6806 493954 -6186 529398
rect -6806 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 -6186 493954
rect -6806 493634 -6186 493718
rect -6806 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 -6186 493634
rect -6806 457954 -6186 493398
rect -6806 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 -6186 457954
rect -6806 457634 -6186 457718
rect -6806 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 -6186 457634
rect -6806 421954 -6186 457398
rect -6806 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 -6186 421954
rect -6806 421634 -6186 421718
rect -6806 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 -6186 421634
rect -6806 385954 -6186 421398
rect -6806 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 -6186 385954
rect -6806 385634 -6186 385718
rect -6806 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 -6186 385634
rect -6806 349954 -6186 385398
rect -6806 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 -6186 349954
rect -6806 349634 -6186 349718
rect -6806 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 -6186 349634
rect -6806 313954 -6186 349398
rect -6806 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 -6186 313954
rect -6806 313634 -6186 313718
rect -6806 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 -6186 313634
rect -6806 277954 -6186 313398
rect -6806 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 -6186 277954
rect -6806 277634 -6186 277718
rect -6806 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 -6186 277634
rect -6806 241954 -6186 277398
rect -6806 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 -6186 241954
rect -6806 241634 -6186 241718
rect -6806 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 -6186 241634
rect -6806 205954 -6186 241398
rect -6806 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 -6186 205954
rect -6806 205634 -6186 205718
rect -6806 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 -6186 205634
rect -6806 169954 -6186 205398
rect -6806 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 -6186 169954
rect -6806 169634 -6186 169718
rect -6806 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 -6186 169634
rect -6806 133954 -6186 169398
rect -6806 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 -6186 133954
rect -6806 133634 -6186 133718
rect -6806 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 -6186 133634
rect -6806 97954 -6186 133398
rect -6806 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 -6186 97954
rect -6806 97634 -6186 97718
rect -6806 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 -6186 97634
rect -6806 61954 -6186 97398
rect -6806 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 -6186 61954
rect -6806 61634 -6186 61718
rect -6806 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 -6186 61634
rect -6806 25954 -6186 61398
rect -6806 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 -6186 25954
rect -6806 25634 -6186 25718
rect -6806 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 -6186 25634
rect -6806 -5146 -6186 25398
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 669454 -5226 708122
rect -5846 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 -5226 669454
rect -5846 669134 -5226 669218
rect -5846 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 -5226 669134
rect -5846 633454 -5226 668898
rect -5846 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 -5226 633454
rect -5846 633134 -5226 633218
rect -5846 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 -5226 633134
rect -5846 597454 -5226 632898
rect -5846 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 -5226 597454
rect -5846 597134 -5226 597218
rect -5846 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 -5226 597134
rect -5846 561454 -5226 596898
rect -5846 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 -5226 561454
rect -5846 561134 -5226 561218
rect -5846 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 -5226 561134
rect -5846 525454 -5226 560898
rect -5846 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 -5226 525454
rect -5846 525134 -5226 525218
rect -5846 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 -5226 525134
rect -5846 489454 -5226 524898
rect -5846 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 -5226 489454
rect -5846 489134 -5226 489218
rect -5846 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 -5226 489134
rect -5846 453454 -5226 488898
rect -5846 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 -5226 453454
rect -5846 453134 -5226 453218
rect -5846 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 -5226 453134
rect -5846 417454 -5226 452898
rect -5846 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 -5226 417454
rect -5846 417134 -5226 417218
rect -5846 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 -5226 417134
rect -5846 381454 -5226 416898
rect -5846 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 -5226 381454
rect -5846 381134 -5226 381218
rect -5846 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 -5226 381134
rect -5846 345454 -5226 380898
rect -5846 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 -5226 345454
rect -5846 345134 -5226 345218
rect -5846 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 -5226 345134
rect -5846 309454 -5226 344898
rect -5846 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 -5226 309454
rect -5846 309134 -5226 309218
rect -5846 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 -5226 309134
rect -5846 273454 -5226 308898
rect -5846 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 -5226 273454
rect -5846 273134 -5226 273218
rect -5846 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 -5226 273134
rect -5846 237454 -5226 272898
rect -5846 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 -5226 237454
rect -5846 237134 -5226 237218
rect -5846 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 -5226 237134
rect -5846 201454 -5226 236898
rect -5846 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 -5226 201454
rect -5846 201134 -5226 201218
rect -5846 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 -5226 201134
rect -5846 165454 -5226 200898
rect -5846 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 -5226 165454
rect -5846 165134 -5226 165218
rect -5846 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 -5226 165134
rect -5846 129454 -5226 164898
rect -5846 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 -5226 129454
rect -5846 129134 -5226 129218
rect -5846 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 -5226 129134
rect -5846 93454 -5226 128898
rect -5846 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 -5226 93454
rect -5846 93134 -5226 93218
rect -5846 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 -5226 93134
rect -5846 57454 -5226 92898
rect -5846 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 -5226 57454
rect -5846 57134 -5226 57218
rect -5846 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 -5226 57134
rect -5846 21454 -5226 56898
rect -5846 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 -5226 21454
rect -5846 21134 -5226 21218
rect -5846 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 -5226 21134
rect -5846 -4186 -5226 20898
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 700954 -4266 707162
rect -4886 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 -4266 700954
rect -4886 700634 -4266 700718
rect -4886 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 -4266 700634
rect -4886 664954 -4266 700398
rect -4886 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 -4266 664954
rect -4886 664634 -4266 664718
rect -4886 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 -4266 664634
rect -4886 628954 -4266 664398
rect -4886 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 -4266 628954
rect -4886 628634 -4266 628718
rect -4886 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 -4266 628634
rect -4886 592954 -4266 628398
rect -4886 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 -4266 592954
rect -4886 592634 -4266 592718
rect -4886 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 -4266 592634
rect -4886 556954 -4266 592398
rect -4886 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 -4266 556954
rect -4886 556634 -4266 556718
rect -4886 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 -4266 556634
rect -4886 520954 -4266 556398
rect -4886 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 -4266 520954
rect -4886 520634 -4266 520718
rect -4886 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 -4266 520634
rect -4886 484954 -4266 520398
rect -4886 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 -4266 484954
rect -4886 484634 -4266 484718
rect -4886 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 -4266 484634
rect -4886 448954 -4266 484398
rect -4886 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 -4266 448954
rect -4886 448634 -4266 448718
rect -4886 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 -4266 448634
rect -4886 412954 -4266 448398
rect -4886 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 -4266 412954
rect -4886 412634 -4266 412718
rect -4886 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 -4266 412634
rect -4886 376954 -4266 412398
rect -4886 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 -4266 376954
rect -4886 376634 -4266 376718
rect -4886 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 -4266 376634
rect -4886 340954 -4266 376398
rect -4886 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 -4266 340954
rect -4886 340634 -4266 340718
rect -4886 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 -4266 340634
rect -4886 304954 -4266 340398
rect -4886 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 -4266 304954
rect -4886 304634 -4266 304718
rect -4886 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 -4266 304634
rect -4886 268954 -4266 304398
rect -4886 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 -4266 268954
rect -4886 268634 -4266 268718
rect -4886 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 -4266 268634
rect -4886 232954 -4266 268398
rect -4886 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 -4266 232954
rect -4886 232634 -4266 232718
rect -4886 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 -4266 232634
rect -4886 196954 -4266 232398
rect -4886 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 -4266 196954
rect -4886 196634 -4266 196718
rect -4886 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 -4266 196634
rect -4886 160954 -4266 196398
rect -4886 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 -4266 160954
rect -4886 160634 -4266 160718
rect -4886 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 -4266 160634
rect -4886 124954 -4266 160398
rect -4886 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 -4266 124954
rect -4886 124634 -4266 124718
rect -4886 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 -4266 124634
rect -4886 88954 -4266 124398
rect -4886 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 -4266 88954
rect -4886 88634 -4266 88718
rect -4886 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 -4266 88634
rect -4886 52954 -4266 88398
rect -4886 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 -4266 52954
rect -4886 52634 -4266 52718
rect -4886 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 -4266 52634
rect -4886 16954 -4266 52398
rect -4886 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 -4266 16954
rect -4886 16634 -4266 16718
rect -4886 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 -4266 16634
rect -4886 -3226 -4266 16398
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 696454 -3306 706202
rect -3926 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 -3306 696454
rect -3926 696134 -3306 696218
rect -3926 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 -3306 696134
rect -3926 660454 -3306 695898
rect -3926 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 -3306 660454
rect -3926 660134 -3306 660218
rect -3926 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 -3306 660134
rect -3926 624454 -3306 659898
rect -3926 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 -3306 624454
rect -3926 624134 -3306 624218
rect -3926 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 -3306 624134
rect -3926 588454 -3306 623898
rect -3926 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 -3306 588454
rect -3926 588134 -3306 588218
rect -3926 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 -3306 588134
rect -3926 552454 -3306 587898
rect -3926 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 -3306 552454
rect -3926 552134 -3306 552218
rect -3926 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 -3306 552134
rect -3926 516454 -3306 551898
rect -3926 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 -3306 516454
rect -3926 516134 -3306 516218
rect -3926 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 -3306 516134
rect -3926 480454 -3306 515898
rect -3926 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 -3306 480454
rect -3926 480134 -3306 480218
rect -3926 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 -3306 480134
rect -3926 444454 -3306 479898
rect -3926 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 -3306 444454
rect -3926 444134 -3306 444218
rect -3926 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 -3306 444134
rect -3926 408454 -3306 443898
rect -3926 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 -3306 408454
rect -3926 408134 -3306 408218
rect -3926 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 -3306 408134
rect -3926 372454 -3306 407898
rect -3926 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 -3306 372454
rect -3926 372134 -3306 372218
rect -3926 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 -3306 372134
rect -3926 336454 -3306 371898
rect -3926 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 -3306 336454
rect -3926 336134 -3306 336218
rect -3926 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 -3306 336134
rect -3926 300454 -3306 335898
rect -3926 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 -3306 300454
rect -3926 300134 -3306 300218
rect -3926 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 -3306 300134
rect -3926 264454 -3306 299898
rect -3926 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 -3306 264454
rect -3926 264134 -3306 264218
rect -3926 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 -3306 264134
rect -3926 228454 -3306 263898
rect -3926 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 -3306 228454
rect -3926 228134 -3306 228218
rect -3926 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 -3306 228134
rect -3926 192454 -3306 227898
rect -3926 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 -3306 192454
rect -3926 192134 -3306 192218
rect -3926 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 -3306 192134
rect -3926 156454 -3306 191898
rect -3926 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 -3306 156454
rect -3926 156134 -3306 156218
rect -3926 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 -3306 156134
rect -3926 120454 -3306 155898
rect -3926 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 -3306 120454
rect -3926 120134 -3306 120218
rect -3926 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 -3306 120134
rect -3926 84454 -3306 119898
rect -3926 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 -3306 84454
rect -3926 84134 -3306 84218
rect -3926 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 -3306 84134
rect -3926 48454 -3306 83898
rect -3926 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 -3306 48454
rect -3926 48134 -3306 48218
rect -3926 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 -3306 48134
rect -3926 12454 -3306 47898
rect -3926 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 -3306 12454
rect -3926 12134 -3306 12218
rect -3926 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 -3306 12134
rect -3926 -2266 -3306 11898
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691954 -2346 705242
rect -2966 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 -2346 691954
rect -2966 691634 -2346 691718
rect -2966 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 -2346 691634
rect -2966 655954 -2346 691398
rect -2966 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 -2346 655954
rect -2966 655634 -2346 655718
rect -2966 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 -2346 655634
rect -2966 619954 -2346 655398
rect -2966 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 -2346 619954
rect -2966 619634 -2346 619718
rect -2966 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 -2346 619634
rect -2966 583954 -2346 619398
rect -2966 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 -2346 583954
rect -2966 583634 -2346 583718
rect -2966 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 -2346 583634
rect -2966 547954 -2346 583398
rect -2966 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 -2346 547954
rect -2966 547634 -2346 547718
rect -2966 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 -2346 547634
rect -2966 511954 -2346 547398
rect -2966 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 -2346 511954
rect -2966 511634 -2346 511718
rect -2966 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 -2346 511634
rect -2966 475954 -2346 511398
rect -2966 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 -2346 475954
rect -2966 475634 -2346 475718
rect -2966 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 -2346 475634
rect -2966 439954 -2346 475398
rect -2966 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 -2346 439954
rect -2966 439634 -2346 439718
rect -2966 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 -2346 439634
rect -2966 403954 -2346 439398
rect -2966 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 -2346 403954
rect -2966 403634 -2346 403718
rect -2966 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 -2346 403634
rect -2966 367954 -2346 403398
rect -2966 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 -2346 367954
rect -2966 367634 -2346 367718
rect -2966 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 -2346 367634
rect -2966 331954 -2346 367398
rect -2966 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 -2346 331954
rect -2966 331634 -2346 331718
rect -2966 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 -2346 331634
rect -2966 295954 -2346 331398
rect -2966 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 -2346 295954
rect -2966 295634 -2346 295718
rect -2966 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 -2346 295634
rect -2966 259954 -2346 295398
rect -2966 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 -2346 259954
rect -2966 259634 -2346 259718
rect -2966 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 -2346 259634
rect -2966 223954 -2346 259398
rect -2966 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 -2346 223954
rect -2966 223634 -2346 223718
rect -2966 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 -2346 223634
rect -2966 187954 -2346 223398
rect -2966 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 -2346 187954
rect -2966 187634 -2346 187718
rect -2966 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 -2346 187634
rect -2966 151954 -2346 187398
rect -2966 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 -2346 151954
rect -2966 151634 -2346 151718
rect -2966 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 -2346 151634
rect -2966 115954 -2346 151398
rect -2966 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 -2346 115954
rect -2966 115634 -2346 115718
rect -2966 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 -2346 115634
rect -2966 79954 -2346 115398
rect -2966 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 -2346 79954
rect -2966 79634 -2346 79718
rect -2966 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 -2346 79634
rect -2966 43954 -2346 79398
rect -2966 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 -2346 43954
rect -2966 43634 -2346 43718
rect -2966 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 -2346 43634
rect -2966 7954 -2346 43398
rect -2966 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 -2346 7954
rect -2966 7634 -2346 7718
rect -2966 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 -2346 7634
rect -2966 -1306 -2346 7398
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 6294 705798 6914 711590
rect 6294 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 6914 705798
rect 6294 705478 6914 705562
rect 6294 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 6914 705478
rect 6294 691954 6914 705242
rect 6294 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 6914 691954
rect 6294 691634 6914 691718
rect 6294 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 6914 691634
rect 6294 655954 6914 691398
rect 6294 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 6914 655954
rect 6294 655634 6914 655718
rect 6294 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 6914 655634
rect 6294 619954 6914 655398
rect 6294 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 6914 619954
rect 6294 619634 6914 619718
rect 6294 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 6914 619634
rect 6294 583954 6914 619398
rect 6294 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 6914 583954
rect 6294 583634 6914 583718
rect 6294 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 6914 583634
rect 6294 547954 6914 583398
rect 6294 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 6914 547954
rect 6294 547634 6914 547718
rect 6294 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 6914 547634
rect 6294 511954 6914 547398
rect 6294 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 6914 511954
rect 6294 511634 6914 511718
rect 6294 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 6914 511634
rect 6294 475954 6914 511398
rect 6294 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 6914 475954
rect 6294 475634 6914 475718
rect 6294 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 6914 475634
rect 6294 439954 6914 475398
rect 6294 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 6914 439954
rect 6294 439634 6914 439718
rect 6294 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 6914 439634
rect 6294 403954 6914 439398
rect 6294 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 6914 403954
rect 6294 403634 6914 403718
rect 6294 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 6914 403634
rect 6294 367954 6914 403398
rect 6294 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 6914 367954
rect 6294 367634 6914 367718
rect 6294 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 6914 367634
rect 6294 331954 6914 367398
rect 6294 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 6914 331954
rect 6294 331634 6914 331718
rect 6294 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 6914 331634
rect 6294 295954 6914 331398
rect 6294 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 6914 295954
rect 6294 295634 6914 295718
rect 6294 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 6914 295634
rect 6294 259954 6914 295398
rect 6294 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 6914 259954
rect 6294 259634 6914 259718
rect 6294 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 6914 259634
rect 6294 223954 6914 259398
rect 6294 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 6914 223954
rect 6294 223634 6914 223718
rect 6294 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 6914 223634
rect 6294 187954 6914 223398
rect 6294 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 6914 187954
rect 6294 187634 6914 187718
rect 6294 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 6914 187634
rect 6294 151954 6914 187398
rect 6294 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 6914 151954
rect 6294 151634 6914 151718
rect 6294 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 6914 151634
rect 6294 115954 6914 151398
rect 6294 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 6914 115954
rect 6294 115634 6914 115718
rect 6294 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 6914 115634
rect 6294 79954 6914 115398
rect 6294 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 6914 79954
rect 6294 79634 6914 79718
rect 6294 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 6914 79634
rect 6294 43954 6914 79398
rect 6294 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 6914 43954
rect 6294 43634 6914 43718
rect 6294 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 6914 43634
rect 6294 7954 6914 43398
rect 6294 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 6914 7954
rect 6294 7634 6914 7718
rect 6294 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 6914 7634
rect 6294 -1306 6914 7398
rect 6294 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 6914 -1306
rect 6294 -1626 6914 -1542
rect 6294 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 6914 -1626
rect 6294 -7654 6914 -1862
rect 10794 706758 11414 711590
rect 10794 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 11414 706758
rect 10794 706438 11414 706522
rect 10794 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 11414 706438
rect 10794 696454 11414 706202
rect 10794 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 11414 696454
rect 10794 696134 11414 696218
rect 10794 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 11414 696134
rect 10794 660454 11414 695898
rect 10794 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 11414 660454
rect 10794 660134 11414 660218
rect 10794 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 11414 660134
rect 10794 624454 11414 659898
rect 10794 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 11414 624454
rect 10794 624134 11414 624218
rect 10794 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 11414 624134
rect 10794 588454 11414 623898
rect 10794 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 11414 588454
rect 10794 588134 11414 588218
rect 10794 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 11414 588134
rect 10794 552454 11414 587898
rect 10794 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 11414 552454
rect 10794 552134 11414 552218
rect 10794 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 11414 552134
rect 10794 516454 11414 551898
rect 10794 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 11414 516454
rect 10794 516134 11414 516218
rect 10794 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 11414 516134
rect 10794 480454 11414 515898
rect 10794 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 11414 480454
rect 10794 480134 11414 480218
rect 10794 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 11414 480134
rect 10794 444454 11414 479898
rect 10794 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 11414 444454
rect 10794 444134 11414 444218
rect 10794 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 11414 444134
rect 10794 408454 11414 443898
rect 10794 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 11414 408454
rect 10794 408134 11414 408218
rect 10794 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 11414 408134
rect 10794 372454 11414 407898
rect 10794 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 11414 372454
rect 10794 372134 11414 372218
rect 10794 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 11414 372134
rect 10794 336454 11414 371898
rect 10794 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 11414 336454
rect 10794 336134 11414 336218
rect 10794 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 11414 336134
rect 10794 300454 11414 335898
rect 10794 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 11414 300454
rect 10794 300134 11414 300218
rect 10794 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 11414 300134
rect 10794 264454 11414 299898
rect 10794 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 11414 264454
rect 10794 264134 11414 264218
rect 10794 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 11414 264134
rect 10794 228454 11414 263898
rect 10794 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 11414 228454
rect 10794 228134 11414 228218
rect 10794 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 11414 228134
rect 10794 192454 11414 227898
rect 10794 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 11414 192454
rect 10794 192134 11414 192218
rect 10794 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 11414 192134
rect 10794 156454 11414 191898
rect 10794 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 11414 156454
rect 10794 156134 11414 156218
rect 10794 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 11414 156134
rect 10794 120454 11414 155898
rect 10794 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 11414 120454
rect 10794 120134 11414 120218
rect 10794 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 11414 120134
rect 10794 84454 11414 119898
rect 10794 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 11414 84454
rect 10794 84134 11414 84218
rect 10794 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 11414 84134
rect 10794 48454 11414 83898
rect 10794 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 11414 48454
rect 10794 48134 11414 48218
rect 10794 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 11414 48134
rect 10794 12454 11414 47898
rect 10794 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 11414 12454
rect 10794 12134 11414 12218
rect 10794 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 11414 12134
rect 10794 -2266 11414 11898
rect 10794 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 11414 -2266
rect 10794 -2586 11414 -2502
rect 10794 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 11414 -2586
rect 10794 -7654 11414 -2822
rect 15294 707718 15914 711590
rect 15294 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 15914 707718
rect 15294 707398 15914 707482
rect 15294 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 15914 707398
rect 15294 700954 15914 707162
rect 15294 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 15914 700954
rect 15294 700634 15914 700718
rect 15294 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 15914 700634
rect 15294 664954 15914 700398
rect 15294 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 15914 664954
rect 15294 664634 15914 664718
rect 15294 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 15914 664634
rect 15294 628954 15914 664398
rect 15294 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 15914 628954
rect 15294 628634 15914 628718
rect 15294 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 15914 628634
rect 15294 592954 15914 628398
rect 15294 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 15914 592954
rect 15294 592634 15914 592718
rect 15294 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 15914 592634
rect 15294 556954 15914 592398
rect 15294 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 15914 556954
rect 15294 556634 15914 556718
rect 15294 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 15914 556634
rect 15294 520954 15914 556398
rect 15294 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 15914 520954
rect 15294 520634 15914 520718
rect 15294 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 15914 520634
rect 15294 484954 15914 520398
rect 15294 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 15914 484954
rect 15294 484634 15914 484718
rect 15294 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 15914 484634
rect 15294 448954 15914 484398
rect 15294 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 15914 448954
rect 15294 448634 15914 448718
rect 15294 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 15914 448634
rect 15294 412954 15914 448398
rect 15294 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 15914 412954
rect 15294 412634 15914 412718
rect 15294 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 15914 412634
rect 15294 376954 15914 412398
rect 15294 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 15914 376954
rect 15294 376634 15914 376718
rect 15294 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 15914 376634
rect 15294 340954 15914 376398
rect 15294 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 15914 340954
rect 15294 340634 15914 340718
rect 15294 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 15914 340634
rect 15294 304954 15914 340398
rect 15294 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 15914 304954
rect 15294 304634 15914 304718
rect 15294 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 15914 304634
rect 15294 268954 15914 304398
rect 15294 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 15914 268954
rect 15294 268634 15914 268718
rect 15294 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 15914 268634
rect 15294 232954 15914 268398
rect 15294 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 15914 232954
rect 15294 232634 15914 232718
rect 15294 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 15914 232634
rect 15294 196954 15914 232398
rect 15294 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 15914 196954
rect 15294 196634 15914 196718
rect 15294 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 15914 196634
rect 15294 160954 15914 196398
rect 15294 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 15914 160954
rect 15294 160634 15914 160718
rect 15294 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 15914 160634
rect 15294 124954 15914 160398
rect 15294 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 15914 124954
rect 15294 124634 15914 124718
rect 15294 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 15914 124634
rect 15294 88954 15914 124398
rect 15294 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 15914 88954
rect 15294 88634 15914 88718
rect 15294 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 15914 88634
rect 15294 52954 15914 88398
rect 15294 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 15914 52954
rect 15294 52634 15914 52718
rect 15294 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 15914 52634
rect 15294 16954 15914 52398
rect 15294 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 15914 16954
rect 15294 16634 15914 16718
rect 15294 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 15914 16634
rect 15294 -3226 15914 16398
rect 15294 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 15914 -3226
rect 15294 -3546 15914 -3462
rect 15294 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 15914 -3546
rect 15294 -7654 15914 -3782
rect 19794 708678 20414 711590
rect 19794 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 20414 708678
rect 19794 708358 20414 708442
rect 19794 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 20414 708358
rect 19794 669454 20414 708122
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -4186 20414 20898
rect 19794 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 20414 -4186
rect 19794 -4506 20414 -4422
rect 19794 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 20414 -4506
rect 19794 -7654 20414 -4742
rect 24294 709638 24914 711590
rect 24294 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 24914 709638
rect 24294 709318 24914 709402
rect 24294 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 24914 709318
rect 24294 673954 24914 709082
rect 24294 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 24914 673954
rect 24294 673634 24914 673718
rect 24294 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 24914 673634
rect 24294 637954 24914 673398
rect 24294 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 24914 637954
rect 24294 637634 24914 637718
rect 24294 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 24914 637634
rect 24294 601954 24914 637398
rect 24294 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 24914 601954
rect 24294 601634 24914 601718
rect 24294 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 24914 601634
rect 24294 565954 24914 601398
rect 24294 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 24914 565954
rect 24294 565634 24914 565718
rect 24294 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 24914 565634
rect 24294 529954 24914 565398
rect 24294 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 24914 529954
rect 24294 529634 24914 529718
rect 24294 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 24914 529634
rect 24294 493954 24914 529398
rect 24294 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 24914 493954
rect 24294 493634 24914 493718
rect 24294 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 24914 493634
rect 24294 457954 24914 493398
rect 24294 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 24914 457954
rect 24294 457634 24914 457718
rect 24294 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 24914 457634
rect 24294 421954 24914 457398
rect 24294 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 24914 421954
rect 24294 421634 24914 421718
rect 24294 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 24914 421634
rect 24294 385954 24914 421398
rect 24294 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 24914 385954
rect 24294 385634 24914 385718
rect 24294 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 24914 385634
rect 24294 349954 24914 385398
rect 24294 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 24914 349954
rect 24294 349634 24914 349718
rect 24294 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 24914 349634
rect 24294 313954 24914 349398
rect 24294 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 24914 313954
rect 24294 313634 24914 313718
rect 24294 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 24914 313634
rect 24294 277954 24914 313398
rect 24294 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 24914 277954
rect 24294 277634 24914 277718
rect 24294 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 24914 277634
rect 24294 241954 24914 277398
rect 24294 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 24914 241954
rect 24294 241634 24914 241718
rect 24294 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 24914 241634
rect 24294 205954 24914 241398
rect 24294 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 24914 205954
rect 24294 205634 24914 205718
rect 24294 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 24914 205634
rect 24294 169954 24914 205398
rect 24294 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 24914 169954
rect 24294 169634 24914 169718
rect 24294 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 24914 169634
rect 24294 133954 24914 169398
rect 24294 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 24914 133954
rect 24294 133634 24914 133718
rect 24294 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 24914 133634
rect 24294 97954 24914 133398
rect 24294 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 24914 97954
rect 24294 97634 24914 97718
rect 24294 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 24914 97634
rect 24294 61954 24914 97398
rect 24294 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 24914 61954
rect 24294 61634 24914 61718
rect 24294 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 24914 61634
rect 24294 25954 24914 61398
rect 24294 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 24914 25954
rect 24294 25634 24914 25718
rect 24294 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 24914 25634
rect 24294 -5146 24914 25398
rect 24294 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 24914 -5146
rect 24294 -5466 24914 -5382
rect 24294 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 24914 -5466
rect 24294 -7654 24914 -5702
rect 28794 710598 29414 711590
rect 28794 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 29414 710598
rect 28794 710278 29414 710362
rect 28794 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 29414 710278
rect 28794 678454 29414 710042
rect 28794 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 29414 678454
rect 28794 678134 29414 678218
rect 28794 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 29414 678134
rect 28794 642454 29414 677898
rect 28794 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 29414 642454
rect 28794 642134 29414 642218
rect 28794 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 29414 642134
rect 28794 606454 29414 641898
rect 28794 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 29414 606454
rect 28794 606134 29414 606218
rect 28794 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 29414 606134
rect 28794 570454 29414 605898
rect 28794 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 29414 570454
rect 28794 570134 29414 570218
rect 28794 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 29414 570134
rect 28794 534454 29414 569898
rect 28794 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 29414 534454
rect 28794 534134 29414 534218
rect 28794 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 29414 534134
rect 28794 498454 29414 533898
rect 28794 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 29414 498454
rect 28794 498134 29414 498218
rect 28794 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 29414 498134
rect 28794 462454 29414 497898
rect 28794 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 29414 462454
rect 28794 462134 29414 462218
rect 28794 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 29414 462134
rect 28794 426454 29414 461898
rect 28794 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 29414 426454
rect 28794 426134 29414 426218
rect 28794 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 29414 426134
rect 28794 390454 29414 425898
rect 28794 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 29414 390454
rect 28794 390134 29414 390218
rect 28794 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 29414 390134
rect 28794 354454 29414 389898
rect 28794 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 29414 354454
rect 28794 354134 29414 354218
rect 28794 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 29414 354134
rect 28794 318454 29414 353898
rect 28794 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 29414 318454
rect 28794 318134 29414 318218
rect 28794 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 29414 318134
rect 28794 282454 29414 317898
rect 28794 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 29414 282454
rect 28794 282134 29414 282218
rect 28794 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 29414 282134
rect 28794 246454 29414 281898
rect 28794 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 29414 246454
rect 28794 246134 29414 246218
rect 28794 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 29414 246134
rect 28794 210454 29414 245898
rect 28794 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 29414 210454
rect 28794 210134 29414 210218
rect 28794 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 29414 210134
rect 28794 174454 29414 209898
rect 28794 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 29414 174454
rect 28794 174134 29414 174218
rect 28794 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 29414 174134
rect 28794 138454 29414 173898
rect 28794 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 29414 138454
rect 28794 138134 29414 138218
rect 28794 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 29414 138134
rect 28794 102454 29414 137898
rect 28794 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 29414 102454
rect 28794 102134 29414 102218
rect 28794 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 29414 102134
rect 28794 66454 29414 101898
rect 28794 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 29414 66454
rect 28794 66134 29414 66218
rect 28794 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 29414 66134
rect 28794 30454 29414 65898
rect 28794 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 29414 30454
rect 28794 30134 29414 30218
rect 28794 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 29414 30134
rect 28794 -6106 29414 29898
rect 28794 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 29414 -6106
rect 28794 -6426 29414 -6342
rect 28794 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 29414 -6426
rect 28794 -7654 29414 -6662
rect 33294 711558 33914 711590
rect 33294 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 33914 711558
rect 33294 711238 33914 711322
rect 33294 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 33914 711238
rect 33294 682954 33914 711002
rect 33294 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 33914 682954
rect 33294 682634 33914 682718
rect 33294 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 33914 682634
rect 33294 646954 33914 682398
rect 33294 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 33914 646954
rect 33294 646634 33914 646718
rect 33294 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 33914 646634
rect 33294 610954 33914 646398
rect 33294 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 33914 610954
rect 33294 610634 33914 610718
rect 33294 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 33914 610634
rect 33294 574954 33914 610398
rect 33294 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 33914 574954
rect 33294 574634 33914 574718
rect 33294 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 33914 574634
rect 33294 538954 33914 574398
rect 33294 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 33914 538954
rect 33294 538634 33914 538718
rect 33294 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 33914 538634
rect 33294 502954 33914 538398
rect 33294 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 33914 502954
rect 33294 502634 33914 502718
rect 33294 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 33914 502634
rect 33294 466954 33914 502398
rect 33294 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 33914 466954
rect 33294 466634 33914 466718
rect 33294 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 33914 466634
rect 33294 430954 33914 466398
rect 33294 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 33914 430954
rect 33294 430634 33914 430718
rect 33294 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 33914 430634
rect 33294 394954 33914 430398
rect 33294 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 33914 394954
rect 33294 394634 33914 394718
rect 33294 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 33914 394634
rect 33294 358954 33914 394398
rect 33294 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 33914 358954
rect 33294 358634 33914 358718
rect 33294 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 33914 358634
rect 33294 322954 33914 358398
rect 33294 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 33914 322954
rect 33294 322634 33914 322718
rect 33294 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 33914 322634
rect 33294 286954 33914 322398
rect 33294 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 33914 286954
rect 33294 286634 33914 286718
rect 33294 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 33914 286634
rect 33294 250954 33914 286398
rect 33294 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 33914 250954
rect 33294 250634 33914 250718
rect 33294 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 33914 250634
rect 33294 214954 33914 250398
rect 33294 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 33914 214954
rect 33294 214634 33914 214718
rect 33294 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 33914 214634
rect 33294 178954 33914 214398
rect 33294 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 33914 178954
rect 33294 178634 33914 178718
rect 33294 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 33914 178634
rect 33294 142954 33914 178398
rect 33294 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 33914 142954
rect 33294 142634 33914 142718
rect 33294 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 33914 142634
rect 33294 106954 33914 142398
rect 33294 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 33914 106954
rect 33294 106634 33914 106718
rect 33294 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 33914 106634
rect 33294 70954 33914 106398
rect 33294 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 33914 70954
rect 33294 70634 33914 70718
rect 33294 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 33914 70634
rect 33294 34954 33914 70398
rect 33294 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 33914 34954
rect 33294 34634 33914 34718
rect 33294 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 33914 34634
rect 33294 -7066 33914 34398
rect 33294 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 33914 -7066
rect 33294 -7386 33914 -7302
rect 33294 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 33914 -7386
rect 33294 -7654 33914 -7622
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 42294 705798 42914 711590
rect 42294 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 42914 705798
rect 42294 705478 42914 705562
rect 42294 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 42914 705478
rect 42294 691954 42914 705242
rect 42294 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 42914 691954
rect 42294 691634 42914 691718
rect 42294 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 42914 691634
rect 42294 655954 42914 691398
rect 42294 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 42914 655954
rect 42294 655634 42914 655718
rect 42294 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 42914 655634
rect 42294 619954 42914 655398
rect 42294 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 42914 619954
rect 42294 619634 42914 619718
rect 42294 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 42914 619634
rect 42294 583954 42914 619398
rect 42294 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 42914 583954
rect 42294 583634 42914 583718
rect 42294 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 42914 583634
rect 42294 547954 42914 583398
rect 42294 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 42914 547954
rect 42294 547634 42914 547718
rect 42294 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 42914 547634
rect 42294 511954 42914 547398
rect 42294 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 42914 511954
rect 42294 511634 42914 511718
rect 42294 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 42914 511634
rect 42294 475954 42914 511398
rect 42294 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 42914 475954
rect 42294 475634 42914 475718
rect 42294 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 42914 475634
rect 42294 439954 42914 475398
rect 42294 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 42914 439954
rect 42294 439634 42914 439718
rect 42294 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 42914 439634
rect 42294 403954 42914 439398
rect 42294 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 42914 403954
rect 42294 403634 42914 403718
rect 42294 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 42914 403634
rect 42294 367954 42914 403398
rect 42294 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 42914 367954
rect 42294 367634 42914 367718
rect 42294 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 42914 367634
rect 42294 331954 42914 367398
rect 42294 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 42914 331954
rect 42294 331634 42914 331718
rect 42294 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 42914 331634
rect 42294 295954 42914 331398
rect 42294 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 42914 295954
rect 42294 295634 42914 295718
rect 42294 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 42914 295634
rect 42294 259954 42914 295398
rect 42294 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 42914 259954
rect 42294 259634 42914 259718
rect 42294 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 42914 259634
rect 42294 223954 42914 259398
rect 42294 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 42914 223954
rect 42294 223634 42914 223718
rect 42294 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 42914 223634
rect 42294 187954 42914 223398
rect 42294 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 42914 187954
rect 42294 187634 42914 187718
rect 42294 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 42914 187634
rect 42294 151954 42914 187398
rect 42294 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 42914 151954
rect 42294 151634 42914 151718
rect 42294 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 42914 151634
rect 42294 115954 42914 151398
rect 42294 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 42914 115954
rect 42294 115634 42914 115718
rect 42294 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 42914 115634
rect 42294 79954 42914 115398
rect 42294 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 42914 79954
rect 42294 79634 42914 79718
rect 42294 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 42914 79634
rect 42294 43954 42914 79398
rect 42294 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 42914 43954
rect 42294 43634 42914 43718
rect 42294 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 42914 43634
rect 42294 7954 42914 43398
rect 42294 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 42914 7954
rect 42294 7634 42914 7718
rect 42294 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 42914 7634
rect 42294 -1306 42914 7398
rect 42294 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 42914 -1306
rect 42294 -1626 42914 -1542
rect 42294 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 42914 -1626
rect 42294 -7654 42914 -1862
rect 46794 706758 47414 711590
rect 46794 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 47414 706758
rect 46794 706438 47414 706522
rect 46794 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 47414 706438
rect 46794 696454 47414 706202
rect 46794 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 47414 696454
rect 46794 696134 47414 696218
rect 46794 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 47414 696134
rect 46794 660454 47414 695898
rect 46794 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 47414 660454
rect 46794 660134 47414 660218
rect 46794 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 47414 660134
rect 46794 624454 47414 659898
rect 46794 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 47414 624454
rect 46794 624134 47414 624218
rect 46794 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 47414 624134
rect 46794 588454 47414 623898
rect 46794 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 47414 588454
rect 46794 588134 47414 588218
rect 46794 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 47414 588134
rect 46794 552454 47414 587898
rect 46794 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 47414 552454
rect 46794 552134 47414 552218
rect 46794 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 47414 552134
rect 46794 516454 47414 551898
rect 46794 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 47414 516454
rect 46794 516134 47414 516218
rect 46794 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 47414 516134
rect 46794 480454 47414 515898
rect 46794 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 47414 480454
rect 46794 480134 47414 480218
rect 46794 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 47414 480134
rect 46794 444454 47414 479898
rect 46794 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 47414 444454
rect 46794 444134 47414 444218
rect 46794 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 47414 444134
rect 46794 408454 47414 443898
rect 46794 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 47414 408454
rect 46794 408134 47414 408218
rect 46794 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 47414 408134
rect 46794 372454 47414 407898
rect 46794 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 47414 372454
rect 46794 372134 47414 372218
rect 46794 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 47414 372134
rect 46794 336454 47414 371898
rect 46794 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 47414 336454
rect 46794 336134 47414 336218
rect 46794 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 47414 336134
rect 46794 300454 47414 335898
rect 46794 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 47414 300454
rect 46794 300134 47414 300218
rect 46794 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 47414 300134
rect 46794 264454 47414 299898
rect 46794 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 47414 264454
rect 46794 264134 47414 264218
rect 46794 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 47414 264134
rect 46794 228454 47414 263898
rect 46794 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 47414 228454
rect 46794 228134 47414 228218
rect 46794 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 47414 228134
rect 46794 192454 47414 227898
rect 46794 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 47414 192454
rect 46794 192134 47414 192218
rect 46794 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 47414 192134
rect 46794 156454 47414 191898
rect 46794 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 47414 156454
rect 46794 156134 47414 156218
rect 46794 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 47414 156134
rect 46794 120454 47414 155898
rect 46794 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 47414 120454
rect 46794 120134 47414 120218
rect 46794 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 47414 120134
rect 46794 84454 47414 119898
rect 46794 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 47414 84454
rect 46794 84134 47414 84218
rect 46794 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 47414 84134
rect 46794 48454 47414 83898
rect 46794 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 47414 48454
rect 46794 48134 47414 48218
rect 46794 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 47414 48134
rect 46794 12454 47414 47898
rect 46794 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 47414 12454
rect 46794 12134 47414 12218
rect 46794 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 47414 12134
rect 46794 -2266 47414 11898
rect 46794 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 47414 -2266
rect 46794 -2586 47414 -2502
rect 46794 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 47414 -2586
rect 46794 -7654 47414 -2822
rect 51294 707718 51914 711590
rect 51294 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 51914 707718
rect 51294 707398 51914 707482
rect 51294 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 51914 707398
rect 51294 700954 51914 707162
rect 51294 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 51914 700954
rect 51294 700634 51914 700718
rect 51294 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 51914 700634
rect 51294 664954 51914 700398
rect 51294 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 51914 664954
rect 51294 664634 51914 664718
rect 51294 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 51914 664634
rect 51294 628954 51914 664398
rect 51294 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 51914 628954
rect 51294 628634 51914 628718
rect 51294 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 51914 628634
rect 51294 592954 51914 628398
rect 51294 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 51914 592954
rect 51294 592634 51914 592718
rect 51294 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 51914 592634
rect 51294 556954 51914 592398
rect 51294 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 51914 556954
rect 51294 556634 51914 556718
rect 51294 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 51914 556634
rect 51294 520954 51914 556398
rect 51294 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 51914 520954
rect 51294 520634 51914 520718
rect 51294 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 51914 520634
rect 51294 484954 51914 520398
rect 51294 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 51914 484954
rect 51294 484634 51914 484718
rect 51294 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 51914 484634
rect 51294 448954 51914 484398
rect 51294 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 51914 448954
rect 51294 448634 51914 448718
rect 51294 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 51914 448634
rect 51294 412954 51914 448398
rect 51294 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 51914 412954
rect 51294 412634 51914 412718
rect 51294 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 51914 412634
rect 51294 376954 51914 412398
rect 51294 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 51914 376954
rect 51294 376634 51914 376718
rect 51294 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 51914 376634
rect 51294 340954 51914 376398
rect 51294 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 51914 340954
rect 51294 340634 51914 340718
rect 51294 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 51914 340634
rect 51294 304954 51914 340398
rect 51294 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 51914 304954
rect 51294 304634 51914 304718
rect 51294 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 51914 304634
rect 51294 268954 51914 304398
rect 51294 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 51914 268954
rect 51294 268634 51914 268718
rect 51294 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 51914 268634
rect 51294 232954 51914 268398
rect 51294 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 51914 232954
rect 51294 232634 51914 232718
rect 51294 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 51914 232634
rect 51294 196954 51914 232398
rect 51294 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 51914 196954
rect 51294 196634 51914 196718
rect 51294 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 51914 196634
rect 51294 160954 51914 196398
rect 51294 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 51914 160954
rect 51294 160634 51914 160718
rect 51294 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 51914 160634
rect 51294 124954 51914 160398
rect 51294 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 51914 124954
rect 51294 124634 51914 124718
rect 51294 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 51914 124634
rect 51294 88954 51914 124398
rect 51294 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 51914 88954
rect 51294 88634 51914 88718
rect 51294 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 51914 88634
rect 51294 52954 51914 88398
rect 51294 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 51914 52954
rect 51294 52634 51914 52718
rect 51294 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 51914 52634
rect 51294 16954 51914 52398
rect 51294 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 51914 16954
rect 51294 16634 51914 16718
rect 51294 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 51914 16634
rect 51294 -3226 51914 16398
rect 51294 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 51914 -3226
rect 51294 -3546 51914 -3462
rect 51294 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 51914 -3546
rect 51294 -7654 51914 -3782
rect 55794 708678 56414 711590
rect 55794 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 56414 708678
rect 55794 708358 56414 708442
rect 55794 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 56414 708358
rect 55794 669454 56414 708122
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -4186 56414 20898
rect 55794 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 56414 -4186
rect 55794 -4506 56414 -4422
rect 55794 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 56414 -4506
rect 55794 -7654 56414 -4742
rect 60294 709638 60914 711590
rect 60294 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 60914 709638
rect 60294 709318 60914 709402
rect 60294 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 60914 709318
rect 60294 673954 60914 709082
rect 60294 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 60914 673954
rect 60294 673634 60914 673718
rect 60294 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 60914 673634
rect 60294 637954 60914 673398
rect 60294 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 60914 637954
rect 60294 637634 60914 637718
rect 60294 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 60914 637634
rect 60294 601954 60914 637398
rect 60294 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 60914 601954
rect 60294 601634 60914 601718
rect 60294 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 60914 601634
rect 60294 565954 60914 601398
rect 60294 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 60914 565954
rect 60294 565634 60914 565718
rect 60294 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 60914 565634
rect 60294 529954 60914 565398
rect 60294 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 60914 529954
rect 60294 529634 60914 529718
rect 60294 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 60914 529634
rect 60294 493954 60914 529398
rect 60294 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 60914 493954
rect 60294 493634 60914 493718
rect 60294 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 60914 493634
rect 60294 457954 60914 493398
rect 60294 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 60914 457954
rect 60294 457634 60914 457718
rect 60294 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 60914 457634
rect 60294 421954 60914 457398
rect 60294 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 60914 421954
rect 60294 421634 60914 421718
rect 60294 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 60914 421634
rect 60294 385954 60914 421398
rect 60294 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 60914 385954
rect 60294 385634 60914 385718
rect 60294 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 60914 385634
rect 60294 349954 60914 385398
rect 60294 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 60914 349954
rect 60294 349634 60914 349718
rect 60294 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 60914 349634
rect 60294 313954 60914 349398
rect 60294 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 60914 313954
rect 60294 313634 60914 313718
rect 60294 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 60914 313634
rect 60294 277954 60914 313398
rect 60294 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 60914 277954
rect 60294 277634 60914 277718
rect 60294 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 60914 277634
rect 60294 241954 60914 277398
rect 60294 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 60914 241954
rect 60294 241634 60914 241718
rect 60294 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 60914 241634
rect 60294 205954 60914 241398
rect 60294 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 60914 205954
rect 60294 205634 60914 205718
rect 60294 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 60914 205634
rect 60294 169954 60914 205398
rect 60294 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 60914 169954
rect 60294 169634 60914 169718
rect 60294 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 60914 169634
rect 60294 133954 60914 169398
rect 60294 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 60914 133954
rect 60294 133634 60914 133718
rect 60294 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 60914 133634
rect 60294 97954 60914 133398
rect 60294 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 60914 97954
rect 60294 97634 60914 97718
rect 60294 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 60914 97634
rect 60294 61954 60914 97398
rect 60294 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 60914 61954
rect 60294 61634 60914 61718
rect 60294 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 60914 61634
rect 60294 25954 60914 61398
rect 60294 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 60914 25954
rect 60294 25634 60914 25718
rect 60294 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 60914 25634
rect 60294 -5146 60914 25398
rect 60294 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 60914 -5146
rect 60294 -5466 60914 -5382
rect 60294 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 60914 -5466
rect 60294 -7654 60914 -5702
rect 64794 710598 65414 711590
rect 64794 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 65414 710598
rect 64794 710278 65414 710362
rect 64794 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 65414 710278
rect 64794 678454 65414 710042
rect 64794 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 65414 678454
rect 64794 678134 65414 678218
rect 64794 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 65414 678134
rect 64794 642454 65414 677898
rect 64794 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 65414 642454
rect 64794 642134 65414 642218
rect 64794 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 65414 642134
rect 64794 606454 65414 641898
rect 64794 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 65414 606454
rect 64794 606134 65414 606218
rect 64794 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 65414 606134
rect 64794 570454 65414 605898
rect 64794 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 65414 570454
rect 64794 570134 65414 570218
rect 64794 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 65414 570134
rect 64794 534454 65414 569898
rect 64794 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 65414 534454
rect 64794 534134 65414 534218
rect 64794 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 65414 534134
rect 64794 498454 65414 533898
rect 64794 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 65414 498454
rect 64794 498134 65414 498218
rect 64794 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 65414 498134
rect 64794 462454 65414 497898
rect 64794 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 65414 462454
rect 64794 462134 65414 462218
rect 64794 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 65414 462134
rect 64794 426454 65414 461898
rect 64794 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 65414 426454
rect 64794 426134 65414 426218
rect 64794 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 65414 426134
rect 64794 390454 65414 425898
rect 64794 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 65414 390454
rect 64794 390134 65414 390218
rect 64794 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 65414 390134
rect 64794 354454 65414 389898
rect 64794 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 65414 354454
rect 64794 354134 65414 354218
rect 64794 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 65414 354134
rect 64794 318454 65414 353898
rect 64794 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 65414 318454
rect 64794 318134 65414 318218
rect 64794 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 65414 318134
rect 64794 282454 65414 317898
rect 64794 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 65414 282454
rect 64794 282134 65414 282218
rect 64794 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 65414 282134
rect 64794 246454 65414 281898
rect 64794 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 65414 246454
rect 64794 246134 65414 246218
rect 64794 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 65414 246134
rect 64794 210454 65414 245898
rect 64794 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 65414 210454
rect 64794 210134 65414 210218
rect 64794 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 65414 210134
rect 64794 174454 65414 209898
rect 64794 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 65414 174454
rect 64794 174134 65414 174218
rect 64794 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 65414 174134
rect 64794 138454 65414 173898
rect 64794 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 65414 138454
rect 64794 138134 65414 138218
rect 64794 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 65414 138134
rect 64794 102454 65414 137898
rect 64794 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 65414 102454
rect 64794 102134 65414 102218
rect 64794 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 65414 102134
rect 64794 66454 65414 101898
rect 64794 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 65414 66454
rect 64794 66134 65414 66218
rect 64794 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 65414 66134
rect 64794 30454 65414 65898
rect 64794 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 65414 30454
rect 64794 30134 65414 30218
rect 64794 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 65414 30134
rect 64794 -6106 65414 29898
rect 64794 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 65414 -6106
rect 64794 -6426 65414 -6342
rect 64794 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 65414 -6426
rect 64794 -7654 65414 -6662
rect 69294 711558 69914 711590
rect 69294 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 69914 711558
rect 69294 711238 69914 711322
rect 69294 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 69914 711238
rect 69294 682954 69914 711002
rect 69294 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 69914 682954
rect 69294 682634 69914 682718
rect 69294 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 69914 682634
rect 69294 646954 69914 682398
rect 69294 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 69914 646954
rect 69294 646634 69914 646718
rect 69294 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 69914 646634
rect 69294 610954 69914 646398
rect 69294 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 69914 610954
rect 69294 610634 69914 610718
rect 69294 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 69914 610634
rect 69294 574954 69914 610398
rect 69294 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 69914 574954
rect 69294 574634 69914 574718
rect 69294 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 69914 574634
rect 69294 538954 69914 574398
rect 69294 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 69914 538954
rect 69294 538634 69914 538718
rect 69294 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 69914 538634
rect 69294 502954 69914 538398
rect 69294 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 69914 502954
rect 69294 502634 69914 502718
rect 69294 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 69914 502634
rect 69294 466954 69914 502398
rect 69294 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 69914 466954
rect 69294 466634 69914 466718
rect 69294 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 69914 466634
rect 69294 430954 69914 466398
rect 69294 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 69914 430954
rect 69294 430634 69914 430718
rect 69294 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 69914 430634
rect 69294 394954 69914 430398
rect 69294 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 69914 394954
rect 69294 394634 69914 394718
rect 69294 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 69914 394634
rect 69294 358954 69914 394398
rect 69294 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 69914 358954
rect 69294 358634 69914 358718
rect 69294 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 69914 358634
rect 69294 322954 69914 358398
rect 69294 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 69914 322954
rect 69294 322634 69914 322718
rect 69294 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 69914 322634
rect 69294 286954 69914 322398
rect 69294 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 69914 286954
rect 69294 286634 69914 286718
rect 69294 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 69914 286634
rect 69294 250954 69914 286398
rect 69294 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 69914 250954
rect 69294 250634 69914 250718
rect 69294 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 69914 250634
rect 69294 214954 69914 250398
rect 69294 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 69914 214954
rect 69294 214634 69914 214718
rect 69294 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 69914 214634
rect 69294 178954 69914 214398
rect 69294 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 69914 178954
rect 69294 178634 69914 178718
rect 69294 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 69914 178634
rect 69294 142954 69914 178398
rect 69294 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 69914 142954
rect 69294 142634 69914 142718
rect 69294 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 69914 142634
rect 69294 106954 69914 142398
rect 69294 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 69914 106954
rect 69294 106634 69914 106718
rect 69294 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 69914 106634
rect 69294 70954 69914 106398
rect 69294 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 69914 70954
rect 69294 70634 69914 70718
rect 69294 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 69914 70634
rect 69294 34954 69914 70398
rect 69294 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 69914 34954
rect 69294 34634 69914 34718
rect 69294 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 69914 34634
rect 69294 -7066 69914 34398
rect 69294 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 69914 -7066
rect 69294 -7386 69914 -7302
rect 69294 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 69914 -7386
rect 69294 -7654 69914 -7622
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 78294 705798 78914 711590
rect 78294 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 78914 705798
rect 78294 705478 78914 705562
rect 78294 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 78914 705478
rect 78294 691954 78914 705242
rect 78294 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 78914 691954
rect 78294 691634 78914 691718
rect 78294 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 78914 691634
rect 78294 655954 78914 691398
rect 78294 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 78914 655954
rect 78294 655634 78914 655718
rect 78294 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 78914 655634
rect 78294 619954 78914 655398
rect 78294 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 78914 619954
rect 78294 619634 78914 619718
rect 78294 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 78914 619634
rect 78294 583954 78914 619398
rect 78294 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 78914 583954
rect 78294 583634 78914 583718
rect 78294 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 78914 583634
rect 78294 547954 78914 583398
rect 78294 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 78914 547954
rect 78294 547634 78914 547718
rect 78294 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 78914 547634
rect 78294 511954 78914 547398
rect 78294 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 78914 511954
rect 78294 511634 78914 511718
rect 78294 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 78914 511634
rect 78294 475954 78914 511398
rect 78294 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 78914 475954
rect 78294 475634 78914 475718
rect 78294 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 78914 475634
rect 78294 439954 78914 475398
rect 78294 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 78914 439954
rect 78294 439634 78914 439718
rect 78294 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 78914 439634
rect 78294 403954 78914 439398
rect 78294 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 78914 403954
rect 78294 403634 78914 403718
rect 78294 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 78914 403634
rect 78294 367954 78914 403398
rect 78294 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 78914 367954
rect 78294 367634 78914 367718
rect 78294 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 78914 367634
rect 78294 331954 78914 367398
rect 78294 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 78914 331954
rect 78294 331634 78914 331718
rect 78294 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 78914 331634
rect 78294 295954 78914 331398
rect 78294 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 78914 295954
rect 78294 295634 78914 295718
rect 78294 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 78914 295634
rect 78294 259954 78914 295398
rect 78294 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 78914 259954
rect 78294 259634 78914 259718
rect 78294 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 78914 259634
rect 78294 223954 78914 259398
rect 78294 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 78914 223954
rect 78294 223634 78914 223718
rect 78294 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 78914 223634
rect 78294 187954 78914 223398
rect 78294 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 78914 187954
rect 78294 187634 78914 187718
rect 78294 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 78914 187634
rect 78294 151954 78914 187398
rect 78294 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 78914 151954
rect 78294 151634 78914 151718
rect 78294 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 78914 151634
rect 78294 115954 78914 151398
rect 78294 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 78914 115954
rect 78294 115634 78914 115718
rect 78294 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 78914 115634
rect 78294 79954 78914 115398
rect 78294 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 78914 79954
rect 78294 79634 78914 79718
rect 78294 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 78914 79634
rect 78294 43954 78914 79398
rect 78294 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 78914 43954
rect 78294 43634 78914 43718
rect 78294 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 78914 43634
rect 78294 7954 78914 43398
rect 78294 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 78914 7954
rect 78294 7634 78914 7718
rect 78294 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 78914 7634
rect 78294 -1306 78914 7398
rect 78294 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 78914 -1306
rect 78294 -1626 78914 -1542
rect 78294 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 78914 -1626
rect 78294 -7654 78914 -1862
rect 82794 706758 83414 711590
rect 82794 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 83414 706758
rect 82794 706438 83414 706522
rect 82794 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 83414 706438
rect 82794 696454 83414 706202
rect 82794 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 83414 696454
rect 82794 696134 83414 696218
rect 82794 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 83414 696134
rect 82794 660454 83414 695898
rect 82794 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 83414 660454
rect 82794 660134 83414 660218
rect 82794 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 83414 660134
rect 82794 624454 83414 659898
rect 82794 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 83414 624454
rect 82794 624134 83414 624218
rect 82794 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 83414 624134
rect 82794 588454 83414 623898
rect 82794 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 83414 588454
rect 82794 588134 83414 588218
rect 82794 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 83414 588134
rect 82794 552454 83414 587898
rect 82794 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 83414 552454
rect 82794 552134 83414 552218
rect 82794 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 83414 552134
rect 82794 516454 83414 551898
rect 82794 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 83414 516454
rect 82794 516134 83414 516218
rect 82794 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 83414 516134
rect 82794 480454 83414 515898
rect 82794 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 83414 480454
rect 82794 480134 83414 480218
rect 82794 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 83414 480134
rect 82794 444454 83414 479898
rect 82794 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 83414 444454
rect 82794 444134 83414 444218
rect 82794 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 83414 444134
rect 82794 408454 83414 443898
rect 82794 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 83414 408454
rect 82794 408134 83414 408218
rect 82794 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 83414 408134
rect 82794 372454 83414 407898
rect 82794 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 83414 372454
rect 82794 372134 83414 372218
rect 82794 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 83414 372134
rect 82794 336454 83414 371898
rect 82794 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 83414 336454
rect 82794 336134 83414 336218
rect 82794 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 83414 336134
rect 82794 300454 83414 335898
rect 82794 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 83414 300454
rect 82794 300134 83414 300218
rect 82794 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 83414 300134
rect 82794 264454 83414 299898
rect 82794 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 83414 264454
rect 82794 264134 83414 264218
rect 82794 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 83414 264134
rect 82794 228454 83414 263898
rect 82794 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 83414 228454
rect 82794 228134 83414 228218
rect 82794 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 83414 228134
rect 82794 192454 83414 227898
rect 82794 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 83414 192454
rect 82794 192134 83414 192218
rect 82794 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 83414 192134
rect 82794 156454 83414 191898
rect 82794 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 83414 156454
rect 82794 156134 83414 156218
rect 82794 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 83414 156134
rect 82794 120454 83414 155898
rect 82794 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 83414 120454
rect 82794 120134 83414 120218
rect 82794 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 83414 120134
rect 82794 84454 83414 119898
rect 82794 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 83414 84454
rect 82794 84134 83414 84218
rect 82794 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 83414 84134
rect 82794 48454 83414 83898
rect 82794 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 83414 48454
rect 82794 48134 83414 48218
rect 82794 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 83414 48134
rect 82794 12454 83414 47898
rect 82794 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 83414 12454
rect 82794 12134 83414 12218
rect 82794 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 83414 12134
rect 82794 -2266 83414 11898
rect 82794 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 83414 -2266
rect 82794 -2586 83414 -2502
rect 82794 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 83414 -2586
rect 82794 -7654 83414 -2822
rect 87294 707718 87914 711590
rect 87294 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 87914 707718
rect 87294 707398 87914 707482
rect 87294 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 87914 707398
rect 87294 700954 87914 707162
rect 87294 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 87914 700954
rect 87294 700634 87914 700718
rect 87294 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 87914 700634
rect 87294 664954 87914 700398
rect 87294 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 87914 664954
rect 87294 664634 87914 664718
rect 87294 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 87914 664634
rect 87294 628954 87914 664398
rect 87294 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 87914 628954
rect 87294 628634 87914 628718
rect 87294 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 87914 628634
rect 87294 592954 87914 628398
rect 87294 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 87914 592954
rect 87294 592634 87914 592718
rect 87294 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 87914 592634
rect 87294 556954 87914 592398
rect 87294 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 87914 556954
rect 87294 556634 87914 556718
rect 87294 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 87914 556634
rect 87294 520954 87914 556398
rect 87294 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 87914 520954
rect 87294 520634 87914 520718
rect 87294 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 87914 520634
rect 87294 484954 87914 520398
rect 87294 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 87914 484954
rect 87294 484634 87914 484718
rect 87294 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 87914 484634
rect 87294 448954 87914 484398
rect 87294 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 87914 448954
rect 87294 448634 87914 448718
rect 87294 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 87914 448634
rect 87294 412954 87914 448398
rect 87294 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 87914 412954
rect 87294 412634 87914 412718
rect 87294 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 87914 412634
rect 87294 376954 87914 412398
rect 87294 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 87914 376954
rect 87294 376634 87914 376718
rect 87294 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 87914 376634
rect 87294 340954 87914 376398
rect 87294 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 87914 340954
rect 87294 340634 87914 340718
rect 87294 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 87914 340634
rect 87294 304954 87914 340398
rect 87294 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 87914 304954
rect 87294 304634 87914 304718
rect 87294 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 87914 304634
rect 87294 268954 87914 304398
rect 87294 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 87914 268954
rect 87294 268634 87914 268718
rect 87294 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 87914 268634
rect 87294 232954 87914 268398
rect 87294 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 87914 232954
rect 87294 232634 87914 232718
rect 87294 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 87914 232634
rect 87294 196954 87914 232398
rect 87294 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 87914 196954
rect 87294 196634 87914 196718
rect 87294 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 87914 196634
rect 87294 160954 87914 196398
rect 87294 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 87914 160954
rect 87294 160634 87914 160718
rect 87294 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 87914 160634
rect 87294 124954 87914 160398
rect 87294 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 87914 124954
rect 87294 124634 87914 124718
rect 87294 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 87914 124634
rect 87294 88954 87914 124398
rect 87294 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 87914 88954
rect 87294 88634 87914 88718
rect 87294 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 87914 88634
rect 87294 52954 87914 88398
rect 87294 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 87914 52954
rect 87294 52634 87914 52718
rect 87294 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 87914 52634
rect 87294 16954 87914 52398
rect 87294 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 87914 16954
rect 87294 16634 87914 16718
rect 87294 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 87914 16634
rect 87294 -3226 87914 16398
rect 87294 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 87914 -3226
rect 87294 -3546 87914 -3462
rect 87294 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 87914 -3546
rect 87294 -7654 87914 -3782
rect 91794 708678 92414 711590
rect 91794 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 92414 708678
rect 91794 708358 92414 708442
rect 91794 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 92414 708358
rect 91794 669454 92414 708122
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 273454 92414 308898
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 237454 92414 272898
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 129454 92414 164898
rect 91794 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 92414 129454
rect 91794 129134 92414 129218
rect 91794 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 92414 129134
rect 91794 93454 92414 128898
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 91794 57454 92414 92898
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -4186 92414 20898
rect 91794 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 92414 -4186
rect 91794 -4506 92414 -4422
rect 91794 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 92414 -4506
rect 91794 -7654 92414 -4742
rect 96294 709638 96914 711590
rect 96294 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 96914 709638
rect 96294 709318 96914 709402
rect 96294 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 96914 709318
rect 96294 673954 96914 709082
rect 96294 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 96914 673954
rect 96294 673634 96914 673718
rect 96294 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 96914 673634
rect 96294 637954 96914 673398
rect 96294 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 96914 637954
rect 96294 637634 96914 637718
rect 96294 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 96914 637634
rect 96294 601954 96914 637398
rect 96294 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 96914 601954
rect 96294 601634 96914 601718
rect 96294 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 96914 601634
rect 96294 565954 96914 601398
rect 96294 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 96914 565954
rect 96294 565634 96914 565718
rect 96294 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 96914 565634
rect 96294 529954 96914 565398
rect 96294 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 96914 529954
rect 96294 529634 96914 529718
rect 96294 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 96914 529634
rect 96294 493954 96914 529398
rect 96294 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 96914 493954
rect 96294 493634 96914 493718
rect 96294 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 96914 493634
rect 96294 457954 96914 493398
rect 96294 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 96914 457954
rect 96294 457634 96914 457718
rect 96294 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 96914 457634
rect 96294 421954 96914 457398
rect 96294 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 96914 421954
rect 96294 421634 96914 421718
rect 96294 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 96914 421634
rect 96294 385954 96914 421398
rect 96294 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 96914 385954
rect 96294 385634 96914 385718
rect 96294 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 96914 385634
rect 96294 349954 96914 385398
rect 96294 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 96914 349954
rect 96294 349634 96914 349718
rect 96294 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 96914 349634
rect 96294 313954 96914 349398
rect 96294 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 96914 313954
rect 96294 313634 96914 313718
rect 96294 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 96914 313634
rect 96294 277954 96914 313398
rect 96294 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 96914 277954
rect 96294 277634 96914 277718
rect 96294 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 96914 277634
rect 96294 241954 96914 277398
rect 96294 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 96914 241954
rect 96294 241634 96914 241718
rect 96294 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 96914 241634
rect 96294 205954 96914 241398
rect 96294 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 96914 205954
rect 96294 205634 96914 205718
rect 96294 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 96914 205634
rect 96294 169954 96914 205398
rect 96294 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 96914 169954
rect 96294 169634 96914 169718
rect 96294 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 96914 169634
rect 96294 133954 96914 169398
rect 96294 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 96914 133954
rect 96294 133634 96914 133718
rect 96294 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 96914 133634
rect 96294 97954 96914 133398
rect 96294 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 96914 97954
rect 96294 97634 96914 97718
rect 96294 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 96914 97634
rect 96294 61954 96914 97398
rect 96294 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 96914 61954
rect 96294 61634 96914 61718
rect 96294 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 96914 61634
rect 96294 25954 96914 61398
rect 96294 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 96914 25954
rect 96294 25634 96914 25718
rect 96294 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 96914 25634
rect 96294 -5146 96914 25398
rect 96294 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 96914 -5146
rect 96294 -5466 96914 -5382
rect 96294 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 96914 -5466
rect 96294 -7654 96914 -5702
rect 100794 710598 101414 711590
rect 100794 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 101414 710598
rect 100794 710278 101414 710362
rect 100794 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 101414 710278
rect 100794 678454 101414 710042
rect 100794 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 101414 678454
rect 100794 678134 101414 678218
rect 100794 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 101414 678134
rect 100794 642454 101414 677898
rect 100794 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 101414 642454
rect 100794 642134 101414 642218
rect 100794 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 101414 642134
rect 100794 606454 101414 641898
rect 100794 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 101414 606454
rect 100794 606134 101414 606218
rect 100794 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 101414 606134
rect 100794 570454 101414 605898
rect 100794 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 101414 570454
rect 100794 570134 101414 570218
rect 100794 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 101414 570134
rect 100794 534454 101414 569898
rect 100794 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 101414 534454
rect 100794 534134 101414 534218
rect 100794 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 101414 534134
rect 100794 498454 101414 533898
rect 100794 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 101414 498454
rect 100794 498134 101414 498218
rect 100794 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 101414 498134
rect 100794 462454 101414 497898
rect 100794 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 101414 462454
rect 100794 462134 101414 462218
rect 100794 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 101414 462134
rect 100794 426454 101414 461898
rect 100794 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 101414 426454
rect 100794 426134 101414 426218
rect 100794 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 101414 426134
rect 100794 390454 101414 425898
rect 100794 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 101414 390454
rect 100794 390134 101414 390218
rect 100794 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 101414 390134
rect 100794 354454 101414 389898
rect 100794 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 101414 354454
rect 100794 354134 101414 354218
rect 100794 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 101414 354134
rect 100794 318454 101414 353898
rect 100794 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 101414 318454
rect 100794 318134 101414 318218
rect 100794 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 101414 318134
rect 100794 282454 101414 317898
rect 100794 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 101414 282454
rect 100794 282134 101414 282218
rect 100794 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 101414 282134
rect 100794 246454 101414 281898
rect 100794 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 101414 246454
rect 100794 246134 101414 246218
rect 100794 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 101414 246134
rect 100794 210454 101414 245898
rect 100794 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 101414 210454
rect 100794 210134 101414 210218
rect 100794 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 101414 210134
rect 100794 174454 101414 209898
rect 100794 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 101414 174454
rect 100794 174134 101414 174218
rect 100794 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 101414 174134
rect 100794 138454 101414 173898
rect 100794 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 101414 138454
rect 100794 138134 101414 138218
rect 100794 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 101414 138134
rect 100794 102454 101414 137898
rect 100794 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 101414 102454
rect 100794 102134 101414 102218
rect 100794 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 101414 102134
rect 100794 66454 101414 101898
rect 100794 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 101414 66454
rect 100794 66134 101414 66218
rect 100794 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 101414 66134
rect 100794 30454 101414 65898
rect 100794 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 101414 30454
rect 100794 30134 101414 30218
rect 100794 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 101414 30134
rect 100794 -6106 101414 29898
rect 100794 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 101414 -6106
rect 100794 -6426 101414 -6342
rect 100794 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 101414 -6426
rect 100794 -7654 101414 -6662
rect 105294 711558 105914 711590
rect 105294 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 105914 711558
rect 105294 711238 105914 711322
rect 105294 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 105914 711238
rect 105294 682954 105914 711002
rect 105294 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 105914 682954
rect 105294 682634 105914 682718
rect 105294 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 105914 682634
rect 105294 646954 105914 682398
rect 105294 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 105914 646954
rect 105294 646634 105914 646718
rect 105294 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 105914 646634
rect 105294 610954 105914 646398
rect 105294 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 105914 610954
rect 105294 610634 105914 610718
rect 105294 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 105914 610634
rect 105294 574954 105914 610398
rect 105294 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 105914 574954
rect 105294 574634 105914 574718
rect 105294 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 105914 574634
rect 105294 538954 105914 574398
rect 105294 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 105914 538954
rect 105294 538634 105914 538718
rect 105294 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 105914 538634
rect 105294 502954 105914 538398
rect 105294 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 105914 502954
rect 105294 502634 105914 502718
rect 105294 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 105914 502634
rect 105294 466954 105914 502398
rect 105294 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 105914 466954
rect 105294 466634 105914 466718
rect 105294 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 105914 466634
rect 105294 430954 105914 466398
rect 105294 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 105914 430954
rect 105294 430634 105914 430718
rect 105294 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 105914 430634
rect 105294 394954 105914 430398
rect 105294 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 105914 394954
rect 105294 394634 105914 394718
rect 105294 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 105914 394634
rect 105294 358954 105914 394398
rect 105294 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 105914 358954
rect 105294 358634 105914 358718
rect 105294 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 105914 358634
rect 105294 322954 105914 358398
rect 105294 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 105914 322954
rect 105294 322634 105914 322718
rect 105294 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 105914 322634
rect 105294 286954 105914 322398
rect 105294 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 105914 286954
rect 105294 286634 105914 286718
rect 105294 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 105914 286634
rect 105294 250954 105914 286398
rect 105294 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 105914 250954
rect 105294 250634 105914 250718
rect 105294 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 105914 250634
rect 105294 214954 105914 250398
rect 105294 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 105914 214954
rect 105294 214634 105914 214718
rect 105294 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 105914 214634
rect 105294 178954 105914 214398
rect 105294 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 105914 178954
rect 105294 178634 105914 178718
rect 105294 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 105914 178634
rect 105294 142954 105914 178398
rect 105294 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 105914 142954
rect 105294 142634 105914 142718
rect 105294 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 105914 142634
rect 105294 106954 105914 142398
rect 105294 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 105914 106954
rect 105294 106634 105914 106718
rect 105294 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 105914 106634
rect 105294 70954 105914 106398
rect 105294 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 105914 70954
rect 105294 70634 105914 70718
rect 105294 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 105914 70634
rect 105294 34954 105914 70398
rect 105294 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 105914 34954
rect 105294 34634 105914 34718
rect 105294 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 105914 34634
rect 105294 -7066 105914 34398
rect 105294 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 105914 -7066
rect 105294 -7386 105914 -7302
rect 105294 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 105914 -7386
rect 105294 -7654 105914 -7622
rect 109794 704838 110414 711590
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 219454 110414 254898
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 114294 705798 114914 711590
rect 114294 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 114914 705798
rect 114294 705478 114914 705562
rect 114294 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 114914 705478
rect 114294 691954 114914 705242
rect 114294 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 114914 691954
rect 114294 691634 114914 691718
rect 114294 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 114914 691634
rect 114294 655954 114914 691398
rect 114294 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 114914 655954
rect 114294 655634 114914 655718
rect 114294 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 114914 655634
rect 114294 619954 114914 655398
rect 114294 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 114914 619954
rect 114294 619634 114914 619718
rect 114294 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 114914 619634
rect 114294 583954 114914 619398
rect 114294 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 114914 583954
rect 114294 583634 114914 583718
rect 114294 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 114914 583634
rect 114294 547954 114914 583398
rect 114294 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 114914 547954
rect 114294 547634 114914 547718
rect 114294 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 114914 547634
rect 114294 511954 114914 547398
rect 114294 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 114914 511954
rect 114294 511634 114914 511718
rect 114294 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 114914 511634
rect 114294 475954 114914 511398
rect 114294 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 114914 475954
rect 114294 475634 114914 475718
rect 114294 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 114914 475634
rect 114294 439954 114914 475398
rect 114294 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 114914 439954
rect 114294 439634 114914 439718
rect 114294 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 114914 439634
rect 114294 403954 114914 439398
rect 114294 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 114914 403954
rect 114294 403634 114914 403718
rect 114294 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 114914 403634
rect 114294 367954 114914 403398
rect 114294 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 114914 367954
rect 114294 367634 114914 367718
rect 114294 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 114914 367634
rect 114294 331954 114914 367398
rect 114294 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 114914 331954
rect 114294 331634 114914 331718
rect 114294 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 114914 331634
rect 114294 295954 114914 331398
rect 114294 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 114914 295954
rect 114294 295634 114914 295718
rect 114294 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 114914 295634
rect 114294 259954 114914 295398
rect 114294 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 114914 259954
rect 114294 259634 114914 259718
rect 114294 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 114914 259634
rect 114294 223954 114914 259398
rect 114294 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 114914 223954
rect 114294 223634 114914 223718
rect 114294 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 114914 223634
rect 114294 187954 114914 223398
rect 114294 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 114914 187954
rect 114294 187634 114914 187718
rect 114294 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 114914 187634
rect 114294 151954 114914 187398
rect 114294 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 114914 151954
rect 114294 151634 114914 151718
rect 114294 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 114914 151634
rect 114294 115954 114914 151398
rect 118794 706758 119414 711590
rect 118794 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 119414 706758
rect 118794 706438 119414 706522
rect 118794 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 119414 706438
rect 118794 696454 119414 706202
rect 118794 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 119414 696454
rect 118794 696134 119414 696218
rect 118794 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 119414 696134
rect 118794 660454 119414 695898
rect 118794 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 119414 660454
rect 118794 660134 119414 660218
rect 118794 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 119414 660134
rect 118794 624454 119414 659898
rect 118794 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 119414 624454
rect 118794 624134 119414 624218
rect 118794 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 119414 624134
rect 118794 588454 119414 623898
rect 118794 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 119414 588454
rect 118794 588134 119414 588218
rect 118794 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 119414 588134
rect 118794 552454 119414 587898
rect 118794 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 119414 552454
rect 118794 552134 119414 552218
rect 118794 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 119414 552134
rect 118794 516454 119414 551898
rect 118794 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 119414 516454
rect 118794 516134 119414 516218
rect 118794 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 119414 516134
rect 118794 480454 119414 515898
rect 118794 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 119414 480454
rect 118794 480134 119414 480218
rect 118794 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 119414 480134
rect 118794 444454 119414 479898
rect 118794 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 119414 444454
rect 118794 444134 119414 444218
rect 118794 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 119414 444134
rect 118794 408454 119414 443898
rect 118794 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 119414 408454
rect 118794 408134 119414 408218
rect 118794 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 119414 408134
rect 118794 372454 119414 407898
rect 118794 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 119414 372454
rect 118794 372134 119414 372218
rect 118794 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 119414 372134
rect 118794 336454 119414 371898
rect 118794 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 119414 336454
rect 118794 336134 119414 336218
rect 118794 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 119414 336134
rect 118794 300454 119414 335898
rect 118794 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 119414 300454
rect 118794 300134 119414 300218
rect 118794 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 119414 300134
rect 118794 264454 119414 299898
rect 118794 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 119414 264454
rect 118794 264134 119414 264218
rect 118794 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 119414 264134
rect 118794 228454 119414 263898
rect 118794 228218 118826 228454
rect 119062 228218 119146 228454
rect 119382 228218 119414 228454
rect 118794 228134 119414 228218
rect 118794 227898 118826 228134
rect 119062 227898 119146 228134
rect 119382 227898 119414 228134
rect 118794 192454 119414 227898
rect 118794 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 119414 192454
rect 118794 192134 119414 192218
rect 118794 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 119414 192134
rect 118794 156454 119414 191898
rect 118794 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 119414 156454
rect 118794 156134 119414 156218
rect 118794 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 119414 156134
rect 118794 142000 119414 155898
rect 123294 707718 123914 711590
rect 123294 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 123914 707718
rect 123294 707398 123914 707482
rect 123294 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 123914 707398
rect 123294 700954 123914 707162
rect 123294 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 123914 700954
rect 123294 700634 123914 700718
rect 123294 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 123914 700634
rect 123294 664954 123914 700398
rect 123294 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 123914 664954
rect 123294 664634 123914 664718
rect 123294 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 123914 664634
rect 123294 628954 123914 664398
rect 123294 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 123914 628954
rect 123294 628634 123914 628718
rect 123294 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 123914 628634
rect 123294 592954 123914 628398
rect 123294 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 123914 592954
rect 123294 592634 123914 592718
rect 123294 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 123914 592634
rect 123294 556954 123914 592398
rect 123294 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 123914 556954
rect 123294 556634 123914 556718
rect 123294 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 123914 556634
rect 123294 520954 123914 556398
rect 123294 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 123914 520954
rect 123294 520634 123914 520718
rect 123294 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 123914 520634
rect 123294 484954 123914 520398
rect 123294 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 123914 484954
rect 123294 484634 123914 484718
rect 123294 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 123914 484634
rect 123294 448954 123914 484398
rect 123294 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 123914 448954
rect 123294 448634 123914 448718
rect 123294 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 123914 448634
rect 123294 412954 123914 448398
rect 123294 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 123914 412954
rect 123294 412634 123914 412718
rect 123294 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 123914 412634
rect 123294 376954 123914 412398
rect 123294 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 123914 376954
rect 123294 376634 123914 376718
rect 123294 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 123914 376634
rect 123294 340954 123914 376398
rect 123294 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 123914 340954
rect 123294 340634 123914 340718
rect 123294 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 123914 340634
rect 123294 304954 123914 340398
rect 123294 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 123914 304954
rect 123294 304634 123914 304718
rect 123294 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 123914 304634
rect 123294 268954 123914 304398
rect 123294 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 123914 268954
rect 123294 268634 123914 268718
rect 123294 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 123914 268634
rect 123294 232954 123914 268398
rect 123294 232718 123326 232954
rect 123562 232718 123646 232954
rect 123882 232718 123914 232954
rect 123294 232634 123914 232718
rect 123294 232398 123326 232634
rect 123562 232398 123646 232634
rect 123882 232398 123914 232634
rect 123294 196954 123914 232398
rect 123294 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 123914 196954
rect 123294 196634 123914 196718
rect 123294 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 123914 196634
rect 123294 160954 123914 196398
rect 123294 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 123914 160954
rect 123294 160634 123914 160718
rect 123294 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 123914 160634
rect 123294 142000 123914 160398
rect 127794 708678 128414 711590
rect 127794 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 128414 708678
rect 127794 708358 128414 708442
rect 127794 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 128414 708358
rect 127794 669454 128414 708122
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 201454 128414 236898
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 127794 165454 128414 200898
rect 127794 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 128414 165454
rect 127794 165134 128414 165218
rect 127794 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 128414 165134
rect 127794 142000 128414 164898
rect 132294 709638 132914 711590
rect 132294 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 132914 709638
rect 132294 709318 132914 709402
rect 132294 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 132914 709318
rect 132294 673954 132914 709082
rect 132294 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 132914 673954
rect 132294 673634 132914 673718
rect 132294 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 132914 673634
rect 132294 637954 132914 673398
rect 132294 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 132914 637954
rect 132294 637634 132914 637718
rect 132294 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 132914 637634
rect 132294 601954 132914 637398
rect 132294 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 132914 601954
rect 132294 601634 132914 601718
rect 132294 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 132914 601634
rect 132294 565954 132914 601398
rect 132294 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 132914 565954
rect 132294 565634 132914 565718
rect 132294 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 132914 565634
rect 132294 529954 132914 565398
rect 132294 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 132914 529954
rect 132294 529634 132914 529718
rect 132294 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 132914 529634
rect 132294 493954 132914 529398
rect 132294 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 132914 493954
rect 132294 493634 132914 493718
rect 132294 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 132914 493634
rect 132294 457954 132914 493398
rect 132294 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 132914 457954
rect 132294 457634 132914 457718
rect 132294 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 132914 457634
rect 132294 421954 132914 457398
rect 132294 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 132914 421954
rect 132294 421634 132914 421718
rect 132294 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 132914 421634
rect 132294 385954 132914 421398
rect 132294 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 132914 385954
rect 132294 385634 132914 385718
rect 132294 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 132914 385634
rect 132294 349954 132914 385398
rect 132294 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 132914 349954
rect 132294 349634 132914 349718
rect 132294 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 132914 349634
rect 132294 313954 132914 349398
rect 132294 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 132914 313954
rect 132294 313634 132914 313718
rect 132294 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 132914 313634
rect 132294 277954 132914 313398
rect 132294 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 132914 277954
rect 132294 277634 132914 277718
rect 132294 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 132914 277634
rect 132294 241954 132914 277398
rect 132294 241718 132326 241954
rect 132562 241718 132646 241954
rect 132882 241718 132914 241954
rect 132294 241634 132914 241718
rect 132294 241398 132326 241634
rect 132562 241398 132646 241634
rect 132882 241398 132914 241634
rect 132294 205954 132914 241398
rect 132294 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205718 132914 205954
rect 132294 205634 132914 205718
rect 132294 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205398 132914 205634
rect 132294 169954 132914 205398
rect 132294 169718 132326 169954
rect 132562 169718 132646 169954
rect 132882 169718 132914 169954
rect 132294 169634 132914 169718
rect 132294 169398 132326 169634
rect 132562 169398 132646 169634
rect 132882 169398 132914 169634
rect 132294 142000 132914 169398
rect 136794 710598 137414 711590
rect 136794 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 137414 710598
rect 136794 710278 137414 710362
rect 136794 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 137414 710278
rect 136794 678454 137414 710042
rect 136794 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 137414 678454
rect 136794 678134 137414 678218
rect 136794 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 137414 678134
rect 136794 642454 137414 677898
rect 136794 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 137414 642454
rect 136794 642134 137414 642218
rect 136794 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 137414 642134
rect 136794 606454 137414 641898
rect 136794 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 137414 606454
rect 136794 606134 137414 606218
rect 136794 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 137414 606134
rect 136794 570454 137414 605898
rect 136794 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 137414 570454
rect 136794 570134 137414 570218
rect 136794 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 137414 570134
rect 136794 534454 137414 569898
rect 136794 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 137414 534454
rect 136794 534134 137414 534218
rect 136794 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 137414 534134
rect 136794 498454 137414 533898
rect 136794 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 137414 498454
rect 136794 498134 137414 498218
rect 136794 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 137414 498134
rect 136794 462454 137414 497898
rect 136794 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 137414 462454
rect 136794 462134 137414 462218
rect 136794 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 137414 462134
rect 136794 426454 137414 461898
rect 136794 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 137414 426454
rect 136794 426134 137414 426218
rect 136794 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 137414 426134
rect 136794 390454 137414 425898
rect 136794 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 137414 390454
rect 136794 390134 137414 390218
rect 136794 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 137414 390134
rect 136794 354454 137414 389898
rect 136794 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 137414 354454
rect 136794 354134 137414 354218
rect 136794 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 137414 354134
rect 136794 318454 137414 353898
rect 136794 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 137414 318454
rect 136794 318134 137414 318218
rect 136794 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 137414 318134
rect 136794 282454 137414 317898
rect 136794 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 137414 282454
rect 136794 282134 137414 282218
rect 136794 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 137414 282134
rect 136794 246454 137414 281898
rect 136794 246218 136826 246454
rect 137062 246218 137146 246454
rect 137382 246218 137414 246454
rect 136794 246134 137414 246218
rect 136794 245898 136826 246134
rect 137062 245898 137146 246134
rect 137382 245898 137414 246134
rect 136794 210454 137414 245898
rect 136794 210218 136826 210454
rect 137062 210218 137146 210454
rect 137382 210218 137414 210454
rect 136794 210134 137414 210218
rect 136794 209898 136826 210134
rect 137062 209898 137146 210134
rect 137382 209898 137414 210134
rect 136794 174454 137414 209898
rect 136794 174218 136826 174454
rect 137062 174218 137146 174454
rect 137382 174218 137414 174454
rect 136794 174134 137414 174218
rect 136794 173898 136826 174134
rect 137062 173898 137146 174134
rect 137382 173898 137414 174134
rect 136794 142000 137414 173898
rect 141294 711558 141914 711590
rect 141294 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 141914 711558
rect 141294 711238 141914 711322
rect 141294 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 141914 711238
rect 141294 682954 141914 711002
rect 141294 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 141914 682954
rect 141294 682634 141914 682718
rect 141294 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 141914 682634
rect 141294 646954 141914 682398
rect 141294 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 141914 646954
rect 141294 646634 141914 646718
rect 141294 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 141914 646634
rect 141294 610954 141914 646398
rect 141294 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 141914 610954
rect 141294 610634 141914 610718
rect 141294 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 141914 610634
rect 141294 574954 141914 610398
rect 141294 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 141914 574954
rect 141294 574634 141914 574718
rect 141294 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 141914 574634
rect 141294 538954 141914 574398
rect 141294 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 141914 538954
rect 141294 538634 141914 538718
rect 141294 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 141914 538634
rect 141294 502954 141914 538398
rect 141294 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 141914 502954
rect 141294 502634 141914 502718
rect 141294 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 141914 502634
rect 141294 466954 141914 502398
rect 141294 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 141914 466954
rect 141294 466634 141914 466718
rect 141294 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 141914 466634
rect 141294 430954 141914 466398
rect 141294 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 141914 430954
rect 141294 430634 141914 430718
rect 141294 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 141914 430634
rect 141294 394954 141914 430398
rect 141294 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 141914 394954
rect 141294 394634 141914 394718
rect 141294 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 141914 394634
rect 141294 358954 141914 394398
rect 141294 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 141914 358954
rect 141294 358634 141914 358718
rect 141294 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 141914 358634
rect 141294 322954 141914 358398
rect 141294 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 141914 322954
rect 141294 322634 141914 322718
rect 141294 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 141914 322634
rect 141294 286954 141914 322398
rect 141294 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 141914 286954
rect 141294 286634 141914 286718
rect 141294 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 141914 286634
rect 141294 250954 141914 286398
rect 141294 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 141914 250954
rect 141294 250634 141914 250718
rect 141294 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 141914 250634
rect 141294 214954 141914 250398
rect 141294 214718 141326 214954
rect 141562 214718 141646 214954
rect 141882 214718 141914 214954
rect 141294 214634 141914 214718
rect 141294 214398 141326 214634
rect 141562 214398 141646 214634
rect 141882 214398 141914 214634
rect 141294 178954 141914 214398
rect 141294 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 141914 178954
rect 141294 178634 141914 178718
rect 141294 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 141914 178634
rect 141294 142954 141914 178398
rect 141294 142718 141326 142954
rect 141562 142718 141646 142954
rect 141882 142718 141914 142954
rect 141294 142634 141914 142718
rect 141294 142398 141326 142634
rect 141562 142398 141646 142634
rect 141882 142398 141914 142634
rect 141294 142000 141914 142398
rect 145794 704838 146414 711590
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 147454 146414 182898
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 142000 146414 146898
rect 150294 705798 150914 711590
rect 150294 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 150914 705798
rect 150294 705478 150914 705562
rect 150294 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 150914 705478
rect 150294 691954 150914 705242
rect 150294 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 150914 691954
rect 150294 691634 150914 691718
rect 150294 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 150914 691634
rect 150294 655954 150914 691398
rect 150294 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 150914 655954
rect 150294 655634 150914 655718
rect 150294 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 150914 655634
rect 150294 619954 150914 655398
rect 150294 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 150914 619954
rect 150294 619634 150914 619718
rect 150294 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 150914 619634
rect 150294 583954 150914 619398
rect 150294 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 150914 583954
rect 150294 583634 150914 583718
rect 150294 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 150914 583634
rect 150294 547954 150914 583398
rect 150294 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 150914 547954
rect 150294 547634 150914 547718
rect 150294 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 150914 547634
rect 150294 511954 150914 547398
rect 150294 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 150914 511954
rect 150294 511634 150914 511718
rect 150294 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 150914 511634
rect 150294 475954 150914 511398
rect 150294 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 150914 475954
rect 150294 475634 150914 475718
rect 150294 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 150914 475634
rect 150294 439954 150914 475398
rect 150294 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 150914 439954
rect 150294 439634 150914 439718
rect 150294 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 150914 439634
rect 150294 403954 150914 439398
rect 150294 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 150914 403954
rect 150294 403634 150914 403718
rect 150294 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 150914 403634
rect 150294 367954 150914 403398
rect 150294 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 150914 367954
rect 150294 367634 150914 367718
rect 150294 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 150914 367634
rect 150294 331954 150914 367398
rect 150294 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 150914 331954
rect 150294 331634 150914 331718
rect 150294 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 150914 331634
rect 150294 295954 150914 331398
rect 150294 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 150914 295954
rect 150294 295634 150914 295718
rect 150294 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 150914 295634
rect 150294 259954 150914 295398
rect 150294 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 150914 259954
rect 150294 259634 150914 259718
rect 150294 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 150914 259634
rect 150294 223954 150914 259398
rect 150294 223718 150326 223954
rect 150562 223718 150646 223954
rect 150882 223718 150914 223954
rect 150294 223634 150914 223718
rect 150294 223398 150326 223634
rect 150562 223398 150646 223634
rect 150882 223398 150914 223634
rect 150294 187954 150914 223398
rect 150294 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 150914 187954
rect 150294 187634 150914 187718
rect 150294 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 150914 187634
rect 150294 151954 150914 187398
rect 150294 151718 150326 151954
rect 150562 151718 150646 151954
rect 150882 151718 150914 151954
rect 150294 151634 150914 151718
rect 150294 151398 150326 151634
rect 150562 151398 150646 151634
rect 150882 151398 150914 151634
rect 150294 142000 150914 151398
rect 154794 706758 155414 711590
rect 154794 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 155414 706758
rect 154794 706438 155414 706522
rect 154794 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 155414 706438
rect 154794 696454 155414 706202
rect 154794 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 155414 696454
rect 154794 696134 155414 696218
rect 154794 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 155414 696134
rect 154794 660454 155414 695898
rect 154794 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 155414 660454
rect 154794 660134 155414 660218
rect 154794 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 155414 660134
rect 154794 624454 155414 659898
rect 154794 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 155414 624454
rect 154794 624134 155414 624218
rect 154794 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 155414 624134
rect 154794 588454 155414 623898
rect 154794 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 155414 588454
rect 154794 588134 155414 588218
rect 154794 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 155414 588134
rect 154794 552454 155414 587898
rect 154794 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 155414 552454
rect 154794 552134 155414 552218
rect 154794 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 155414 552134
rect 154794 516454 155414 551898
rect 154794 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 155414 516454
rect 154794 516134 155414 516218
rect 154794 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 155414 516134
rect 154794 480454 155414 515898
rect 154794 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 155414 480454
rect 154794 480134 155414 480218
rect 154794 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 155414 480134
rect 154794 444454 155414 479898
rect 154794 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 155414 444454
rect 154794 444134 155414 444218
rect 154794 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 155414 444134
rect 154794 408454 155414 443898
rect 154794 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 155414 408454
rect 154794 408134 155414 408218
rect 154794 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 155414 408134
rect 154794 372454 155414 407898
rect 154794 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 155414 372454
rect 154794 372134 155414 372218
rect 154794 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 155414 372134
rect 154794 336454 155414 371898
rect 154794 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 155414 336454
rect 154794 336134 155414 336218
rect 154794 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 155414 336134
rect 154794 300454 155414 335898
rect 154794 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 155414 300454
rect 154794 300134 155414 300218
rect 154794 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 155414 300134
rect 154794 264454 155414 299898
rect 154794 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 155414 264454
rect 154794 264134 155414 264218
rect 154794 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 155414 264134
rect 154794 228454 155414 263898
rect 154794 228218 154826 228454
rect 155062 228218 155146 228454
rect 155382 228218 155414 228454
rect 154794 228134 155414 228218
rect 154794 227898 154826 228134
rect 155062 227898 155146 228134
rect 155382 227898 155414 228134
rect 154794 192454 155414 227898
rect 154794 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 155414 192454
rect 154794 192134 155414 192218
rect 154794 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 155414 192134
rect 154794 156454 155414 191898
rect 154794 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 155414 156454
rect 154794 156134 155414 156218
rect 154794 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 155414 156134
rect 154794 142000 155414 155898
rect 159294 707718 159914 711590
rect 159294 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 159914 707718
rect 159294 707398 159914 707482
rect 159294 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 159914 707398
rect 159294 700954 159914 707162
rect 159294 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 159914 700954
rect 159294 700634 159914 700718
rect 159294 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 159914 700634
rect 159294 664954 159914 700398
rect 159294 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 159914 664954
rect 159294 664634 159914 664718
rect 159294 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 159914 664634
rect 159294 628954 159914 664398
rect 159294 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 159914 628954
rect 159294 628634 159914 628718
rect 159294 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 159914 628634
rect 159294 592954 159914 628398
rect 159294 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 159914 592954
rect 159294 592634 159914 592718
rect 159294 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 159914 592634
rect 159294 556954 159914 592398
rect 159294 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 159914 556954
rect 159294 556634 159914 556718
rect 159294 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 159914 556634
rect 159294 520954 159914 556398
rect 159294 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 159914 520954
rect 159294 520634 159914 520718
rect 159294 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 159914 520634
rect 159294 484954 159914 520398
rect 159294 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 159914 484954
rect 159294 484634 159914 484718
rect 159294 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 159914 484634
rect 159294 448954 159914 484398
rect 159294 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 159914 448954
rect 159294 448634 159914 448718
rect 159294 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 159914 448634
rect 159294 412954 159914 448398
rect 159294 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 159914 412954
rect 159294 412634 159914 412718
rect 159294 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 159914 412634
rect 159294 376954 159914 412398
rect 159294 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 159914 376954
rect 159294 376634 159914 376718
rect 159294 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 159914 376634
rect 159294 340954 159914 376398
rect 159294 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 159914 340954
rect 159294 340634 159914 340718
rect 159294 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 159914 340634
rect 159294 304954 159914 340398
rect 159294 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 159914 304954
rect 159294 304634 159914 304718
rect 159294 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 159914 304634
rect 159294 268954 159914 304398
rect 159294 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 159914 268954
rect 159294 268634 159914 268718
rect 159294 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 159914 268634
rect 159294 232954 159914 268398
rect 159294 232718 159326 232954
rect 159562 232718 159646 232954
rect 159882 232718 159914 232954
rect 159294 232634 159914 232718
rect 159294 232398 159326 232634
rect 159562 232398 159646 232634
rect 159882 232398 159914 232634
rect 159294 196954 159914 232398
rect 159294 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 159914 196954
rect 159294 196634 159914 196718
rect 159294 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 159914 196634
rect 159294 160954 159914 196398
rect 159294 160718 159326 160954
rect 159562 160718 159646 160954
rect 159882 160718 159914 160954
rect 159294 160634 159914 160718
rect 159294 160398 159326 160634
rect 159562 160398 159646 160634
rect 159882 160398 159914 160634
rect 159294 142000 159914 160398
rect 163794 708678 164414 711590
rect 163794 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 164414 708678
rect 163794 708358 164414 708442
rect 163794 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 164414 708358
rect 163794 669454 164414 708122
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 201454 164414 236898
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 163794 165454 164414 200898
rect 163794 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 164414 165454
rect 163794 165134 164414 165218
rect 163794 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 164414 165134
rect 163794 142000 164414 164898
rect 168294 709638 168914 711590
rect 168294 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 168914 709638
rect 168294 709318 168914 709402
rect 168294 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 168914 709318
rect 168294 673954 168914 709082
rect 168294 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 168914 673954
rect 168294 673634 168914 673718
rect 168294 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 168914 673634
rect 168294 637954 168914 673398
rect 168294 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 168914 637954
rect 168294 637634 168914 637718
rect 168294 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 168914 637634
rect 168294 601954 168914 637398
rect 168294 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 168914 601954
rect 168294 601634 168914 601718
rect 168294 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 168914 601634
rect 168294 565954 168914 601398
rect 168294 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 168914 565954
rect 168294 565634 168914 565718
rect 168294 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 168914 565634
rect 168294 529954 168914 565398
rect 168294 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 168914 529954
rect 168294 529634 168914 529718
rect 168294 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 168914 529634
rect 168294 493954 168914 529398
rect 168294 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 168914 493954
rect 168294 493634 168914 493718
rect 168294 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 168914 493634
rect 168294 457954 168914 493398
rect 168294 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 168914 457954
rect 168294 457634 168914 457718
rect 168294 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 168914 457634
rect 168294 421954 168914 457398
rect 168294 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 168914 421954
rect 168294 421634 168914 421718
rect 168294 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 168914 421634
rect 168294 385954 168914 421398
rect 168294 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 168914 385954
rect 168294 385634 168914 385718
rect 168294 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 168914 385634
rect 168294 349954 168914 385398
rect 168294 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 168914 349954
rect 168294 349634 168914 349718
rect 168294 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 168914 349634
rect 168294 313954 168914 349398
rect 168294 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 168914 313954
rect 168294 313634 168914 313718
rect 168294 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 168914 313634
rect 168294 277954 168914 313398
rect 168294 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 168914 277954
rect 168294 277634 168914 277718
rect 168294 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 168914 277634
rect 168294 241954 168914 277398
rect 168294 241718 168326 241954
rect 168562 241718 168646 241954
rect 168882 241718 168914 241954
rect 168294 241634 168914 241718
rect 168294 241398 168326 241634
rect 168562 241398 168646 241634
rect 168882 241398 168914 241634
rect 168294 205954 168914 241398
rect 168294 205718 168326 205954
rect 168562 205718 168646 205954
rect 168882 205718 168914 205954
rect 168294 205634 168914 205718
rect 168294 205398 168326 205634
rect 168562 205398 168646 205634
rect 168882 205398 168914 205634
rect 168294 169954 168914 205398
rect 168294 169718 168326 169954
rect 168562 169718 168646 169954
rect 168882 169718 168914 169954
rect 168294 169634 168914 169718
rect 168294 169398 168326 169634
rect 168562 169398 168646 169634
rect 168882 169398 168914 169634
rect 168294 142000 168914 169398
rect 172794 710598 173414 711590
rect 172794 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 173414 710598
rect 172794 710278 173414 710362
rect 172794 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 173414 710278
rect 172794 678454 173414 710042
rect 172794 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 173414 678454
rect 172794 678134 173414 678218
rect 172794 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 173414 678134
rect 172794 642454 173414 677898
rect 172794 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 173414 642454
rect 172794 642134 173414 642218
rect 172794 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 173414 642134
rect 172794 606454 173414 641898
rect 172794 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 173414 606454
rect 172794 606134 173414 606218
rect 172794 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 173414 606134
rect 172794 570454 173414 605898
rect 172794 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 173414 570454
rect 172794 570134 173414 570218
rect 172794 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 173414 570134
rect 172794 534454 173414 569898
rect 172794 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 173414 534454
rect 172794 534134 173414 534218
rect 172794 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 173414 534134
rect 172794 498454 173414 533898
rect 172794 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 173414 498454
rect 172794 498134 173414 498218
rect 172794 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 173414 498134
rect 172794 462454 173414 497898
rect 172794 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 173414 462454
rect 172794 462134 173414 462218
rect 172794 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 173414 462134
rect 172794 426454 173414 461898
rect 172794 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 173414 426454
rect 172794 426134 173414 426218
rect 172794 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 173414 426134
rect 172794 390454 173414 425898
rect 172794 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 173414 390454
rect 172794 390134 173414 390218
rect 172794 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 173414 390134
rect 172794 354454 173414 389898
rect 172794 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 173414 354454
rect 172794 354134 173414 354218
rect 172794 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 173414 354134
rect 172794 318454 173414 353898
rect 172794 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 173414 318454
rect 172794 318134 173414 318218
rect 172794 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 173414 318134
rect 172794 282454 173414 317898
rect 172794 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 173414 282454
rect 172794 282134 173414 282218
rect 172794 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 173414 282134
rect 172794 246454 173414 281898
rect 172794 246218 172826 246454
rect 173062 246218 173146 246454
rect 173382 246218 173414 246454
rect 172794 246134 173414 246218
rect 172794 245898 172826 246134
rect 173062 245898 173146 246134
rect 173382 245898 173414 246134
rect 172794 210454 173414 245898
rect 172794 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 173414 210454
rect 172794 210134 173414 210218
rect 172794 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 173414 210134
rect 172794 174454 173414 209898
rect 172794 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 173414 174454
rect 172794 174134 173414 174218
rect 172794 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 173414 174134
rect 172794 142000 173414 173898
rect 177294 711558 177914 711590
rect 177294 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 177914 711558
rect 177294 711238 177914 711322
rect 177294 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 177914 711238
rect 177294 682954 177914 711002
rect 177294 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 177914 682954
rect 177294 682634 177914 682718
rect 177294 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 177914 682634
rect 177294 646954 177914 682398
rect 177294 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 177914 646954
rect 177294 646634 177914 646718
rect 177294 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 177914 646634
rect 177294 610954 177914 646398
rect 177294 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 177914 610954
rect 177294 610634 177914 610718
rect 177294 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 177914 610634
rect 177294 574954 177914 610398
rect 177294 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 177914 574954
rect 177294 574634 177914 574718
rect 177294 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 177914 574634
rect 177294 538954 177914 574398
rect 177294 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 177914 538954
rect 177294 538634 177914 538718
rect 177294 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 177914 538634
rect 177294 502954 177914 538398
rect 177294 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 177914 502954
rect 177294 502634 177914 502718
rect 177294 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 177914 502634
rect 177294 466954 177914 502398
rect 177294 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 177914 466954
rect 177294 466634 177914 466718
rect 177294 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 177914 466634
rect 177294 430954 177914 466398
rect 177294 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 177914 430954
rect 177294 430634 177914 430718
rect 177294 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 177914 430634
rect 177294 394954 177914 430398
rect 177294 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 177914 394954
rect 177294 394634 177914 394718
rect 177294 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 177914 394634
rect 177294 358954 177914 394398
rect 177294 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 177914 358954
rect 177294 358634 177914 358718
rect 177294 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 177914 358634
rect 177294 322954 177914 358398
rect 177294 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 177914 322954
rect 177294 322634 177914 322718
rect 177294 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 177914 322634
rect 177294 286954 177914 322398
rect 177294 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 177914 286954
rect 177294 286634 177914 286718
rect 177294 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 177914 286634
rect 177294 250954 177914 286398
rect 177294 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 177914 250954
rect 177294 250634 177914 250718
rect 177294 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 177914 250634
rect 177294 214954 177914 250398
rect 177294 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 177914 214954
rect 177294 214634 177914 214718
rect 177294 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 177914 214634
rect 177294 178954 177914 214398
rect 177294 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 177914 178954
rect 177294 178634 177914 178718
rect 177294 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 177914 178634
rect 177294 142954 177914 178398
rect 177294 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 177914 142954
rect 177294 142634 177914 142718
rect 177294 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 177914 142634
rect 177294 142000 177914 142398
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 142000 182414 146898
rect 186294 705798 186914 711590
rect 186294 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 186914 705798
rect 186294 705478 186914 705562
rect 186294 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 186914 705478
rect 186294 691954 186914 705242
rect 186294 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 186914 691954
rect 186294 691634 186914 691718
rect 186294 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 186914 691634
rect 186294 655954 186914 691398
rect 186294 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 186914 655954
rect 186294 655634 186914 655718
rect 186294 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 186914 655634
rect 186294 619954 186914 655398
rect 186294 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 186914 619954
rect 186294 619634 186914 619718
rect 186294 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 186914 619634
rect 186294 583954 186914 619398
rect 186294 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 186914 583954
rect 186294 583634 186914 583718
rect 186294 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 186914 583634
rect 186294 547954 186914 583398
rect 186294 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 186914 547954
rect 186294 547634 186914 547718
rect 186294 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 186914 547634
rect 186294 511954 186914 547398
rect 186294 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 186914 511954
rect 186294 511634 186914 511718
rect 186294 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 186914 511634
rect 186294 475954 186914 511398
rect 186294 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 186914 475954
rect 186294 475634 186914 475718
rect 186294 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 186914 475634
rect 186294 439954 186914 475398
rect 186294 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 186914 439954
rect 186294 439634 186914 439718
rect 186294 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 186914 439634
rect 186294 403954 186914 439398
rect 186294 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 186914 403954
rect 186294 403634 186914 403718
rect 186294 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 186914 403634
rect 186294 367954 186914 403398
rect 186294 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 186914 367954
rect 186294 367634 186914 367718
rect 186294 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 186914 367634
rect 186294 331954 186914 367398
rect 186294 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 186914 331954
rect 186294 331634 186914 331718
rect 186294 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 186914 331634
rect 186294 295954 186914 331398
rect 186294 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 186914 295954
rect 186294 295634 186914 295718
rect 186294 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 186914 295634
rect 186294 259954 186914 295398
rect 186294 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 186914 259954
rect 186294 259634 186914 259718
rect 186294 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 186914 259634
rect 186294 223954 186914 259398
rect 186294 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 186914 223954
rect 186294 223634 186914 223718
rect 186294 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 186914 223634
rect 186294 187954 186914 223398
rect 186294 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 186914 187954
rect 186294 187634 186914 187718
rect 186294 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 186914 187634
rect 186294 151954 186914 187398
rect 186294 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 186914 151954
rect 186294 151634 186914 151718
rect 186294 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 186914 151634
rect 186294 142000 186914 151398
rect 190794 706758 191414 711590
rect 190794 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 191414 706758
rect 190794 706438 191414 706522
rect 190794 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 191414 706438
rect 190794 696454 191414 706202
rect 190794 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 191414 696454
rect 190794 696134 191414 696218
rect 190794 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 191414 696134
rect 190794 660454 191414 695898
rect 190794 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 191414 660454
rect 190794 660134 191414 660218
rect 190794 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 191414 660134
rect 190794 624454 191414 659898
rect 190794 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 191414 624454
rect 190794 624134 191414 624218
rect 190794 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 191414 624134
rect 190794 588454 191414 623898
rect 190794 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 191414 588454
rect 190794 588134 191414 588218
rect 190794 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 191414 588134
rect 190794 552454 191414 587898
rect 190794 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 191414 552454
rect 190794 552134 191414 552218
rect 190794 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 191414 552134
rect 190794 516454 191414 551898
rect 190794 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 191414 516454
rect 190794 516134 191414 516218
rect 190794 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 191414 516134
rect 190794 480454 191414 515898
rect 190794 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 191414 480454
rect 190794 480134 191414 480218
rect 190794 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 191414 480134
rect 190794 444454 191414 479898
rect 190794 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 191414 444454
rect 190794 444134 191414 444218
rect 190794 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 191414 444134
rect 190794 408454 191414 443898
rect 190794 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 191414 408454
rect 190794 408134 191414 408218
rect 190794 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 191414 408134
rect 190794 372454 191414 407898
rect 190794 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 191414 372454
rect 190794 372134 191414 372218
rect 190794 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 191414 372134
rect 190794 336454 191414 371898
rect 190794 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 191414 336454
rect 190794 336134 191414 336218
rect 190794 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 191414 336134
rect 190794 300454 191414 335898
rect 190794 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 191414 300454
rect 190794 300134 191414 300218
rect 190794 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 191414 300134
rect 190794 264454 191414 299898
rect 190794 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 191414 264454
rect 190794 264134 191414 264218
rect 190794 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 191414 264134
rect 190794 228454 191414 263898
rect 190794 228218 190826 228454
rect 191062 228218 191146 228454
rect 191382 228218 191414 228454
rect 190794 228134 191414 228218
rect 190794 227898 190826 228134
rect 191062 227898 191146 228134
rect 191382 227898 191414 228134
rect 190794 192454 191414 227898
rect 190794 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 191414 192454
rect 190794 192134 191414 192218
rect 190794 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 191414 192134
rect 190794 156454 191414 191898
rect 190794 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 191414 156454
rect 190794 156134 191414 156218
rect 190794 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 191414 156134
rect 190794 142000 191414 155898
rect 195294 707718 195914 711590
rect 195294 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 195914 707718
rect 195294 707398 195914 707482
rect 195294 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 195914 707398
rect 195294 700954 195914 707162
rect 195294 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 195914 700954
rect 195294 700634 195914 700718
rect 195294 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 195914 700634
rect 195294 664954 195914 700398
rect 195294 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 195914 664954
rect 195294 664634 195914 664718
rect 195294 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 195914 664634
rect 195294 628954 195914 664398
rect 195294 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 195914 628954
rect 195294 628634 195914 628718
rect 195294 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 195914 628634
rect 195294 592954 195914 628398
rect 195294 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 195914 592954
rect 195294 592634 195914 592718
rect 195294 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 195914 592634
rect 195294 556954 195914 592398
rect 195294 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 195914 556954
rect 195294 556634 195914 556718
rect 195294 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 195914 556634
rect 195294 520954 195914 556398
rect 195294 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 195914 520954
rect 195294 520634 195914 520718
rect 195294 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 195914 520634
rect 195294 484954 195914 520398
rect 195294 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 195914 484954
rect 195294 484634 195914 484718
rect 195294 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 195914 484634
rect 195294 448954 195914 484398
rect 195294 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 195914 448954
rect 195294 448634 195914 448718
rect 195294 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 195914 448634
rect 195294 412954 195914 448398
rect 195294 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 195914 412954
rect 195294 412634 195914 412718
rect 195294 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 195914 412634
rect 195294 376954 195914 412398
rect 195294 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 195914 376954
rect 195294 376634 195914 376718
rect 195294 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 195914 376634
rect 195294 340954 195914 376398
rect 195294 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 195914 340954
rect 195294 340634 195914 340718
rect 195294 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 195914 340634
rect 195294 304954 195914 340398
rect 195294 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 195914 304954
rect 195294 304634 195914 304718
rect 195294 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 195914 304634
rect 195294 268954 195914 304398
rect 195294 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 195914 268954
rect 195294 268634 195914 268718
rect 195294 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 195914 268634
rect 195294 232954 195914 268398
rect 195294 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 195914 232954
rect 195294 232634 195914 232718
rect 195294 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 195914 232634
rect 195294 196954 195914 232398
rect 195294 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 195914 196954
rect 195294 196634 195914 196718
rect 195294 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 195914 196634
rect 195294 160954 195914 196398
rect 195294 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 195914 160954
rect 195294 160634 195914 160718
rect 195294 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 195914 160634
rect 195294 124954 195914 160398
rect 195294 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 195914 124954
rect 195294 124634 195914 124718
rect 195294 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 195914 124634
rect 114294 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 114914 115954
rect 114294 115634 114914 115718
rect 114294 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 114914 115634
rect 114294 79954 114914 115398
rect 139568 115954 139888 115986
rect 139568 115718 139610 115954
rect 139846 115718 139888 115954
rect 139568 115634 139888 115718
rect 139568 115398 139610 115634
rect 139846 115398 139888 115634
rect 139568 115366 139888 115398
rect 170288 115954 170608 115986
rect 170288 115718 170330 115954
rect 170566 115718 170608 115954
rect 170288 115634 170608 115718
rect 170288 115398 170330 115634
rect 170566 115398 170608 115634
rect 170288 115366 170608 115398
rect 124208 111454 124528 111486
rect 124208 111218 124250 111454
rect 124486 111218 124528 111454
rect 124208 111134 124528 111218
rect 124208 110898 124250 111134
rect 124486 110898 124528 111134
rect 124208 110866 124528 110898
rect 154928 111454 155248 111486
rect 154928 111218 154970 111454
rect 155206 111218 155248 111454
rect 154928 111134 155248 111218
rect 154928 110898 154970 111134
rect 155206 110898 155248 111134
rect 154928 110866 155248 110898
rect 185648 111454 185968 111486
rect 185648 111218 185690 111454
rect 185926 111218 185968 111454
rect 185648 111134 185968 111218
rect 185648 110898 185690 111134
rect 185926 110898 185968 111134
rect 185648 110866 185968 110898
rect 195294 88954 195914 124398
rect 195294 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 195914 88954
rect 195294 88634 195914 88718
rect 195294 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 195914 88634
rect 176699 81020 176765 81021
rect 176699 80956 176700 81020
rect 176764 80956 176765 81020
rect 176699 80955 176765 80956
rect 175227 80476 175293 80477
rect 175227 80412 175228 80476
rect 175292 80412 175293 80476
rect 175227 80411 175293 80412
rect 134011 80204 134077 80205
rect 134011 80140 134012 80204
rect 134076 80140 134077 80204
rect 134011 80139 134077 80140
rect 143211 80204 143277 80205
rect 143211 80140 143212 80204
rect 143276 80140 143277 80204
rect 143211 80139 143277 80140
rect 149651 80204 149717 80205
rect 149651 80140 149652 80204
rect 149716 80140 149717 80204
rect 149651 80139 149717 80140
rect 170627 80204 170693 80205
rect 170627 80140 170628 80204
rect 170692 80140 170693 80204
rect 170627 80139 170693 80140
rect 133275 80068 133341 80069
rect 133275 80004 133276 80068
rect 133340 80004 133341 80068
rect 133275 80003 133341 80004
rect 114294 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 114914 79954
rect 131435 79932 131501 79933
rect 131435 79868 131436 79932
rect 131500 79930 131501 79932
rect 132723 79932 132789 79933
rect 131500 79870 131682 79930
rect 131500 79868 131501 79870
rect 131435 79867 131501 79868
rect 131435 79796 131501 79797
rect 131435 79732 131436 79796
rect 131500 79732 131501 79796
rect 131435 79731 131501 79732
rect 114294 79634 114914 79718
rect 114294 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 114914 79634
rect 114294 43954 114914 79398
rect 131251 78980 131317 78981
rect 131251 78916 131252 78980
rect 131316 78916 131317 78980
rect 131251 78915 131317 78916
rect 131067 78028 131133 78029
rect 114294 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 114914 43954
rect 114294 43634 114914 43718
rect 114294 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 114914 43634
rect 114294 7954 114914 43398
rect 114294 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 114914 7954
rect 114294 7634 114914 7718
rect 114294 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 114914 7634
rect 114294 -1306 114914 7398
rect 114294 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 114914 -1306
rect 114294 -1626 114914 -1542
rect 114294 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 114914 -1626
rect 114294 -7654 114914 -1862
rect 118794 48454 119414 78000
rect 118794 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 119414 48454
rect 118794 48134 119414 48218
rect 118794 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 119414 48134
rect 118794 12454 119414 47898
rect 118794 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 119414 12454
rect 118794 12134 119414 12218
rect 118794 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 119414 12134
rect 118794 -2266 119414 11898
rect 118794 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 119414 -2266
rect 118794 -2586 119414 -2502
rect 118794 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 119414 -2586
rect 118794 -7654 119414 -2822
rect 123294 52954 123914 78000
rect 123294 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 123914 52954
rect 123294 52634 123914 52718
rect 123294 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 123914 52634
rect 123294 16954 123914 52398
rect 123294 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 123914 16954
rect 123294 16634 123914 16718
rect 123294 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 123914 16634
rect 123294 -3226 123914 16398
rect 123294 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 123914 -3226
rect 123294 -3546 123914 -3462
rect 123294 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 123914 -3546
rect 123294 -7654 123914 -3782
rect 127794 57454 128414 78000
rect 131067 77964 131068 78028
rect 131132 77964 131133 78028
rect 131067 77963 131133 77964
rect 131070 75173 131130 77963
rect 131067 75172 131133 75173
rect 131067 75108 131068 75172
rect 131132 75108 131133 75172
rect 131067 75107 131133 75108
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -4186 128414 20898
rect 131254 8941 131314 78915
rect 131438 76533 131498 79731
rect 131435 76532 131501 76533
rect 131435 76468 131436 76532
rect 131500 76468 131501 76532
rect 131435 76467 131501 76468
rect 131251 8940 131317 8941
rect 131251 8876 131252 8940
rect 131316 8876 131317 8940
rect 131251 8875 131317 8876
rect 131622 4861 131682 79870
rect 132723 79868 132724 79932
rect 132788 79930 132789 79932
rect 132788 79870 133154 79930
rect 132788 79868 132789 79870
rect 132723 79867 132789 79868
rect 132294 61954 132914 78000
rect 132294 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 132914 61954
rect 132294 61634 132914 61718
rect 132294 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 132914 61634
rect 132294 25954 132914 61398
rect 132294 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 132914 25954
rect 132294 25634 132914 25718
rect 132294 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 132914 25634
rect 131619 4860 131685 4861
rect 131619 4796 131620 4860
rect 131684 4796 131685 4860
rect 131619 4795 131685 4796
rect 127794 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 128414 -4186
rect 127794 -4506 128414 -4422
rect 127794 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 128414 -4506
rect 127794 -7654 128414 -4742
rect 132294 -5146 132914 25398
rect 133094 7581 133154 79870
rect 133278 9077 133338 80003
rect 133643 79660 133709 79661
rect 133643 79596 133644 79660
rect 133708 79596 133709 79660
rect 133643 79595 133709 79596
rect 133459 78708 133525 78709
rect 133459 78644 133460 78708
rect 133524 78644 133525 78708
rect 133459 78643 133525 78644
rect 133462 73813 133522 78643
rect 133646 78437 133706 79595
rect 133643 78436 133709 78437
rect 133643 78372 133644 78436
rect 133708 78372 133709 78436
rect 133643 78371 133709 78372
rect 134014 75930 134074 80139
rect 134563 79932 134629 79933
rect 134563 79868 134564 79932
rect 134628 79868 134629 79932
rect 134563 79867 134629 79868
rect 135299 79932 135365 79933
rect 135299 79868 135300 79932
rect 135364 79868 135365 79932
rect 135299 79867 135365 79868
rect 137507 79932 137573 79933
rect 137507 79868 137508 79932
rect 137572 79868 137573 79932
rect 137507 79867 137573 79868
rect 137875 79932 137941 79933
rect 137875 79868 137876 79932
rect 137940 79868 137941 79932
rect 137875 79867 137941 79868
rect 141923 79932 141989 79933
rect 141923 79868 141924 79932
rect 141988 79868 141989 79932
rect 141923 79867 141989 79868
rect 134195 79796 134261 79797
rect 134195 79732 134196 79796
rect 134260 79794 134261 79796
rect 134260 79734 134442 79794
rect 134260 79732 134261 79734
rect 134195 79731 134261 79732
rect 134195 78028 134261 78029
rect 134195 77964 134196 78028
rect 134260 77964 134261 78028
rect 134195 77963 134261 77964
rect 133830 75870 134074 75930
rect 133830 75309 133890 75870
rect 133827 75308 133893 75309
rect 133827 75244 133828 75308
rect 133892 75244 133893 75308
rect 133827 75243 133893 75244
rect 134198 73949 134258 77963
rect 134195 73948 134261 73949
rect 134195 73884 134196 73948
rect 134260 73884 134261 73948
rect 134195 73883 134261 73884
rect 133459 73812 133525 73813
rect 133459 73748 133460 73812
rect 133524 73748 133525 73812
rect 133459 73747 133525 73748
rect 134382 9213 134442 79734
rect 134566 78165 134626 79867
rect 135302 79525 135362 79867
rect 135483 79796 135549 79797
rect 135483 79732 135484 79796
rect 135548 79732 135549 79796
rect 135483 79731 135549 79732
rect 135299 79524 135365 79525
rect 135299 79460 135300 79524
rect 135364 79460 135365 79524
rect 135299 79459 135365 79460
rect 134563 78164 134629 78165
rect 134563 78100 134564 78164
rect 134628 78100 134629 78164
rect 134563 78099 134629 78100
rect 135299 78028 135365 78029
rect 135299 77964 135300 78028
rect 135364 77964 135365 78028
rect 135299 77963 135365 77964
rect 134379 9212 134445 9213
rect 134379 9148 134380 9212
rect 134444 9148 134445 9212
rect 134379 9147 134445 9148
rect 133275 9076 133341 9077
rect 133275 9012 133276 9076
rect 133340 9012 133341 9076
rect 133275 9011 133341 9012
rect 133091 7580 133157 7581
rect 133091 7516 133092 7580
rect 133156 7516 133157 7580
rect 133091 7515 133157 7516
rect 135302 6221 135362 77963
rect 135486 9349 135546 79731
rect 135667 78028 135733 78029
rect 135667 77964 135668 78028
rect 135732 77964 135733 78028
rect 135667 77963 135733 77964
rect 135670 22677 135730 77963
rect 136794 66454 137414 78000
rect 136794 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 137414 66454
rect 136794 66134 137414 66218
rect 136794 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 137414 66134
rect 136794 30454 137414 65898
rect 136794 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 137414 30454
rect 136794 30134 137414 30218
rect 136794 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 137414 30134
rect 135667 22676 135733 22677
rect 135667 22612 135668 22676
rect 135732 22612 135733 22676
rect 135667 22611 135733 22612
rect 135483 9348 135549 9349
rect 135483 9284 135484 9348
rect 135548 9284 135549 9348
rect 135483 9283 135549 9284
rect 135299 6220 135365 6221
rect 135299 6156 135300 6220
rect 135364 6156 135365 6220
rect 135299 6155 135365 6156
rect 132294 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 132914 -5146
rect 132294 -5466 132914 -5382
rect 132294 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 132914 -5466
rect 132294 -7654 132914 -5702
rect 136794 -6106 137414 29898
rect 137510 9485 137570 79867
rect 137878 78437 137938 79867
rect 138059 79796 138125 79797
rect 138059 79732 138060 79796
rect 138124 79732 138125 79796
rect 138059 79731 138125 79732
rect 138427 79796 138493 79797
rect 138427 79732 138428 79796
rect 138492 79732 138493 79796
rect 138427 79731 138493 79732
rect 137875 78436 137941 78437
rect 137875 78372 137876 78436
rect 137940 78372 137941 78436
rect 137875 78371 137941 78372
rect 138062 76805 138122 79731
rect 138243 78708 138309 78709
rect 138243 78644 138244 78708
rect 138308 78644 138309 78708
rect 138243 78643 138309 78644
rect 138059 76804 138125 76805
rect 138059 76740 138060 76804
rect 138124 76740 138125 76804
rect 138059 76739 138125 76740
rect 138246 21317 138306 78643
rect 138243 21316 138309 21317
rect 138243 21252 138244 21316
rect 138308 21252 138309 21316
rect 138243 21251 138309 21252
rect 137507 9484 137573 9485
rect 137507 9420 137508 9484
rect 137572 9420 137573 9484
rect 137507 9419 137573 9420
rect 138430 4997 138490 79731
rect 139715 79660 139781 79661
rect 139715 79596 139716 79660
rect 139780 79596 139781 79660
rect 139715 79595 139781 79596
rect 139899 79660 139965 79661
rect 139899 79596 139900 79660
rect 139964 79596 139965 79660
rect 139899 79595 139965 79596
rect 139163 78028 139229 78029
rect 139163 77964 139164 78028
rect 139228 77964 139229 78028
rect 139163 77963 139229 77964
rect 138427 4996 138493 4997
rect 138427 4932 138428 4996
rect 138492 4932 138493 4996
rect 138427 4931 138493 4932
rect 139166 3637 139226 77963
rect 139531 75308 139597 75309
rect 139531 75244 139532 75308
rect 139596 75244 139597 75308
rect 139531 75243 139597 75244
rect 139534 7717 139594 75243
rect 139718 10301 139778 79595
rect 139715 10300 139781 10301
rect 139715 10236 139716 10300
rect 139780 10236 139781 10300
rect 139715 10235 139781 10236
rect 139531 7716 139597 7717
rect 139531 7652 139532 7716
rect 139596 7652 139597 7716
rect 139531 7651 139597 7652
rect 139163 3636 139229 3637
rect 139163 3572 139164 3636
rect 139228 3572 139229 3636
rect 139163 3571 139229 3572
rect 139902 3365 139962 79595
rect 141926 78981 141986 79867
rect 142107 79660 142173 79661
rect 142107 79596 142108 79660
rect 142172 79596 142173 79660
rect 142107 79595 142173 79596
rect 141923 78980 141989 78981
rect 141923 78916 141924 78980
rect 141988 78916 141989 78980
rect 141923 78915 141989 78916
rect 141003 76532 141069 76533
rect 141003 76468 141004 76532
rect 141068 76468 141069 76532
rect 141003 76467 141069 76468
rect 140819 75308 140885 75309
rect 140819 75244 140820 75308
rect 140884 75244 140885 75308
rect 140819 75243 140885 75244
rect 140822 44301 140882 75243
rect 140819 44300 140885 44301
rect 140819 44236 140820 44300
rect 140884 44236 140885 44300
rect 140819 44235 140885 44236
rect 141006 3501 141066 76467
rect 141294 70954 141914 78000
rect 142110 75037 142170 79595
rect 143027 76804 143093 76805
rect 143027 76740 143028 76804
rect 143092 76740 143093 76804
rect 143027 76739 143093 76740
rect 142843 76668 142909 76669
rect 142843 76604 142844 76668
rect 142908 76604 142909 76668
rect 142843 76603 142909 76604
rect 142107 75036 142173 75037
rect 142107 74972 142108 75036
rect 142172 74972 142173 75036
rect 142107 74971 142173 74972
rect 141294 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 141914 70954
rect 141294 70634 141914 70718
rect 141294 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 141914 70634
rect 141294 34954 141914 70398
rect 142846 66197 142906 76603
rect 142843 66196 142909 66197
rect 142843 66132 142844 66196
rect 142908 66132 142909 66196
rect 142843 66131 142909 66132
rect 141294 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 141914 34954
rect 141294 34634 141914 34718
rect 141294 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 141914 34634
rect 141003 3500 141069 3501
rect 141003 3436 141004 3500
rect 141068 3436 141069 3500
rect 141003 3435 141069 3436
rect 139899 3364 139965 3365
rect 139899 3300 139900 3364
rect 139964 3300 139965 3364
rect 139899 3299 139965 3300
rect 136794 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 137414 -6106
rect 136794 -6426 137414 -6342
rect 136794 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 137414 -6426
rect 136794 -7654 137414 -6662
rect 141294 -7066 141914 34398
rect 143030 4997 143090 76739
rect 143027 4996 143093 4997
rect 143027 4932 143028 4996
rect 143092 4932 143093 4996
rect 143027 4931 143093 4932
rect 143214 4861 143274 80139
rect 143763 79932 143829 79933
rect 143763 79868 143764 79932
rect 143828 79868 143829 79932
rect 143763 79867 143829 79868
rect 144499 79932 144565 79933
rect 144499 79868 144500 79932
rect 144564 79868 144565 79932
rect 144499 79867 144565 79868
rect 146891 79932 146957 79933
rect 146891 79868 146892 79932
rect 146956 79868 146957 79932
rect 146891 79867 146957 79868
rect 147995 79932 148061 79933
rect 147995 79868 147996 79932
rect 148060 79868 148061 79932
rect 147995 79867 148061 79868
rect 148179 79932 148245 79933
rect 148179 79868 148180 79932
rect 148244 79868 148245 79932
rect 148915 79932 148981 79933
rect 148915 79930 148916 79932
rect 148179 79867 148245 79868
rect 148734 79870 148916 79930
rect 143395 79796 143461 79797
rect 143395 79732 143396 79796
rect 143460 79732 143461 79796
rect 143395 79731 143461 79732
rect 143211 4860 143277 4861
rect 143211 4796 143212 4860
rect 143276 4796 143277 4860
rect 143211 4795 143277 4796
rect 143398 3365 143458 79731
rect 143766 78165 143826 79867
rect 144502 78437 144562 79867
rect 144683 79660 144749 79661
rect 144683 79596 144684 79660
rect 144748 79596 144749 79660
rect 144683 79595 144749 79596
rect 144499 78436 144565 78437
rect 144499 78372 144500 78436
rect 144564 78372 144565 78436
rect 144499 78371 144565 78372
rect 144686 78298 144746 79595
rect 144502 78238 144746 78298
rect 143763 78164 143829 78165
rect 143763 78100 143764 78164
rect 143828 78100 143829 78164
rect 143763 78099 143829 78100
rect 144315 76668 144381 76669
rect 144315 76604 144316 76668
rect 144380 76604 144381 76668
rect 144315 76603 144381 76604
rect 144318 69597 144378 76603
rect 144315 69596 144381 69597
rect 144315 69532 144316 69596
rect 144380 69532 144381 69596
rect 144315 69531 144381 69532
rect 144502 65517 144562 78238
rect 144683 78164 144749 78165
rect 144683 78100 144684 78164
rect 144748 78100 144749 78164
rect 144683 78099 144749 78100
rect 144499 65516 144565 65517
rect 144499 65452 144500 65516
rect 144564 65452 144565 65516
rect 144499 65451 144565 65452
rect 144686 25669 144746 78099
rect 145419 77484 145485 77485
rect 145419 77420 145420 77484
rect 145484 77420 145485 77484
rect 145419 77419 145485 77420
rect 145235 77348 145301 77349
rect 145235 77284 145236 77348
rect 145300 77284 145301 77348
rect 145235 77283 145301 77284
rect 145238 62797 145298 77283
rect 145235 62796 145301 62797
rect 145235 62732 145236 62796
rect 145300 62732 145301 62796
rect 145235 62731 145301 62732
rect 144683 25668 144749 25669
rect 144683 25604 144684 25668
rect 144748 25604 144749 25668
rect 144683 25603 144749 25604
rect 145422 24445 145482 77419
rect 145794 75454 146414 78000
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145603 75172 145669 75173
rect 145603 75108 145604 75172
rect 145668 75108 145669 75172
rect 145603 75107 145669 75108
rect 145794 75134 146414 75218
rect 145419 24444 145485 24445
rect 145419 24380 145420 24444
rect 145484 24380 145485 24444
rect 145419 24379 145485 24380
rect 145606 6901 145666 75107
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145603 6900 145669 6901
rect 145603 6836 145604 6900
rect 145668 6836 145669 6900
rect 145603 6835 145669 6836
rect 145794 3454 146414 38898
rect 146894 3773 146954 79867
rect 147075 77484 147141 77485
rect 147075 77420 147076 77484
rect 147140 77420 147141 77484
rect 147075 77419 147141 77420
rect 147078 28253 147138 77419
rect 147259 77348 147325 77349
rect 147259 77284 147260 77348
rect 147324 77284 147325 77348
rect 147259 77283 147325 77284
rect 147075 28252 147141 28253
rect 147075 28188 147076 28252
rect 147140 28188 147141 28252
rect 147075 28187 147141 28188
rect 147262 18733 147322 77283
rect 147998 76669 148058 79867
rect 147995 76668 148061 76669
rect 147995 76604 147996 76668
rect 148060 76604 148061 76668
rect 147995 76603 148061 76604
rect 148182 75445 148242 79867
rect 148547 76668 148613 76669
rect 148547 76604 148548 76668
rect 148612 76604 148613 76668
rect 148547 76603 148613 76604
rect 148179 75444 148245 75445
rect 148179 75380 148180 75444
rect 148244 75380 148245 75444
rect 148179 75379 148245 75380
rect 148550 29613 148610 76603
rect 148547 29612 148613 29613
rect 148547 29548 148548 29612
rect 148612 29548 148613 29612
rect 148547 29547 148613 29548
rect 147259 18732 147325 18733
rect 147259 18668 147260 18732
rect 147324 18668 147325 18732
rect 147259 18667 147325 18668
rect 148734 6085 148794 79870
rect 148915 79868 148916 79870
rect 148980 79868 148981 79932
rect 148915 79867 148981 79868
rect 148915 79796 148981 79797
rect 148915 79732 148916 79796
rect 148980 79732 148981 79796
rect 148915 79731 148981 79732
rect 148731 6084 148797 6085
rect 148731 6020 148732 6084
rect 148796 6020 148797 6084
rect 148731 6019 148797 6020
rect 148918 5269 148978 79731
rect 149654 73949 149714 80139
rect 161243 80068 161309 80069
rect 161243 80004 161244 80068
rect 161308 80004 161309 80068
rect 166763 80068 166829 80069
rect 166763 80066 166764 80068
rect 161243 80003 161309 80004
rect 166582 80006 166764 80066
rect 151123 79932 151189 79933
rect 151123 79868 151124 79932
rect 151188 79868 151189 79932
rect 151123 79867 151189 79868
rect 151491 79932 151557 79933
rect 151491 79868 151492 79932
rect 151556 79868 151557 79932
rect 151491 79867 151557 79868
rect 151675 79932 151741 79933
rect 151675 79868 151676 79932
rect 151740 79868 151741 79932
rect 151675 79867 151741 79868
rect 152779 79932 152845 79933
rect 152779 79868 152780 79932
rect 152844 79930 152845 79932
rect 153699 79932 153765 79933
rect 152844 79870 153026 79930
rect 152844 79868 152845 79870
rect 152779 79867 152845 79868
rect 150203 79796 150269 79797
rect 150203 79794 150204 79796
rect 149838 79734 150204 79794
rect 149651 73948 149717 73949
rect 149651 73884 149652 73948
rect 149716 73884 149717 73948
rect 149651 73883 149717 73884
rect 149838 7581 149898 79734
rect 150203 79732 150204 79734
rect 150268 79732 150269 79796
rect 150203 79731 150269 79732
rect 150019 78708 150085 78709
rect 150019 78644 150020 78708
rect 150084 78644 150085 78708
rect 150019 78643 150085 78644
rect 149835 7580 149901 7581
rect 149835 7516 149836 7580
rect 149900 7516 149901 7580
rect 149835 7515 149901 7516
rect 150022 6765 150082 78643
rect 150294 43954 150914 78000
rect 151126 76669 151186 79867
rect 151307 79796 151373 79797
rect 151307 79732 151308 79796
rect 151372 79732 151373 79796
rect 151307 79731 151373 79732
rect 151123 76668 151189 76669
rect 151123 76604 151124 76668
rect 151188 76604 151189 76668
rect 151123 76603 151189 76604
rect 150294 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 150914 43954
rect 150294 43634 150914 43718
rect 150294 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 150914 43634
rect 150294 7954 150914 43398
rect 151310 30973 151370 79731
rect 151494 78437 151554 79867
rect 151491 78436 151557 78437
rect 151491 78372 151492 78436
rect 151556 78372 151557 78436
rect 151491 78371 151557 78372
rect 151491 76668 151557 76669
rect 151491 76604 151492 76668
rect 151556 76604 151557 76668
rect 151491 76603 151557 76604
rect 151307 30972 151373 30973
rect 151307 30908 151308 30972
rect 151372 30908 151373 30972
rect 151307 30907 151373 30908
rect 151494 20229 151554 76603
rect 151491 20228 151557 20229
rect 151491 20164 151492 20228
rect 151556 20164 151557 20228
rect 151491 20163 151557 20164
rect 151678 9213 151738 79867
rect 152411 77484 152477 77485
rect 152411 77420 152412 77484
rect 152476 77420 152477 77484
rect 152411 77419 152477 77420
rect 152414 73813 152474 77419
rect 152779 77348 152845 77349
rect 152779 77284 152780 77348
rect 152844 77284 152845 77348
rect 152779 77283 152845 77284
rect 152411 73812 152477 73813
rect 152411 73748 152412 73812
rect 152476 73748 152477 73812
rect 152411 73747 152477 73748
rect 152782 26893 152842 77283
rect 152779 26892 152845 26893
rect 152779 26828 152780 26892
rect 152844 26828 152845 26892
rect 152779 26827 152845 26828
rect 152966 10437 153026 79870
rect 153699 79868 153700 79932
rect 153764 79868 153765 79932
rect 153699 79867 153765 79868
rect 154435 79932 154501 79933
rect 154435 79868 154436 79932
rect 154500 79868 154501 79932
rect 154435 79867 154501 79868
rect 154619 79932 154685 79933
rect 154619 79868 154620 79932
rect 154684 79868 154685 79932
rect 154619 79867 154685 79868
rect 155355 79932 155421 79933
rect 155355 79868 155356 79932
rect 155420 79868 155421 79932
rect 155355 79867 155421 79868
rect 155539 79932 155605 79933
rect 155539 79868 155540 79932
rect 155604 79868 155605 79932
rect 155539 79867 155605 79868
rect 156275 79932 156341 79933
rect 156275 79868 156276 79932
rect 156340 79868 156341 79932
rect 156275 79867 156341 79868
rect 156827 79932 156893 79933
rect 156827 79868 156828 79932
rect 156892 79868 156893 79932
rect 156827 79867 156893 79868
rect 158115 79932 158181 79933
rect 158115 79868 158116 79932
rect 158180 79868 158181 79932
rect 158115 79867 158181 79868
rect 159587 79932 159653 79933
rect 159587 79868 159588 79932
rect 159652 79868 159653 79932
rect 159587 79867 159653 79868
rect 160691 79932 160757 79933
rect 160691 79868 160692 79932
rect 160756 79868 160757 79932
rect 160691 79867 160757 79868
rect 153702 77349 153762 79867
rect 154067 79796 154133 79797
rect 154067 79732 154068 79796
rect 154132 79732 154133 79796
rect 154067 79731 154133 79732
rect 154070 77482 154130 79731
rect 153886 77422 154130 77482
rect 154251 77484 154317 77485
rect 153699 77348 153765 77349
rect 153699 77284 153700 77348
rect 153764 77284 153765 77348
rect 153699 77283 153765 77284
rect 152963 10436 153029 10437
rect 152963 10372 152964 10436
rect 153028 10372 153029 10436
rect 152963 10371 153029 10372
rect 151675 9212 151741 9213
rect 151675 9148 151676 9212
rect 151740 9148 151741 9212
rect 151675 9147 151741 9148
rect 150294 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 150914 7954
rect 150294 7634 150914 7718
rect 150294 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 150914 7634
rect 150019 6764 150085 6765
rect 150019 6700 150020 6764
rect 150084 6700 150085 6764
rect 150019 6699 150085 6700
rect 148915 5268 148981 5269
rect 148915 5204 148916 5268
rect 148980 5204 148981 5268
rect 148915 5203 148981 5204
rect 146891 3772 146957 3773
rect 146891 3708 146892 3772
rect 146956 3708 146957 3772
rect 146891 3707 146957 3708
rect 143395 3364 143461 3365
rect 143395 3300 143396 3364
rect 143460 3300 143461 3364
rect 143395 3299 143461 3300
rect 141294 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 141914 -7066
rect 141294 -7386 141914 -7302
rect 141294 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 141914 -7386
rect 141294 -7654 141914 -7622
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 150294 -1306 150914 7398
rect 153886 6629 153946 77422
rect 154251 77420 154252 77484
rect 154316 77420 154317 77484
rect 154251 77419 154317 77420
rect 154067 77348 154133 77349
rect 154067 77284 154068 77348
rect 154132 77284 154133 77348
rect 154067 77283 154133 77284
rect 154070 55861 154130 77283
rect 154067 55860 154133 55861
rect 154067 55796 154068 55860
rect 154132 55796 154133 55860
rect 154067 55795 154133 55796
rect 154254 16149 154314 77419
rect 154438 76669 154498 79867
rect 154622 77349 154682 79867
rect 155358 78165 155418 79867
rect 155355 78164 155421 78165
rect 155355 78100 155356 78164
rect 155420 78100 155421 78164
rect 155355 78099 155421 78100
rect 154619 77348 154685 77349
rect 154619 77284 154620 77348
rect 154684 77284 154685 77348
rect 154619 77283 154685 77284
rect 154435 76668 154501 76669
rect 154435 76604 154436 76668
rect 154500 76604 154501 76668
rect 154435 76603 154501 76604
rect 154794 48454 155414 78000
rect 154794 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 155414 48454
rect 154794 48134 155414 48218
rect 154794 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 155414 48134
rect 154251 16148 154317 16149
rect 154251 16084 154252 16148
rect 154316 16084 154317 16148
rect 154251 16083 154317 16084
rect 154794 12454 155414 47898
rect 154794 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 155414 12454
rect 155542 12341 155602 79867
rect 156278 77349 156338 79867
rect 156643 77620 156709 77621
rect 156643 77556 156644 77620
rect 156708 77556 156709 77620
rect 156643 77555 156709 77556
rect 156275 77348 156341 77349
rect 156275 77284 156276 77348
rect 156340 77284 156341 77348
rect 156275 77283 156341 77284
rect 156646 13157 156706 77555
rect 156643 13156 156709 13157
rect 156643 13092 156644 13156
rect 156708 13092 156709 13156
rect 156643 13091 156709 13092
rect 155539 12340 155605 12341
rect 155539 12276 155540 12340
rect 155604 12276 155605 12340
rect 155539 12275 155605 12276
rect 154794 12134 155414 12218
rect 156830 12205 156890 79867
rect 157195 79524 157261 79525
rect 157195 79460 157196 79524
rect 157260 79460 157261 79524
rect 157195 79459 157261 79460
rect 157011 77484 157077 77485
rect 157011 77420 157012 77484
rect 157076 77420 157077 77484
rect 157011 77419 157077 77420
rect 156827 12204 156893 12205
rect 156827 12140 156828 12204
rect 156892 12140 156893 12204
rect 156827 12139 156893 12140
rect 154794 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 155414 12134
rect 153883 6628 153949 6629
rect 153883 6564 153884 6628
rect 153948 6564 153949 6628
rect 153883 6563 153949 6564
rect 150294 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 150914 -1306
rect 150294 -1626 150914 -1542
rect 150294 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 150914 -1626
rect 150294 -7654 150914 -1862
rect 154794 -2266 155414 11898
rect 157014 9077 157074 77419
rect 157011 9076 157077 9077
rect 157011 9012 157012 9076
rect 157076 9012 157077 9076
rect 157011 9011 157077 9012
rect 157198 5133 157258 79459
rect 157931 78708 157997 78709
rect 157931 78644 157932 78708
rect 157996 78644 157997 78708
rect 157931 78643 157997 78644
rect 157934 20093 157994 78643
rect 157931 20092 157997 20093
rect 157931 20028 157932 20092
rect 157996 20028 157997 20092
rect 157931 20027 157997 20028
rect 158118 14925 158178 79867
rect 158299 79796 158365 79797
rect 158299 79732 158300 79796
rect 158364 79732 158365 79796
rect 158299 79731 158365 79732
rect 158115 14924 158181 14925
rect 158115 14860 158116 14924
rect 158180 14860 158181 14924
rect 158115 14859 158181 14860
rect 158302 14789 158362 79731
rect 158851 79660 158917 79661
rect 158851 79596 158852 79660
rect 158916 79596 158917 79660
rect 158851 79595 158917 79596
rect 158483 77348 158549 77349
rect 158483 77284 158484 77348
rect 158548 77284 158549 77348
rect 158483 77283 158549 77284
rect 158299 14788 158365 14789
rect 158299 14724 158300 14788
rect 158364 14724 158365 14788
rect 158299 14723 158365 14724
rect 158486 12069 158546 77283
rect 158854 68237 158914 79595
rect 159590 79525 159650 79867
rect 159587 79524 159653 79525
rect 159587 79460 159588 79524
rect 159652 79460 159653 79524
rect 159587 79459 159653 79460
rect 159035 77348 159101 77349
rect 159035 77284 159036 77348
rect 159100 77284 159101 77348
rect 159035 77283 159101 77284
rect 158851 68236 158917 68237
rect 158851 68172 158852 68236
rect 158916 68172 158917 68236
rect 158851 68171 158917 68172
rect 159038 23085 159098 77283
rect 159294 52954 159914 78000
rect 160694 76533 160754 79867
rect 161059 79796 161125 79797
rect 161059 79732 161060 79796
rect 161124 79732 161125 79796
rect 161059 79731 161125 79732
rect 160875 79524 160941 79525
rect 160875 79460 160876 79524
rect 160940 79460 160941 79524
rect 160875 79459 160941 79460
rect 160691 76532 160757 76533
rect 160691 76468 160692 76532
rect 160756 76468 160757 76532
rect 160691 76467 160757 76468
rect 159294 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 159914 52954
rect 159294 52634 159914 52718
rect 159294 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 159914 52634
rect 159035 23084 159101 23085
rect 159035 23020 159036 23084
rect 159100 23020 159101 23084
rect 159035 23019 159101 23020
rect 159294 16954 159914 52398
rect 159294 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 159914 16954
rect 159294 16634 159914 16718
rect 159294 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 159914 16634
rect 158483 12068 158549 12069
rect 158483 12004 158484 12068
rect 158548 12004 158549 12068
rect 158483 12003 158549 12004
rect 157195 5132 157261 5133
rect 157195 5068 157196 5132
rect 157260 5068 157261 5132
rect 157195 5067 157261 5068
rect 154794 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 155414 -2266
rect 154794 -2586 155414 -2502
rect 154794 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 155414 -2586
rect 154794 -7654 155414 -2822
rect 159294 -3226 159914 16398
rect 160878 16013 160938 79459
rect 160875 16012 160941 16013
rect 160875 15948 160876 16012
rect 160940 15948 160941 16012
rect 160875 15947 160941 15948
rect 161062 14653 161122 79731
rect 161059 14652 161125 14653
rect 161059 14588 161060 14652
rect 161124 14588 161125 14652
rect 161059 14587 161125 14588
rect 161246 11933 161306 80003
rect 161979 79932 162045 79933
rect 161979 79868 161980 79932
rect 162044 79868 162045 79932
rect 161979 79867 162045 79868
rect 162347 79932 162413 79933
rect 162347 79868 162348 79932
rect 162412 79868 162413 79932
rect 162347 79867 162413 79868
rect 163267 79932 163333 79933
rect 163267 79868 163268 79932
rect 163332 79868 163333 79932
rect 163267 79867 163333 79868
rect 164739 79932 164805 79933
rect 164739 79868 164740 79932
rect 164804 79868 164805 79932
rect 164739 79867 164805 79868
rect 161982 77621 162042 79867
rect 161979 77620 162045 77621
rect 161979 77556 161980 77620
rect 162044 77556 162045 77620
rect 161979 77555 162045 77556
rect 162163 76260 162229 76261
rect 162163 76196 162164 76260
rect 162228 76196 162229 76260
rect 162163 76195 162229 76196
rect 162166 22949 162226 76195
rect 162163 22948 162229 22949
rect 162163 22884 162164 22948
rect 162228 22884 162229 22948
rect 162163 22883 162229 22884
rect 162350 17645 162410 79867
rect 162531 78300 162597 78301
rect 162531 78236 162532 78300
rect 162596 78236 162597 78300
rect 162531 78235 162597 78236
rect 162534 17781 162594 78235
rect 162715 76124 162781 76125
rect 162715 76060 162716 76124
rect 162780 76060 162781 76124
rect 162715 76059 162781 76060
rect 162531 17780 162597 17781
rect 162531 17716 162532 17780
rect 162596 17716 162597 17780
rect 162531 17715 162597 17716
rect 162347 17644 162413 17645
rect 162347 17580 162348 17644
rect 162412 17580 162413 17644
rect 162347 17579 162413 17580
rect 162718 15877 162778 76059
rect 163270 75445 163330 79867
rect 164003 79796 164069 79797
rect 164003 79732 164004 79796
rect 164068 79732 164069 79796
rect 164003 79731 164069 79732
rect 163635 78980 163701 78981
rect 163635 78916 163636 78980
rect 163700 78916 163701 78980
rect 163635 78915 163701 78916
rect 163451 78708 163517 78709
rect 163451 78644 163452 78708
rect 163516 78644 163517 78708
rect 163451 78643 163517 78644
rect 163267 75444 163333 75445
rect 163267 75380 163268 75444
rect 163332 75380 163333 75444
rect 163267 75379 163333 75380
rect 163454 36549 163514 78643
rect 163451 36548 163517 36549
rect 163451 36484 163452 36548
rect 163516 36484 163517 36548
rect 163451 36483 163517 36484
rect 163638 18597 163698 78915
rect 164006 78301 164066 79731
rect 164555 79524 164621 79525
rect 164555 79460 164556 79524
rect 164620 79460 164621 79524
rect 164555 79459 164621 79460
rect 164003 78300 164069 78301
rect 164003 78236 164004 78300
rect 164068 78236 164069 78300
rect 164003 78235 164069 78236
rect 163794 57454 164414 78000
rect 164558 77893 164618 79459
rect 164555 77892 164621 77893
rect 164555 77828 164556 77892
rect 164620 77828 164621 77892
rect 164555 77827 164621 77828
rect 164742 76261 164802 79867
rect 165107 79796 165173 79797
rect 165107 79732 165108 79796
rect 165172 79732 165173 79796
rect 165475 79796 165541 79797
rect 165475 79794 165476 79796
rect 165107 79731 165173 79732
rect 165294 79734 165476 79794
rect 164923 78028 164989 78029
rect 164923 77964 164924 78028
rect 164988 77964 164989 78028
rect 164923 77963 164989 77964
rect 164739 76260 164805 76261
rect 164739 76196 164740 76260
rect 164804 76196 164805 76260
rect 164739 76195 164805 76196
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163635 18596 163701 18597
rect 163635 18532 163636 18596
rect 163700 18532 163701 18596
rect 163635 18531 163701 18532
rect 162715 15876 162781 15877
rect 162715 15812 162716 15876
rect 162780 15812 162781 15876
rect 162715 15811 162781 15812
rect 161243 11932 161309 11933
rect 161243 11868 161244 11932
rect 161308 11868 161309 11932
rect 161243 11867 161309 11868
rect 159294 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 159914 -3226
rect 159294 -3546 159914 -3462
rect 159294 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 159914 -3546
rect 159294 -7654 159914 -3782
rect 163794 -4186 164414 20898
rect 164926 19957 164986 77963
rect 164923 19956 164989 19957
rect 164923 19892 164924 19956
rect 164988 19892 164989 19956
rect 164923 19891 164989 19892
rect 165110 11797 165170 79731
rect 165107 11796 165173 11797
rect 165107 11732 165108 11796
rect 165172 11732 165173 11796
rect 165107 11731 165173 11732
rect 165294 6493 165354 79734
rect 165475 79732 165476 79734
rect 165540 79732 165541 79796
rect 165475 79731 165541 79732
rect 165475 78028 165541 78029
rect 165475 77964 165476 78028
rect 165540 77964 165541 78028
rect 165475 77963 165541 77964
rect 165291 6492 165357 6493
rect 165291 6428 165292 6492
rect 165356 6428 165357 6492
rect 165291 6427 165357 6428
rect 165478 4997 165538 77963
rect 166395 77620 166461 77621
rect 166395 77556 166396 77620
rect 166460 77556 166461 77620
rect 166395 77555 166461 77556
rect 166211 77348 166277 77349
rect 166211 77284 166212 77348
rect 166276 77284 166277 77348
rect 166211 77283 166277 77284
rect 166214 8941 166274 77283
rect 166398 17509 166458 77555
rect 166395 17508 166461 17509
rect 166395 17444 166396 17508
rect 166460 17444 166461 17508
rect 166395 17443 166461 17444
rect 166582 14517 166642 80006
rect 166763 80004 166764 80006
rect 166828 80004 166829 80068
rect 166763 80003 166829 80004
rect 167315 79932 167381 79933
rect 167315 79868 167316 79932
rect 167380 79868 167381 79932
rect 167315 79867 167381 79868
rect 168051 79932 168117 79933
rect 168051 79868 168052 79932
rect 168116 79868 168117 79932
rect 168051 79867 168117 79868
rect 168971 79932 169037 79933
rect 168971 79868 168972 79932
rect 169036 79868 169037 79932
rect 168971 79867 169037 79868
rect 170259 79932 170325 79933
rect 170259 79868 170260 79932
rect 170324 79868 170325 79932
rect 170259 79867 170325 79868
rect 166763 77484 166829 77485
rect 166763 77420 166764 77484
rect 166828 77420 166829 77484
rect 166763 77419 166829 77420
rect 166766 75717 166826 77419
rect 167318 77349 167378 79867
rect 167683 79796 167749 79797
rect 167683 79732 167684 79796
rect 167748 79732 167749 79796
rect 167683 79731 167749 79732
rect 167315 77348 167381 77349
rect 167315 77284 167316 77348
rect 167380 77284 167381 77348
rect 167315 77283 167381 77284
rect 166763 75716 166829 75717
rect 166763 75652 166764 75716
rect 166828 75652 166829 75716
rect 166763 75651 166829 75652
rect 167686 64293 167746 79731
rect 167867 79524 167933 79525
rect 167867 79460 167868 79524
rect 167932 79460 167933 79524
rect 167867 79459 167933 79460
rect 167683 64292 167749 64293
rect 167683 64228 167684 64292
rect 167748 64228 167749 64292
rect 167683 64227 167749 64228
rect 166579 14516 166645 14517
rect 166579 14452 166580 14516
rect 166644 14452 166645 14516
rect 166579 14451 166645 14452
rect 167870 13021 167930 79459
rect 167867 13020 167933 13021
rect 167867 12956 167868 13020
rect 167932 12956 167933 13020
rect 167867 12955 167933 12956
rect 168054 10301 168114 79867
rect 168974 78709 169034 79867
rect 169339 79524 169405 79525
rect 169339 79460 169340 79524
rect 169404 79460 169405 79524
rect 169339 79459 169405 79460
rect 169523 79524 169589 79525
rect 169523 79460 169524 79524
rect 169588 79460 169589 79524
rect 169523 79459 169589 79460
rect 168971 78708 169037 78709
rect 168971 78644 168972 78708
rect 169036 78644 169037 78708
rect 168971 78643 169037 78644
rect 168294 61954 168914 78000
rect 169342 63613 169402 79459
rect 169339 63612 169405 63613
rect 169339 63548 169340 63612
rect 169404 63548 169405 63612
rect 169339 63547 169405 63548
rect 168294 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 168914 61954
rect 168294 61634 168914 61718
rect 168294 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 168914 61634
rect 168294 25954 168914 61398
rect 168294 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 168914 25954
rect 168294 25634 168914 25718
rect 168294 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 168914 25634
rect 168051 10300 168117 10301
rect 168051 10236 168052 10300
rect 168116 10236 168117 10300
rect 168051 10235 168117 10236
rect 166211 8940 166277 8941
rect 166211 8876 166212 8940
rect 166276 8876 166277 8940
rect 166211 8875 166277 8876
rect 165475 4996 165541 4997
rect 165475 4932 165476 4996
rect 165540 4932 165541 4996
rect 165475 4931 165541 4932
rect 163794 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 164414 -4186
rect 163794 -4506 164414 -4422
rect 163794 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 164414 -4506
rect 163794 -7654 164414 -4742
rect 168294 -5146 168914 25398
rect 169526 22813 169586 79459
rect 170262 77757 170322 79867
rect 170443 79524 170509 79525
rect 170443 79460 170444 79524
rect 170508 79460 170509 79524
rect 170443 79459 170509 79460
rect 170259 77756 170325 77757
rect 170259 77692 170260 77756
rect 170324 77692 170325 77756
rect 170259 77691 170325 77692
rect 170446 61437 170506 79459
rect 170443 61436 170509 61437
rect 170443 61372 170444 61436
rect 170508 61372 170509 61436
rect 170443 61371 170509 61372
rect 169523 22812 169589 22813
rect 169523 22748 169524 22812
rect 169588 22748 169589 22812
rect 169523 22747 169589 22748
rect 170630 22677 170690 80139
rect 171547 80068 171613 80069
rect 171547 80004 171548 80068
rect 171612 80004 171613 80068
rect 171547 80003 171613 80004
rect 170811 79796 170877 79797
rect 170811 79732 170812 79796
rect 170876 79732 170877 79796
rect 170811 79731 170877 79732
rect 170627 22676 170693 22677
rect 170627 22612 170628 22676
rect 170692 22612 170693 22676
rect 170627 22611 170693 22612
rect 170814 17373 170874 79731
rect 170995 78708 171061 78709
rect 170995 78644 170996 78708
rect 171060 78644 171061 78708
rect 170995 78643 171061 78644
rect 170811 17372 170877 17373
rect 170811 17308 170812 17372
rect 170876 17308 170877 17372
rect 170811 17307 170877 17308
rect 170998 11661 171058 78643
rect 171550 77310 171610 80003
rect 171731 79932 171797 79933
rect 171731 79868 171732 79932
rect 171796 79868 171797 79932
rect 171731 79867 171797 79868
rect 172651 79932 172717 79933
rect 172651 79868 172652 79932
rect 172716 79868 172717 79932
rect 172651 79867 172717 79868
rect 173203 79932 173269 79933
rect 173203 79868 173204 79932
rect 173268 79868 173269 79932
rect 173203 79867 173269 79868
rect 174675 79932 174741 79933
rect 174675 79868 174676 79932
rect 174740 79868 174741 79932
rect 174675 79867 174741 79868
rect 171734 78301 171794 79867
rect 172099 79660 172165 79661
rect 172099 79596 172100 79660
rect 172164 79596 172165 79660
rect 172099 79595 172165 79596
rect 171731 78300 171797 78301
rect 171731 78236 171732 78300
rect 171796 78236 171797 78300
rect 171731 78235 171797 78236
rect 172102 77754 172162 79595
rect 172654 78165 172714 79867
rect 173206 78165 173266 79867
rect 173387 79796 173453 79797
rect 173387 79732 173388 79796
rect 173452 79732 173453 79796
rect 173387 79731 173453 79732
rect 173390 78709 173450 79731
rect 173571 78980 173637 78981
rect 173571 78916 173572 78980
rect 173636 78916 173637 78980
rect 173571 78915 173637 78916
rect 173387 78708 173453 78709
rect 173387 78644 173388 78708
rect 173452 78644 173453 78708
rect 173387 78643 173453 78644
rect 172283 78164 172349 78165
rect 172283 78100 172284 78164
rect 172348 78100 172349 78164
rect 172283 78099 172349 78100
rect 172651 78164 172717 78165
rect 172651 78100 172652 78164
rect 172716 78100 172717 78164
rect 172651 78099 172717 78100
rect 173203 78164 173269 78165
rect 173203 78100 173204 78164
rect 173268 78100 173269 78164
rect 173203 78099 173269 78100
rect 171918 77694 172162 77754
rect 171550 77250 171794 77310
rect 171734 24173 171794 77250
rect 171918 65517 171978 77694
rect 172099 77484 172165 77485
rect 172099 77420 172100 77484
rect 172164 77420 172165 77484
rect 172099 77419 172165 77420
rect 171915 65516 171981 65517
rect 171915 65452 171916 65516
rect 171980 65452 171981 65516
rect 171915 65451 171981 65452
rect 172102 24309 172162 77419
rect 172286 75173 172346 78099
rect 172283 75172 172349 75173
rect 172283 75108 172284 75172
rect 172348 75108 172349 75172
rect 172283 75107 172349 75108
rect 172794 66454 173414 78000
rect 172794 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 173414 66454
rect 172794 66134 173414 66218
rect 172794 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 173414 66134
rect 172794 30454 173414 65898
rect 173574 64157 173634 78915
rect 173755 78708 173821 78709
rect 173755 78644 173756 78708
rect 173820 78644 173821 78708
rect 173755 78643 173821 78644
rect 173571 64156 173637 64157
rect 173571 64092 173572 64156
rect 173636 64092 173637 64156
rect 173571 64091 173637 64092
rect 173758 46205 173818 78643
rect 173755 46204 173821 46205
rect 173755 46140 173756 46204
rect 173820 46140 173821 46204
rect 173755 46139 173821 46140
rect 172794 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 173414 30454
rect 172794 30134 173414 30218
rect 172794 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 173414 30134
rect 172099 24308 172165 24309
rect 172099 24244 172100 24308
rect 172164 24244 172165 24308
rect 172099 24243 172165 24244
rect 171731 24172 171797 24173
rect 171731 24108 171732 24172
rect 171796 24108 171797 24172
rect 171731 24107 171797 24108
rect 170995 11660 171061 11661
rect 170995 11596 170996 11660
rect 171060 11596 171061 11660
rect 170995 11595 171061 11596
rect 168294 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 168914 -5146
rect 168294 -5466 168914 -5382
rect 168294 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 168914 -5466
rect 168294 -7654 168914 -5702
rect 172794 -6106 173414 29898
rect 174678 6221 174738 79867
rect 175230 79661 175290 80411
rect 176331 79932 176397 79933
rect 176331 79868 176332 79932
rect 176396 79868 176397 79932
rect 176331 79867 176397 79868
rect 176147 79796 176213 79797
rect 176147 79732 176148 79796
rect 176212 79732 176213 79796
rect 176147 79731 176213 79732
rect 175043 79660 175109 79661
rect 175043 79596 175044 79660
rect 175108 79596 175109 79660
rect 175043 79595 175109 79596
rect 175227 79660 175293 79661
rect 175227 79596 175228 79660
rect 175292 79596 175293 79660
rect 175227 79595 175293 79596
rect 174859 78708 174925 78709
rect 174859 78644 174860 78708
rect 174924 78644 174925 78708
rect 174859 78643 174925 78644
rect 174862 6357 174922 78643
rect 174859 6356 174925 6357
rect 174859 6292 174860 6356
rect 174924 6292 174925 6356
rect 174859 6291 174925 6292
rect 174675 6220 174741 6221
rect 174675 6156 174676 6220
rect 174740 6156 174741 6220
rect 174675 6155 174741 6156
rect 175046 4861 175106 79595
rect 176150 78981 176210 79731
rect 175227 78980 175293 78981
rect 175227 78916 175228 78980
rect 175292 78916 175293 78980
rect 175227 78915 175293 78916
rect 175779 78980 175845 78981
rect 175779 78916 175780 78980
rect 175844 78916 175845 78980
rect 175779 78915 175845 78916
rect 176147 78980 176213 78981
rect 176147 78916 176148 78980
rect 176212 78916 176213 78980
rect 176147 78915 176213 78916
rect 175230 71093 175290 78915
rect 175782 74493 175842 78915
rect 176147 78708 176213 78709
rect 176147 78644 176148 78708
rect 176212 78644 176213 78708
rect 176147 78643 176213 78644
rect 175779 74492 175845 74493
rect 175779 74428 175780 74492
rect 175844 74428 175845 74492
rect 175779 74427 175845 74428
rect 175227 71092 175293 71093
rect 175227 71028 175228 71092
rect 175292 71028 175293 71092
rect 175227 71027 175293 71028
rect 176150 66877 176210 78643
rect 176147 66876 176213 66877
rect 176147 66812 176148 66876
rect 176212 66812 176213 66876
rect 176147 66811 176213 66812
rect 176334 25533 176394 79867
rect 176702 79389 176762 80955
rect 176883 80884 176949 80885
rect 176883 80820 176884 80884
rect 176948 80820 176949 80884
rect 176883 80819 176949 80820
rect 176886 79797 176946 80819
rect 177435 80612 177501 80613
rect 177435 80548 177436 80612
rect 177500 80548 177501 80612
rect 177435 80547 177501 80548
rect 176883 79796 176949 79797
rect 176883 79732 176884 79796
rect 176948 79732 176949 79796
rect 176883 79731 176949 79732
rect 177438 79661 177498 80547
rect 177803 80204 177869 80205
rect 177803 80140 177804 80204
rect 177868 80140 177869 80204
rect 177803 80139 177869 80140
rect 177806 79933 177866 80139
rect 177803 79932 177869 79933
rect 177803 79868 177804 79932
rect 177868 79868 177869 79932
rect 177803 79867 177869 79868
rect 178355 79932 178421 79933
rect 178355 79868 178356 79932
rect 178420 79868 178421 79932
rect 178355 79867 178421 79868
rect 177435 79660 177501 79661
rect 177435 79596 177436 79660
rect 177500 79596 177501 79660
rect 177435 79595 177501 79596
rect 177067 79524 177133 79525
rect 177067 79460 177068 79524
rect 177132 79460 177133 79524
rect 177067 79459 177133 79460
rect 176699 79388 176765 79389
rect 176699 79324 176700 79388
rect 176764 79324 176765 79388
rect 176699 79323 176765 79324
rect 176515 78980 176581 78981
rect 176515 78916 176516 78980
rect 176580 78916 176581 78980
rect 176515 78915 176581 78916
rect 176331 25532 176397 25533
rect 176331 25468 176332 25532
rect 176396 25468 176397 25532
rect 176331 25467 176397 25468
rect 176518 17237 176578 78915
rect 176515 17236 176581 17237
rect 176515 17172 176516 17236
rect 176580 17172 176581 17236
rect 176515 17171 176581 17172
rect 175043 4860 175109 4861
rect 175043 4796 175044 4860
rect 175108 4796 175109 4860
rect 175043 4795 175109 4796
rect 177070 3365 177130 79459
rect 178358 79253 178418 79867
rect 178355 79252 178421 79253
rect 178355 79188 178356 79252
rect 178420 79188 178421 79252
rect 178355 79187 178421 79188
rect 177294 70954 177914 78000
rect 177294 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 177914 70954
rect 177294 70634 177914 70718
rect 177294 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 177914 70634
rect 177294 34954 177914 70398
rect 177294 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 177914 34954
rect 177294 34634 177914 34718
rect 177294 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 177914 34634
rect 177067 3364 177133 3365
rect 177067 3300 177068 3364
rect 177132 3300 177133 3364
rect 177067 3299 177133 3300
rect 172794 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 173414 -6106
rect 172794 -6426 173414 -6342
rect 172794 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 173414 -6426
rect 172794 -7654 173414 -6662
rect 177294 -7066 177914 34398
rect 177294 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 177914 -7066
rect 177294 -7386 177914 -7302
rect 177294 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 177914 -7386
rect 177294 -7654 177914 -7622
rect 181794 75454 182414 78000
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 186294 43954 186914 78000
rect 186294 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 186914 43954
rect 186294 43634 186914 43718
rect 186294 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 186914 43634
rect 186294 7954 186914 43398
rect 186294 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 186914 7954
rect 186294 7634 186914 7718
rect 186294 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 186914 7634
rect 186294 -1306 186914 7398
rect 186294 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 186914 -1306
rect 186294 -1626 186914 -1542
rect 186294 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 186914 -1626
rect 186294 -7654 186914 -1862
rect 190794 48454 191414 78000
rect 190794 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 191414 48454
rect 190794 48134 191414 48218
rect 190794 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 191414 48134
rect 190794 12454 191414 47898
rect 190794 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 191414 12454
rect 190794 12134 191414 12218
rect 190794 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 191414 12134
rect 190794 -2266 191414 11898
rect 190794 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 191414 -2266
rect 190794 -2586 191414 -2502
rect 190794 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 191414 -2586
rect 190794 -7654 191414 -2822
rect 195294 52954 195914 88398
rect 195294 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 195914 52954
rect 195294 52634 195914 52718
rect 195294 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 195914 52634
rect 195294 16954 195914 52398
rect 195294 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 195914 16954
rect 195294 16634 195914 16718
rect 195294 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 195914 16634
rect 195294 -3226 195914 16398
rect 195294 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 195914 -3226
rect 195294 -3546 195914 -3462
rect 195294 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 195914 -3546
rect 195294 -7654 195914 -3782
rect 199794 708678 200414 711590
rect 199794 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 200414 708678
rect 199794 708358 200414 708442
rect 199794 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 200414 708358
rect 199794 669454 200414 708122
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199794 237454 200414 272898
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -4186 200414 20898
rect 199794 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 200414 -4186
rect 199794 -4506 200414 -4422
rect 199794 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 200414 -4506
rect 199794 -7654 200414 -4742
rect 204294 709638 204914 711590
rect 204294 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 204914 709638
rect 204294 709318 204914 709402
rect 204294 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 204914 709318
rect 204294 673954 204914 709082
rect 204294 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 204914 673954
rect 204294 673634 204914 673718
rect 204294 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 204914 673634
rect 204294 637954 204914 673398
rect 204294 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 204914 637954
rect 204294 637634 204914 637718
rect 204294 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 204914 637634
rect 204294 601954 204914 637398
rect 204294 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 204914 601954
rect 204294 601634 204914 601718
rect 204294 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 204914 601634
rect 204294 565954 204914 601398
rect 204294 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 204914 565954
rect 204294 565634 204914 565718
rect 204294 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 204914 565634
rect 204294 529954 204914 565398
rect 204294 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 204914 529954
rect 204294 529634 204914 529718
rect 204294 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 204914 529634
rect 204294 493954 204914 529398
rect 204294 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 204914 493954
rect 204294 493634 204914 493718
rect 204294 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 204914 493634
rect 204294 457954 204914 493398
rect 204294 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 204914 457954
rect 204294 457634 204914 457718
rect 204294 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 204914 457634
rect 204294 421954 204914 457398
rect 204294 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 204914 421954
rect 204294 421634 204914 421718
rect 204294 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 204914 421634
rect 204294 385954 204914 421398
rect 204294 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 204914 385954
rect 204294 385634 204914 385718
rect 204294 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 204914 385634
rect 204294 349954 204914 385398
rect 204294 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 204914 349954
rect 204294 349634 204914 349718
rect 204294 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 204914 349634
rect 204294 313954 204914 349398
rect 204294 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 204914 313954
rect 204294 313634 204914 313718
rect 204294 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 204914 313634
rect 204294 277954 204914 313398
rect 204294 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 204914 277954
rect 204294 277634 204914 277718
rect 204294 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 204914 277634
rect 204294 241954 204914 277398
rect 204294 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 204914 241954
rect 204294 241634 204914 241718
rect 204294 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 204914 241634
rect 204294 205954 204914 241398
rect 204294 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 204914 205954
rect 204294 205634 204914 205718
rect 204294 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 204914 205634
rect 204294 169954 204914 205398
rect 204294 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 204914 169954
rect 204294 169634 204914 169718
rect 204294 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 204914 169634
rect 204294 133954 204914 169398
rect 204294 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 204914 133954
rect 204294 133634 204914 133718
rect 204294 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 204914 133634
rect 204294 97954 204914 133398
rect 204294 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 204914 97954
rect 204294 97634 204914 97718
rect 204294 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 204914 97634
rect 204294 61954 204914 97398
rect 204294 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 204914 61954
rect 204294 61634 204914 61718
rect 204294 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 204914 61634
rect 204294 25954 204914 61398
rect 204294 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 204914 25954
rect 204294 25634 204914 25718
rect 204294 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 204914 25634
rect 204294 -5146 204914 25398
rect 204294 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 204914 -5146
rect 204294 -5466 204914 -5382
rect 204294 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 204914 -5466
rect 204294 -7654 204914 -5702
rect 208794 710598 209414 711590
rect 208794 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 209414 710598
rect 208794 710278 209414 710362
rect 208794 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 209414 710278
rect 208794 678454 209414 710042
rect 208794 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 209414 678454
rect 208794 678134 209414 678218
rect 208794 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 209414 678134
rect 208794 642454 209414 677898
rect 208794 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 209414 642454
rect 208794 642134 209414 642218
rect 208794 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 209414 642134
rect 208794 606454 209414 641898
rect 208794 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 209414 606454
rect 208794 606134 209414 606218
rect 208794 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 209414 606134
rect 208794 570454 209414 605898
rect 208794 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 209414 570454
rect 208794 570134 209414 570218
rect 208794 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 209414 570134
rect 208794 534454 209414 569898
rect 208794 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 209414 534454
rect 208794 534134 209414 534218
rect 208794 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 209414 534134
rect 208794 498454 209414 533898
rect 208794 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 209414 498454
rect 208794 498134 209414 498218
rect 208794 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 209414 498134
rect 208794 462454 209414 497898
rect 208794 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 209414 462454
rect 208794 462134 209414 462218
rect 208794 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 209414 462134
rect 208794 426454 209414 461898
rect 208794 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 209414 426454
rect 208794 426134 209414 426218
rect 208794 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 209414 426134
rect 208794 390454 209414 425898
rect 208794 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 209414 390454
rect 208794 390134 209414 390218
rect 208794 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 209414 390134
rect 208794 354454 209414 389898
rect 208794 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 209414 354454
rect 208794 354134 209414 354218
rect 208794 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 209414 354134
rect 208794 318454 209414 353898
rect 208794 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 209414 318454
rect 208794 318134 209414 318218
rect 208794 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 209414 318134
rect 208794 282454 209414 317898
rect 208794 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 209414 282454
rect 208794 282134 209414 282218
rect 208794 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 209414 282134
rect 208794 246454 209414 281898
rect 208794 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 209414 246454
rect 208794 246134 209414 246218
rect 208794 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 209414 246134
rect 208794 210454 209414 245898
rect 208794 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 209414 210454
rect 208794 210134 209414 210218
rect 208794 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 209414 210134
rect 208794 174454 209414 209898
rect 208794 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 209414 174454
rect 208794 174134 209414 174218
rect 208794 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 209414 174134
rect 208794 138454 209414 173898
rect 208794 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 209414 138454
rect 208794 138134 209414 138218
rect 208794 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 209414 138134
rect 208794 102454 209414 137898
rect 208794 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 209414 102454
rect 208794 102134 209414 102218
rect 208794 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 209414 102134
rect 208794 66454 209414 101898
rect 208794 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 209414 66454
rect 208794 66134 209414 66218
rect 208794 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 209414 66134
rect 208794 30454 209414 65898
rect 208794 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 209414 30454
rect 208794 30134 209414 30218
rect 208794 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 209414 30134
rect 208794 -6106 209414 29898
rect 208794 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 209414 -6106
rect 208794 -6426 209414 -6342
rect 208794 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 209414 -6426
rect 208794 -7654 209414 -6662
rect 213294 711558 213914 711590
rect 213294 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 213914 711558
rect 213294 711238 213914 711322
rect 213294 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 213914 711238
rect 213294 682954 213914 711002
rect 213294 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 213914 682954
rect 213294 682634 213914 682718
rect 213294 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 213914 682634
rect 213294 646954 213914 682398
rect 213294 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 213914 646954
rect 213294 646634 213914 646718
rect 213294 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 213914 646634
rect 213294 610954 213914 646398
rect 213294 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 213914 610954
rect 213294 610634 213914 610718
rect 213294 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 213914 610634
rect 213294 574954 213914 610398
rect 213294 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 213914 574954
rect 213294 574634 213914 574718
rect 213294 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 213914 574634
rect 213294 538954 213914 574398
rect 213294 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 213914 538954
rect 213294 538634 213914 538718
rect 213294 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 213914 538634
rect 213294 502954 213914 538398
rect 213294 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 213914 502954
rect 213294 502634 213914 502718
rect 213294 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 213914 502634
rect 213294 466954 213914 502398
rect 213294 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 213914 466954
rect 213294 466634 213914 466718
rect 213294 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 213914 466634
rect 213294 430954 213914 466398
rect 213294 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 213914 430954
rect 213294 430634 213914 430718
rect 213294 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 213914 430634
rect 213294 394954 213914 430398
rect 213294 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 213914 394954
rect 213294 394634 213914 394718
rect 213294 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 213914 394634
rect 213294 358954 213914 394398
rect 213294 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 213914 358954
rect 213294 358634 213914 358718
rect 213294 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 213914 358634
rect 213294 322954 213914 358398
rect 213294 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 213914 322954
rect 213294 322634 213914 322718
rect 213294 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 213914 322634
rect 213294 286954 213914 322398
rect 213294 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 213914 286954
rect 213294 286634 213914 286718
rect 213294 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 213914 286634
rect 213294 250954 213914 286398
rect 213294 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 213914 250954
rect 213294 250634 213914 250718
rect 213294 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 213914 250634
rect 213294 214954 213914 250398
rect 213294 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 213914 214954
rect 213294 214634 213914 214718
rect 213294 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 213914 214634
rect 213294 178954 213914 214398
rect 213294 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 213914 178954
rect 213294 178634 213914 178718
rect 213294 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 213914 178634
rect 213294 142954 213914 178398
rect 213294 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 213914 142954
rect 213294 142634 213914 142718
rect 213294 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 213914 142634
rect 213294 106954 213914 142398
rect 213294 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 213914 106954
rect 213294 106634 213914 106718
rect 213294 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 213914 106634
rect 213294 70954 213914 106398
rect 213294 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 213914 70954
rect 213294 70634 213914 70718
rect 213294 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 213914 70634
rect 213294 34954 213914 70398
rect 213294 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 213914 34954
rect 213294 34634 213914 34718
rect 213294 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 213914 34634
rect 213294 -7066 213914 34398
rect 213294 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 213914 -7066
rect 213294 -7386 213914 -7302
rect 213294 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 213914 -7386
rect 213294 -7654 213914 -7622
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 219454 218414 254898
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 147454 218414 182898
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 222294 705798 222914 711590
rect 222294 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 222914 705798
rect 222294 705478 222914 705562
rect 222294 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 222914 705478
rect 222294 691954 222914 705242
rect 222294 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 222914 691954
rect 222294 691634 222914 691718
rect 222294 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 222914 691634
rect 222294 655954 222914 691398
rect 222294 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 222914 655954
rect 222294 655634 222914 655718
rect 222294 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 222914 655634
rect 222294 619954 222914 655398
rect 222294 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 222914 619954
rect 222294 619634 222914 619718
rect 222294 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 222914 619634
rect 222294 583954 222914 619398
rect 222294 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 222914 583954
rect 222294 583634 222914 583718
rect 222294 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 222914 583634
rect 222294 547954 222914 583398
rect 222294 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 222914 547954
rect 222294 547634 222914 547718
rect 222294 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 222914 547634
rect 222294 511954 222914 547398
rect 222294 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 222914 511954
rect 222294 511634 222914 511718
rect 222294 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 222914 511634
rect 222294 475954 222914 511398
rect 222294 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 222914 475954
rect 222294 475634 222914 475718
rect 222294 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 222914 475634
rect 222294 439954 222914 475398
rect 222294 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 222914 439954
rect 222294 439634 222914 439718
rect 222294 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 222914 439634
rect 222294 403954 222914 439398
rect 222294 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 222914 403954
rect 222294 403634 222914 403718
rect 222294 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 222914 403634
rect 222294 367954 222914 403398
rect 222294 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 222914 367954
rect 222294 367634 222914 367718
rect 222294 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 222914 367634
rect 222294 331954 222914 367398
rect 222294 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 222914 331954
rect 222294 331634 222914 331718
rect 222294 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 222914 331634
rect 222294 295954 222914 331398
rect 222294 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 222914 295954
rect 222294 295634 222914 295718
rect 222294 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 222914 295634
rect 222294 259954 222914 295398
rect 222294 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 222914 259954
rect 222294 259634 222914 259718
rect 222294 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 222914 259634
rect 222294 223954 222914 259398
rect 222294 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 222914 223954
rect 222294 223634 222914 223718
rect 222294 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 222914 223634
rect 222294 187954 222914 223398
rect 222294 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 222914 187954
rect 222294 187634 222914 187718
rect 222294 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 222914 187634
rect 222294 151954 222914 187398
rect 222294 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 222914 151954
rect 222294 151634 222914 151718
rect 222294 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 222914 151634
rect 222294 115954 222914 151398
rect 222294 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 222914 115954
rect 222294 115634 222914 115718
rect 222294 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 222914 115634
rect 222294 79954 222914 115398
rect 222294 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 222914 79954
rect 222294 79634 222914 79718
rect 222294 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 222914 79634
rect 222294 43954 222914 79398
rect 222294 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 222914 43954
rect 222294 43634 222914 43718
rect 222294 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 222914 43634
rect 222294 7954 222914 43398
rect 222294 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 222914 7954
rect 222294 7634 222914 7718
rect 222294 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 222914 7634
rect 222294 -1306 222914 7398
rect 222294 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 222914 -1306
rect 222294 -1626 222914 -1542
rect 222294 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 222914 -1626
rect 222294 -7654 222914 -1862
rect 226794 706758 227414 711590
rect 226794 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 227414 706758
rect 226794 706438 227414 706522
rect 226794 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 227414 706438
rect 226794 696454 227414 706202
rect 226794 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 227414 696454
rect 226794 696134 227414 696218
rect 226794 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 227414 696134
rect 226794 660454 227414 695898
rect 226794 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 227414 660454
rect 226794 660134 227414 660218
rect 226794 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 227414 660134
rect 226794 624454 227414 659898
rect 226794 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 227414 624454
rect 226794 624134 227414 624218
rect 226794 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 227414 624134
rect 226794 588454 227414 623898
rect 226794 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 227414 588454
rect 226794 588134 227414 588218
rect 226794 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 227414 588134
rect 226794 552454 227414 587898
rect 226794 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 227414 552454
rect 226794 552134 227414 552218
rect 226794 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 227414 552134
rect 226794 516454 227414 551898
rect 226794 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 227414 516454
rect 226794 516134 227414 516218
rect 226794 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 227414 516134
rect 226794 480454 227414 515898
rect 226794 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 227414 480454
rect 226794 480134 227414 480218
rect 226794 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 227414 480134
rect 226794 444454 227414 479898
rect 226794 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 227414 444454
rect 226794 444134 227414 444218
rect 226794 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 227414 444134
rect 226794 408454 227414 443898
rect 226794 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 227414 408454
rect 226794 408134 227414 408218
rect 226794 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 227414 408134
rect 226794 372454 227414 407898
rect 226794 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 227414 372454
rect 226794 372134 227414 372218
rect 226794 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 227414 372134
rect 226794 336454 227414 371898
rect 226794 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 227414 336454
rect 226794 336134 227414 336218
rect 226794 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 227414 336134
rect 226794 300454 227414 335898
rect 226794 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 227414 300454
rect 226794 300134 227414 300218
rect 226794 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 227414 300134
rect 226794 264454 227414 299898
rect 226794 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 227414 264454
rect 226794 264134 227414 264218
rect 226794 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 227414 264134
rect 226794 228454 227414 263898
rect 226794 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 227414 228454
rect 226794 228134 227414 228218
rect 226794 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 227414 228134
rect 226794 192454 227414 227898
rect 226794 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 227414 192454
rect 226794 192134 227414 192218
rect 226794 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 227414 192134
rect 226794 156454 227414 191898
rect 226794 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 227414 156454
rect 226794 156134 227414 156218
rect 226794 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 227414 156134
rect 226794 120454 227414 155898
rect 226794 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 227414 120454
rect 226794 120134 227414 120218
rect 226794 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 227414 120134
rect 226794 84454 227414 119898
rect 226794 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 227414 84454
rect 226794 84134 227414 84218
rect 226794 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 227414 84134
rect 226794 48454 227414 83898
rect 226794 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 227414 48454
rect 226794 48134 227414 48218
rect 226794 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 227414 48134
rect 226794 12454 227414 47898
rect 226794 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 227414 12454
rect 226794 12134 227414 12218
rect 226794 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 227414 12134
rect 226794 -2266 227414 11898
rect 226794 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 227414 -2266
rect 226794 -2586 227414 -2502
rect 226794 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 227414 -2586
rect 226794 -7654 227414 -2822
rect 231294 707718 231914 711590
rect 231294 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 231914 707718
rect 231294 707398 231914 707482
rect 231294 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 231914 707398
rect 231294 700954 231914 707162
rect 231294 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 231914 700954
rect 231294 700634 231914 700718
rect 231294 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 231914 700634
rect 231294 664954 231914 700398
rect 231294 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 231914 664954
rect 231294 664634 231914 664718
rect 231294 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 231914 664634
rect 231294 628954 231914 664398
rect 231294 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 231914 628954
rect 231294 628634 231914 628718
rect 231294 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 231914 628634
rect 231294 592954 231914 628398
rect 231294 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 231914 592954
rect 231294 592634 231914 592718
rect 231294 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 231914 592634
rect 231294 556954 231914 592398
rect 231294 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 231914 556954
rect 231294 556634 231914 556718
rect 231294 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 231914 556634
rect 231294 520954 231914 556398
rect 231294 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 231914 520954
rect 231294 520634 231914 520718
rect 231294 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 231914 520634
rect 231294 484954 231914 520398
rect 231294 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 231914 484954
rect 231294 484634 231914 484718
rect 231294 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 231914 484634
rect 231294 448954 231914 484398
rect 231294 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 231914 448954
rect 231294 448634 231914 448718
rect 231294 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 231914 448634
rect 231294 412954 231914 448398
rect 231294 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 231914 412954
rect 231294 412634 231914 412718
rect 231294 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 231914 412634
rect 231294 376954 231914 412398
rect 231294 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 231914 376954
rect 231294 376634 231914 376718
rect 231294 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 231914 376634
rect 231294 340954 231914 376398
rect 231294 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 231914 340954
rect 231294 340634 231914 340718
rect 231294 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 231914 340634
rect 231294 304954 231914 340398
rect 231294 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 231914 304954
rect 231294 304634 231914 304718
rect 231294 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 231914 304634
rect 231294 268954 231914 304398
rect 231294 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 231914 268954
rect 231294 268634 231914 268718
rect 231294 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 231914 268634
rect 231294 232954 231914 268398
rect 231294 232718 231326 232954
rect 231562 232718 231646 232954
rect 231882 232718 231914 232954
rect 231294 232634 231914 232718
rect 231294 232398 231326 232634
rect 231562 232398 231646 232634
rect 231882 232398 231914 232634
rect 231294 196954 231914 232398
rect 231294 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 231914 196954
rect 231294 196634 231914 196718
rect 231294 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 231914 196634
rect 231294 160954 231914 196398
rect 231294 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 231914 160954
rect 231294 160634 231914 160718
rect 231294 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 231914 160634
rect 231294 124954 231914 160398
rect 231294 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 231914 124954
rect 231294 124634 231914 124718
rect 231294 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 231914 124634
rect 231294 88954 231914 124398
rect 231294 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 231914 88954
rect 231294 88634 231914 88718
rect 231294 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 231914 88634
rect 231294 52954 231914 88398
rect 231294 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 231914 52954
rect 231294 52634 231914 52718
rect 231294 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 231914 52634
rect 231294 16954 231914 52398
rect 231294 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 231914 16954
rect 231294 16634 231914 16718
rect 231294 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 231914 16634
rect 231294 -3226 231914 16398
rect 231294 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 231914 -3226
rect 231294 -3546 231914 -3462
rect 231294 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 231914 -3546
rect 231294 -7654 231914 -3782
rect 235794 708678 236414 711590
rect 235794 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 236414 708678
rect 235794 708358 236414 708442
rect 235794 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 236414 708358
rect 235794 669454 236414 708122
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381454 236414 416898
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 273454 236414 308898
rect 235794 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 236414 273454
rect 235794 273134 236414 273218
rect 235794 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 236414 273134
rect 235794 237454 236414 272898
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 235794 201454 236414 236898
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 165454 236414 200898
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 235794 129454 236414 164898
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -4186 236414 20898
rect 235794 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 236414 -4186
rect 235794 -4506 236414 -4422
rect 235794 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 236414 -4506
rect 235794 -7654 236414 -4742
rect 240294 709638 240914 711590
rect 240294 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 240914 709638
rect 240294 709318 240914 709402
rect 240294 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 240914 709318
rect 240294 673954 240914 709082
rect 240294 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 240914 673954
rect 240294 673634 240914 673718
rect 240294 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 240914 673634
rect 240294 637954 240914 673398
rect 240294 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 240914 637954
rect 240294 637634 240914 637718
rect 240294 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 240914 637634
rect 240294 601954 240914 637398
rect 240294 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 240914 601954
rect 240294 601634 240914 601718
rect 240294 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 240914 601634
rect 240294 565954 240914 601398
rect 240294 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 240914 565954
rect 240294 565634 240914 565718
rect 240294 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 240914 565634
rect 240294 529954 240914 565398
rect 240294 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 240914 529954
rect 240294 529634 240914 529718
rect 240294 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 240914 529634
rect 240294 493954 240914 529398
rect 240294 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 240914 493954
rect 240294 493634 240914 493718
rect 240294 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 240914 493634
rect 240294 457954 240914 493398
rect 240294 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 240914 457954
rect 240294 457634 240914 457718
rect 240294 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 240914 457634
rect 240294 421954 240914 457398
rect 240294 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 240914 421954
rect 240294 421634 240914 421718
rect 240294 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 240914 421634
rect 240294 385954 240914 421398
rect 240294 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 240914 385954
rect 240294 385634 240914 385718
rect 240294 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 240914 385634
rect 240294 349954 240914 385398
rect 240294 349718 240326 349954
rect 240562 349718 240646 349954
rect 240882 349718 240914 349954
rect 240294 349634 240914 349718
rect 240294 349398 240326 349634
rect 240562 349398 240646 349634
rect 240882 349398 240914 349634
rect 240294 313954 240914 349398
rect 240294 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 240914 313954
rect 240294 313634 240914 313718
rect 240294 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 240914 313634
rect 240294 277954 240914 313398
rect 240294 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 240914 277954
rect 240294 277634 240914 277718
rect 240294 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 240914 277634
rect 240294 241954 240914 277398
rect 240294 241718 240326 241954
rect 240562 241718 240646 241954
rect 240882 241718 240914 241954
rect 240294 241634 240914 241718
rect 240294 241398 240326 241634
rect 240562 241398 240646 241634
rect 240882 241398 240914 241634
rect 240294 205954 240914 241398
rect 240294 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 240914 205954
rect 240294 205634 240914 205718
rect 240294 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 240914 205634
rect 240294 169954 240914 205398
rect 240294 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 240914 169954
rect 240294 169634 240914 169718
rect 240294 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 240914 169634
rect 240294 133954 240914 169398
rect 240294 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 240914 133954
rect 240294 133634 240914 133718
rect 240294 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 240914 133634
rect 240294 97954 240914 133398
rect 240294 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 240914 97954
rect 240294 97634 240914 97718
rect 240294 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 240914 97634
rect 240294 61954 240914 97398
rect 240294 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 240914 61954
rect 240294 61634 240914 61718
rect 240294 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 240914 61634
rect 240294 25954 240914 61398
rect 240294 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 240914 25954
rect 240294 25634 240914 25718
rect 240294 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 240914 25634
rect 240294 -5146 240914 25398
rect 240294 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 240914 -5146
rect 240294 -5466 240914 -5382
rect 240294 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 240914 -5466
rect 240294 -7654 240914 -5702
rect 244794 710598 245414 711590
rect 244794 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 245414 710598
rect 244794 710278 245414 710362
rect 244794 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 245414 710278
rect 244794 678454 245414 710042
rect 244794 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 245414 678454
rect 244794 678134 245414 678218
rect 244794 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 245414 678134
rect 244794 642454 245414 677898
rect 244794 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 245414 642454
rect 244794 642134 245414 642218
rect 244794 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 245414 642134
rect 244794 606454 245414 641898
rect 244794 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 245414 606454
rect 244794 606134 245414 606218
rect 244794 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 245414 606134
rect 244794 570454 245414 605898
rect 244794 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 245414 570454
rect 244794 570134 245414 570218
rect 244794 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 245414 570134
rect 244794 534454 245414 569898
rect 244794 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 245414 534454
rect 244794 534134 245414 534218
rect 244794 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 245414 534134
rect 244794 498454 245414 533898
rect 244794 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 245414 498454
rect 244794 498134 245414 498218
rect 244794 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 245414 498134
rect 244794 462454 245414 497898
rect 244794 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 245414 462454
rect 244794 462134 245414 462218
rect 244794 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 245414 462134
rect 244794 426454 245414 461898
rect 244794 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 245414 426454
rect 244794 426134 245414 426218
rect 244794 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 245414 426134
rect 244794 390454 245414 425898
rect 244794 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 245414 390454
rect 244794 390134 245414 390218
rect 244794 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 245414 390134
rect 244794 354454 245414 389898
rect 244794 354218 244826 354454
rect 245062 354218 245146 354454
rect 245382 354218 245414 354454
rect 244794 354134 245414 354218
rect 244794 353898 244826 354134
rect 245062 353898 245146 354134
rect 245382 353898 245414 354134
rect 244794 318454 245414 353898
rect 244794 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 245414 318454
rect 244794 318134 245414 318218
rect 244794 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 245414 318134
rect 244794 282454 245414 317898
rect 244794 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 245414 282454
rect 244794 282134 245414 282218
rect 244794 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 245414 282134
rect 244794 246454 245414 281898
rect 244794 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 245414 246454
rect 244794 246134 245414 246218
rect 244794 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 245414 246134
rect 244794 210454 245414 245898
rect 244794 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 245414 210454
rect 244794 210134 245414 210218
rect 244794 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 245414 210134
rect 244794 174454 245414 209898
rect 244794 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 245414 174454
rect 244794 174134 245414 174218
rect 244794 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 245414 174134
rect 244794 138454 245414 173898
rect 244794 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 245414 138454
rect 244794 138134 245414 138218
rect 244794 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 245414 138134
rect 244794 102454 245414 137898
rect 244794 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 245414 102454
rect 244794 102134 245414 102218
rect 244794 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 245414 102134
rect 244794 66454 245414 101898
rect 244794 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 245414 66454
rect 244794 66134 245414 66218
rect 244794 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 245414 66134
rect 244794 30454 245414 65898
rect 244794 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 245414 30454
rect 244794 30134 245414 30218
rect 244794 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 245414 30134
rect 244794 -6106 245414 29898
rect 244794 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 245414 -6106
rect 244794 -6426 245414 -6342
rect 244794 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 245414 -6426
rect 244794 -7654 245414 -6662
rect 249294 711558 249914 711590
rect 249294 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 249914 711558
rect 249294 711238 249914 711322
rect 249294 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 249914 711238
rect 249294 682954 249914 711002
rect 249294 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 249914 682954
rect 249294 682634 249914 682718
rect 249294 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 249914 682634
rect 249294 646954 249914 682398
rect 249294 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 249914 646954
rect 249294 646634 249914 646718
rect 249294 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 249914 646634
rect 249294 610954 249914 646398
rect 249294 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 249914 610954
rect 249294 610634 249914 610718
rect 249294 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 249914 610634
rect 249294 574954 249914 610398
rect 249294 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 249914 574954
rect 249294 574634 249914 574718
rect 249294 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 249914 574634
rect 249294 538954 249914 574398
rect 249294 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 249914 538954
rect 249294 538634 249914 538718
rect 249294 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 249914 538634
rect 249294 502954 249914 538398
rect 249294 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 249914 502954
rect 249294 502634 249914 502718
rect 249294 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 249914 502634
rect 249294 466954 249914 502398
rect 249294 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 249914 466954
rect 249294 466634 249914 466718
rect 249294 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 249914 466634
rect 249294 430954 249914 466398
rect 249294 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 249914 430954
rect 249294 430634 249914 430718
rect 249294 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 249914 430634
rect 249294 394954 249914 430398
rect 249294 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 249914 394954
rect 249294 394634 249914 394718
rect 249294 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 249914 394634
rect 249294 358954 249914 394398
rect 249294 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 249914 358954
rect 249294 358634 249914 358718
rect 249294 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 249914 358634
rect 249294 322954 249914 358398
rect 249294 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 249914 322954
rect 249294 322634 249914 322718
rect 249294 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 249914 322634
rect 249294 286954 249914 322398
rect 249294 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 249914 286954
rect 249294 286634 249914 286718
rect 249294 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 249914 286634
rect 249294 250954 249914 286398
rect 249294 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 249914 250954
rect 249294 250634 249914 250718
rect 249294 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 249914 250634
rect 249294 214954 249914 250398
rect 249294 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 249914 214954
rect 249294 214634 249914 214718
rect 249294 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 249914 214634
rect 249294 178954 249914 214398
rect 249294 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 249914 178954
rect 249294 178634 249914 178718
rect 249294 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 249914 178634
rect 249294 142954 249914 178398
rect 249294 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 249914 142954
rect 249294 142634 249914 142718
rect 249294 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 249914 142634
rect 249294 106954 249914 142398
rect 249294 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 249914 106954
rect 249294 106634 249914 106718
rect 249294 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 249914 106634
rect 249294 70954 249914 106398
rect 249294 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 249914 70954
rect 249294 70634 249914 70718
rect 249294 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 249914 70634
rect 249294 34954 249914 70398
rect 249294 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 249914 34954
rect 249294 34634 249914 34718
rect 249294 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 249914 34634
rect 249294 -7066 249914 34398
rect 249294 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 249914 -7066
rect 249294 -7386 249914 -7302
rect 249294 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 249914 -7386
rect 249294 -7654 249914 -7622
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 291454 254414 326898
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 219454 254414 254898
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 258294 705798 258914 711590
rect 258294 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 258914 705798
rect 258294 705478 258914 705562
rect 258294 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 258914 705478
rect 258294 691954 258914 705242
rect 258294 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 258914 691954
rect 258294 691634 258914 691718
rect 258294 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 258914 691634
rect 258294 655954 258914 691398
rect 258294 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 258914 655954
rect 258294 655634 258914 655718
rect 258294 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 258914 655634
rect 258294 619954 258914 655398
rect 258294 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 258914 619954
rect 258294 619634 258914 619718
rect 258294 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 258914 619634
rect 258294 583954 258914 619398
rect 258294 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 258914 583954
rect 258294 583634 258914 583718
rect 258294 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 258914 583634
rect 258294 547954 258914 583398
rect 258294 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 258914 547954
rect 258294 547634 258914 547718
rect 258294 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 258914 547634
rect 258294 511954 258914 547398
rect 258294 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 258914 511954
rect 258294 511634 258914 511718
rect 258294 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 258914 511634
rect 258294 475954 258914 511398
rect 258294 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 258914 475954
rect 258294 475634 258914 475718
rect 258294 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 258914 475634
rect 258294 439954 258914 475398
rect 258294 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 258914 439954
rect 258294 439634 258914 439718
rect 258294 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 258914 439634
rect 258294 403954 258914 439398
rect 258294 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 258914 403954
rect 258294 403634 258914 403718
rect 258294 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 258914 403634
rect 258294 367954 258914 403398
rect 258294 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 258914 367954
rect 258294 367634 258914 367718
rect 258294 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 258914 367634
rect 258294 331954 258914 367398
rect 258294 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 258914 331954
rect 258294 331634 258914 331718
rect 258294 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 258914 331634
rect 258294 295954 258914 331398
rect 258294 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 258914 295954
rect 258294 295634 258914 295718
rect 258294 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 258914 295634
rect 258294 259954 258914 295398
rect 258294 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 258914 259954
rect 258294 259634 258914 259718
rect 258294 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 258914 259634
rect 258294 223954 258914 259398
rect 258294 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 258914 223954
rect 258294 223634 258914 223718
rect 258294 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 258914 223634
rect 258294 187954 258914 223398
rect 258294 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 258914 187954
rect 258294 187634 258914 187718
rect 258294 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 258914 187634
rect 258294 151954 258914 187398
rect 258294 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 258914 151954
rect 258294 151634 258914 151718
rect 258294 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 258914 151634
rect 258294 115954 258914 151398
rect 258294 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 258914 115954
rect 258294 115634 258914 115718
rect 258294 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 258914 115634
rect 258294 79954 258914 115398
rect 258294 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 258914 79954
rect 258294 79634 258914 79718
rect 258294 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 258914 79634
rect 258294 43954 258914 79398
rect 258294 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 258914 43954
rect 258294 43634 258914 43718
rect 258294 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 258914 43634
rect 258294 7954 258914 43398
rect 258294 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 258914 7954
rect 258294 7634 258914 7718
rect 258294 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 258914 7634
rect 258294 -1306 258914 7398
rect 258294 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 258914 -1306
rect 258294 -1626 258914 -1542
rect 258294 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 258914 -1626
rect 258294 -7654 258914 -1862
rect 262794 706758 263414 711590
rect 262794 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 263414 706758
rect 262794 706438 263414 706522
rect 262794 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 263414 706438
rect 262794 696454 263414 706202
rect 262794 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 263414 696454
rect 262794 696134 263414 696218
rect 262794 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 263414 696134
rect 262794 660454 263414 695898
rect 262794 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 263414 660454
rect 262794 660134 263414 660218
rect 262794 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 263414 660134
rect 262794 624454 263414 659898
rect 262794 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 263414 624454
rect 262794 624134 263414 624218
rect 262794 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 263414 624134
rect 262794 588454 263414 623898
rect 262794 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 263414 588454
rect 262794 588134 263414 588218
rect 262794 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 263414 588134
rect 262794 552454 263414 587898
rect 262794 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 263414 552454
rect 262794 552134 263414 552218
rect 262794 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 263414 552134
rect 262794 516454 263414 551898
rect 262794 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 263414 516454
rect 262794 516134 263414 516218
rect 262794 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 263414 516134
rect 262794 480454 263414 515898
rect 262794 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 263414 480454
rect 262794 480134 263414 480218
rect 262794 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 263414 480134
rect 262794 444454 263414 479898
rect 262794 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 263414 444454
rect 262794 444134 263414 444218
rect 262794 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 263414 444134
rect 262794 408454 263414 443898
rect 262794 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 263414 408454
rect 262794 408134 263414 408218
rect 262794 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 263414 408134
rect 262794 372454 263414 407898
rect 262794 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 263414 372454
rect 262794 372134 263414 372218
rect 262794 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 263414 372134
rect 262794 336454 263414 371898
rect 262794 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 263414 336454
rect 262794 336134 263414 336218
rect 262794 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 263414 336134
rect 262794 300454 263414 335898
rect 262794 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 263414 300454
rect 262794 300134 263414 300218
rect 262794 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 263414 300134
rect 262794 264454 263414 299898
rect 262794 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 263414 264454
rect 262794 264134 263414 264218
rect 262794 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 263414 264134
rect 262794 228454 263414 263898
rect 262794 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 263414 228454
rect 262794 228134 263414 228218
rect 262794 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 263414 228134
rect 262794 192454 263414 227898
rect 262794 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 263414 192454
rect 262794 192134 263414 192218
rect 262794 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 263414 192134
rect 262794 156454 263414 191898
rect 262794 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 263414 156454
rect 262794 156134 263414 156218
rect 262794 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 263414 156134
rect 262794 120454 263414 155898
rect 262794 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 263414 120454
rect 262794 120134 263414 120218
rect 262794 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 263414 120134
rect 262794 84454 263414 119898
rect 262794 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 263414 84454
rect 262794 84134 263414 84218
rect 262794 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 263414 84134
rect 262794 48454 263414 83898
rect 262794 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 263414 48454
rect 262794 48134 263414 48218
rect 262794 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 263414 48134
rect 262794 12454 263414 47898
rect 262794 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 263414 12454
rect 262794 12134 263414 12218
rect 262794 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 263414 12134
rect 262794 -2266 263414 11898
rect 262794 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 263414 -2266
rect 262794 -2586 263414 -2502
rect 262794 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 263414 -2586
rect 262794 -7654 263414 -2822
rect 267294 707718 267914 711590
rect 267294 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 267914 707718
rect 267294 707398 267914 707482
rect 267294 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 267914 707398
rect 267294 700954 267914 707162
rect 267294 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 267914 700954
rect 267294 700634 267914 700718
rect 267294 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 267914 700634
rect 267294 664954 267914 700398
rect 267294 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 267914 664954
rect 267294 664634 267914 664718
rect 267294 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 267914 664634
rect 267294 628954 267914 664398
rect 267294 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 267914 628954
rect 267294 628634 267914 628718
rect 267294 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 267914 628634
rect 267294 592954 267914 628398
rect 267294 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 267914 592954
rect 267294 592634 267914 592718
rect 267294 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 267914 592634
rect 267294 556954 267914 592398
rect 267294 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 267914 556954
rect 267294 556634 267914 556718
rect 267294 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 267914 556634
rect 267294 520954 267914 556398
rect 267294 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 267914 520954
rect 267294 520634 267914 520718
rect 267294 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 267914 520634
rect 267294 484954 267914 520398
rect 267294 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 267914 484954
rect 267294 484634 267914 484718
rect 267294 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 267914 484634
rect 267294 448954 267914 484398
rect 267294 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 267914 448954
rect 267294 448634 267914 448718
rect 267294 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 267914 448634
rect 267294 412954 267914 448398
rect 267294 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 267914 412954
rect 267294 412634 267914 412718
rect 267294 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 267914 412634
rect 267294 376954 267914 412398
rect 267294 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 267914 376954
rect 267294 376634 267914 376718
rect 267294 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 267914 376634
rect 267294 340954 267914 376398
rect 267294 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 267914 340954
rect 267294 340634 267914 340718
rect 267294 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 267914 340634
rect 267294 304954 267914 340398
rect 267294 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 267914 304954
rect 267294 304634 267914 304718
rect 267294 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 267914 304634
rect 267294 268954 267914 304398
rect 267294 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 267914 268954
rect 267294 268634 267914 268718
rect 267294 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 267914 268634
rect 267294 232954 267914 268398
rect 267294 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 267914 232954
rect 267294 232634 267914 232718
rect 267294 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 267914 232634
rect 267294 196954 267914 232398
rect 267294 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 267914 196954
rect 267294 196634 267914 196718
rect 267294 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 267914 196634
rect 267294 160954 267914 196398
rect 267294 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 267914 160954
rect 267294 160634 267914 160718
rect 267294 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 267914 160634
rect 267294 124954 267914 160398
rect 267294 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 267914 124954
rect 267294 124634 267914 124718
rect 267294 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 267914 124634
rect 267294 88954 267914 124398
rect 267294 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 267914 88954
rect 267294 88634 267914 88718
rect 267294 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 267914 88634
rect 267294 52954 267914 88398
rect 267294 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 267914 52954
rect 267294 52634 267914 52718
rect 267294 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 267914 52634
rect 267294 16954 267914 52398
rect 267294 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 267914 16954
rect 267294 16634 267914 16718
rect 267294 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 267914 16634
rect 267294 -3226 267914 16398
rect 267294 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 267914 -3226
rect 267294 -3546 267914 -3462
rect 267294 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 267914 -3546
rect 267294 -7654 267914 -3782
rect 271794 708678 272414 711590
rect 271794 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 272414 708678
rect 271794 708358 272414 708442
rect 271794 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 272414 708358
rect 271794 669454 272414 708122
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 345454 272414 380898
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 273454 272414 308898
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 237454 272414 272898
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 271794 201454 272414 236898
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -4186 272414 20898
rect 271794 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 272414 -4186
rect 271794 -4506 272414 -4422
rect 271794 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 272414 -4506
rect 271794 -7654 272414 -4742
rect 276294 709638 276914 711590
rect 276294 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 276914 709638
rect 276294 709318 276914 709402
rect 276294 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 276914 709318
rect 276294 673954 276914 709082
rect 276294 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 276914 673954
rect 276294 673634 276914 673718
rect 276294 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 276914 673634
rect 276294 637954 276914 673398
rect 276294 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 276914 637954
rect 276294 637634 276914 637718
rect 276294 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 276914 637634
rect 276294 601954 276914 637398
rect 276294 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 276914 601954
rect 276294 601634 276914 601718
rect 276294 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 276914 601634
rect 276294 565954 276914 601398
rect 276294 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 276914 565954
rect 276294 565634 276914 565718
rect 276294 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 276914 565634
rect 276294 529954 276914 565398
rect 276294 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 276914 529954
rect 276294 529634 276914 529718
rect 276294 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 276914 529634
rect 276294 493954 276914 529398
rect 276294 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 276914 493954
rect 276294 493634 276914 493718
rect 276294 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 276914 493634
rect 276294 457954 276914 493398
rect 276294 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 276914 457954
rect 276294 457634 276914 457718
rect 276294 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 276914 457634
rect 276294 421954 276914 457398
rect 276294 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 276914 421954
rect 276294 421634 276914 421718
rect 276294 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 276914 421634
rect 276294 385954 276914 421398
rect 276294 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 276914 385954
rect 276294 385634 276914 385718
rect 276294 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 276914 385634
rect 276294 349954 276914 385398
rect 276294 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 276914 349954
rect 276294 349634 276914 349718
rect 276294 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 276914 349634
rect 276294 313954 276914 349398
rect 276294 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 276914 313954
rect 276294 313634 276914 313718
rect 276294 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 276914 313634
rect 276294 277954 276914 313398
rect 276294 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 276914 277954
rect 276294 277634 276914 277718
rect 276294 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 276914 277634
rect 276294 241954 276914 277398
rect 276294 241718 276326 241954
rect 276562 241718 276646 241954
rect 276882 241718 276914 241954
rect 276294 241634 276914 241718
rect 276294 241398 276326 241634
rect 276562 241398 276646 241634
rect 276882 241398 276914 241634
rect 276294 205954 276914 241398
rect 276294 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 276914 205954
rect 276294 205634 276914 205718
rect 276294 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 276914 205634
rect 276294 169954 276914 205398
rect 276294 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 276914 169954
rect 276294 169634 276914 169718
rect 276294 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 276914 169634
rect 276294 133954 276914 169398
rect 276294 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 276914 133954
rect 276294 133634 276914 133718
rect 276294 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 276914 133634
rect 276294 97954 276914 133398
rect 276294 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 276914 97954
rect 276294 97634 276914 97718
rect 276294 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 276914 97634
rect 276294 61954 276914 97398
rect 276294 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 276914 61954
rect 276294 61634 276914 61718
rect 276294 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 276914 61634
rect 276294 25954 276914 61398
rect 276294 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 276914 25954
rect 276294 25634 276914 25718
rect 276294 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 276914 25634
rect 276294 -5146 276914 25398
rect 276294 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 276914 -5146
rect 276294 -5466 276914 -5382
rect 276294 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 276914 -5466
rect 276294 -7654 276914 -5702
rect 280794 710598 281414 711590
rect 280794 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 281414 710598
rect 280794 710278 281414 710362
rect 280794 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 281414 710278
rect 280794 678454 281414 710042
rect 280794 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 281414 678454
rect 280794 678134 281414 678218
rect 280794 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 281414 678134
rect 280794 642454 281414 677898
rect 280794 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 281414 642454
rect 280794 642134 281414 642218
rect 280794 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 281414 642134
rect 280794 606454 281414 641898
rect 280794 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 281414 606454
rect 280794 606134 281414 606218
rect 280794 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 281414 606134
rect 280794 570454 281414 605898
rect 280794 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 281414 570454
rect 280794 570134 281414 570218
rect 280794 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 281414 570134
rect 280794 534454 281414 569898
rect 280794 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 281414 534454
rect 280794 534134 281414 534218
rect 280794 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 281414 534134
rect 280794 498454 281414 533898
rect 280794 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 281414 498454
rect 280794 498134 281414 498218
rect 280794 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 281414 498134
rect 280794 462454 281414 497898
rect 280794 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 281414 462454
rect 280794 462134 281414 462218
rect 280794 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 281414 462134
rect 280794 426454 281414 461898
rect 280794 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 281414 426454
rect 280794 426134 281414 426218
rect 280794 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 281414 426134
rect 280794 390454 281414 425898
rect 280794 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 281414 390454
rect 280794 390134 281414 390218
rect 280794 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 281414 390134
rect 280794 354454 281414 389898
rect 280794 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 281414 354454
rect 280794 354134 281414 354218
rect 280794 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 281414 354134
rect 280794 318454 281414 353898
rect 280794 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 281414 318454
rect 280794 318134 281414 318218
rect 280794 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 281414 318134
rect 280794 282454 281414 317898
rect 280794 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 281414 282454
rect 280794 282134 281414 282218
rect 280794 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 281414 282134
rect 280794 246454 281414 281898
rect 280794 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 281414 246454
rect 280794 246134 281414 246218
rect 280794 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 281414 246134
rect 280794 210454 281414 245898
rect 280794 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 281414 210454
rect 280794 210134 281414 210218
rect 280794 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 281414 210134
rect 280794 174454 281414 209898
rect 280794 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 281414 174454
rect 280794 174134 281414 174218
rect 280794 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 281414 174134
rect 280794 138454 281414 173898
rect 280794 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 281414 138454
rect 280794 138134 281414 138218
rect 280794 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 281414 138134
rect 280794 102454 281414 137898
rect 280794 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 281414 102454
rect 280794 102134 281414 102218
rect 280794 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 281414 102134
rect 280794 66454 281414 101898
rect 280794 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 281414 66454
rect 280794 66134 281414 66218
rect 280794 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 281414 66134
rect 280794 30454 281414 65898
rect 280794 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 281414 30454
rect 280794 30134 281414 30218
rect 280794 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 281414 30134
rect 280794 -6106 281414 29898
rect 280794 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 281414 -6106
rect 280794 -6426 281414 -6342
rect 280794 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 281414 -6426
rect 280794 -7654 281414 -6662
rect 285294 711558 285914 711590
rect 285294 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 285914 711558
rect 285294 711238 285914 711322
rect 285294 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 285914 711238
rect 285294 682954 285914 711002
rect 285294 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 285914 682954
rect 285294 682634 285914 682718
rect 285294 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 285914 682634
rect 285294 646954 285914 682398
rect 285294 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 285914 646954
rect 285294 646634 285914 646718
rect 285294 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 285914 646634
rect 285294 610954 285914 646398
rect 285294 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 285914 610954
rect 285294 610634 285914 610718
rect 285294 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 285914 610634
rect 285294 574954 285914 610398
rect 285294 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 285914 574954
rect 285294 574634 285914 574718
rect 285294 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 285914 574634
rect 285294 538954 285914 574398
rect 285294 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 285914 538954
rect 285294 538634 285914 538718
rect 285294 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 285914 538634
rect 285294 502954 285914 538398
rect 285294 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 285914 502954
rect 285294 502634 285914 502718
rect 285294 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 285914 502634
rect 285294 466954 285914 502398
rect 285294 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 285914 466954
rect 285294 466634 285914 466718
rect 285294 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 285914 466634
rect 285294 430954 285914 466398
rect 285294 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 285914 430954
rect 285294 430634 285914 430718
rect 285294 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 285914 430634
rect 285294 394954 285914 430398
rect 285294 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 285914 394954
rect 285294 394634 285914 394718
rect 285294 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 285914 394634
rect 285294 358954 285914 394398
rect 285294 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 285914 358954
rect 285294 358634 285914 358718
rect 285294 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 285914 358634
rect 285294 322954 285914 358398
rect 285294 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 285914 322954
rect 285294 322634 285914 322718
rect 285294 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 285914 322634
rect 285294 286954 285914 322398
rect 285294 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 285914 286954
rect 285294 286634 285914 286718
rect 285294 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 285914 286634
rect 285294 250954 285914 286398
rect 285294 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 285914 250954
rect 285294 250634 285914 250718
rect 285294 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 285914 250634
rect 285294 214954 285914 250398
rect 285294 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 285914 214954
rect 285294 214634 285914 214718
rect 285294 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 285914 214634
rect 285294 178954 285914 214398
rect 285294 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 285914 178954
rect 285294 178634 285914 178718
rect 285294 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 285914 178634
rect 285294 142954 285914 178398
rect 285294 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 285914 142954
rect 285294 142634 285914 142718
rect 285294 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 285914 142634
rect 285294 106954 285914 142398
rect 285294 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 285914 106954
rect 285294 106634 285914 106718
rect 285294 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 285914 106634
rect 285294 70954 285914 106398
rect 285294 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 285914 70954
rect 285294 70634 285914 70718
rect 285294 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 285914 70634
rect 285294 34954 285914 70398
rect 285294 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 285914 34954
rect 285294 34634 285914 34718
rect 285294 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 285914 34634
rect 285294 -7066 285914 34398
rect 285294 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 285914 -7066
rect 285294 -7386 285914 -7302
rect 285294 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 285914 -7386
rect 285294 -7654 285914 -7622
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 219454 290414 254898
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 294294 705798 294914 711590
rect 294294 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 294914 705798
rect 294294 705478 294914 705562
rect 294294 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 294914 705478
rect 294294 691954 294914 705242
rect 294294 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 294914 691954
rect 294294 691634 294914 691718
rect 294294 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 294914 691634
rect 294294 655954 294914 691398
rect 294294 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 294914 655954
rect 294294 655634 294914 655718
rect 294294 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 294914 655634
rect 294294 619954 294914 655398
rect 294294 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 294914 619954
rect 294294 619634 294914 619718
rect 294294 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 294914 619634
rect 294294 583954 294914 619398
rect 294294 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 294914 583954
rect 294294 583634 294914 583718
rect 294294 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 294914 583634
rect 294294 547954 294914 583398
rect 294294 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 294914 547954
rect 294294 547634 294914 547718
rect 294294 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 294914 547634
rect 294294 511954 294914 547398
rect 294294 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 294914 511954
rect 294294 511634 294914 511718
rect 294294 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 294914 511634
rect 294294 475954 294914 511398
rect 294294 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 294914 475954
rect 294294 475634 294914 475718
rect 294294 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 294914 475634
rect 294294 439954 294914 475398
rect 294294 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 294914 439954
rect 294294 439634 294914 439718
rect 294294 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 294914 439634
rect 294294 403954 294914 439398
rect 294294 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 294914 403954
rect 294294 403634 294914 403718
rect 294294 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 294914 403634
rect 294294 367954 294914 403398
rect 294294 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 294914 367954
rect 294294 367634 294914 367718
rect 294294 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 294914 367634
rect 294294 331954 294914 367398
rect 294294 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 294914 331954
rect 294294 331634 294914 331718
rect 294294 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 294914 331634
rect 294294 295954 294914 331398
rect 294294 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 294914 295954
rect 294294 295634 294914 295718
rect 294294 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 294914 295634
rect 294294 259954 294914 295398
rect 294294 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 294914 259954
rect 294294 259634 294914 259718
rect 294294 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 294914 259634
rect 294294 223954 294914 259398
rect 294294 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 294914 223954
rect 294294 223634 294914 223718
rect 294294 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 294914 223634
rect 294294 187954 294914 223398
rect 294294 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 294914 187954
rect 294294 187634 294914 187718
rect 294294 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 294914 187634
rect 294294 151954 294914 187398
rect 294294 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 294914 151954
rect 294294 151634 294914 151718
rect 294294 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 294914 151634
rect 294294 115954 294914 151398
rect 294294 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 294914 115954
rect 294294 115634 294914 115718
rect 294294 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 294914 115634
rect 294294 79954 294914 115398
rect 294294 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 294914 79954
rect 294294 79634 294914 79718
rect 294294 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 294914 79634
rect 294294 43954 294914 79398
rect 294294 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 294914 43954
rect 294294 43634 294914 43718
rect 294294 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 294914 43634
rect 294294 7954 294914 43398
rect 294294 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 294914 7954
rect 294294 7634 294914 7718
rect 294294 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 294914 7634
rect 294294 -1306 294914 7398
rect 294294 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 294914 -1306
rect 294294 -1626 294914 -1542
rect 294294 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 294914 -1626
rect 294294 -7654 294914 -1862
rect 298794 706758 299414 711590
rect 298794 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 299414 706758
rect 298794 706438 299414 706522
rect 298794 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 299414 706438
rect 298794 696454 299414 706202
rect 298794 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 299414 696454
rect 298794 696134 299414 696218
rect 298794 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 299414 696134
rect 298794 660454 299414 695898
rect 298794 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 299414 660454
rect 298794 660134 299414 660218
rect 298794 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 299414 660134
rect 298794 624454 299414 659898
rect 298794 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 299414 624454
rect 298794 624134 299414 624218
rect 298794 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 299414 624134
rect 298794 588454 299414 623898
rect 298794 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 299414 588454
rect 298794 588134 299414 588218
rect 298794 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 299414 588134
rect 298794 552454 299414 587898
rect 298794 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 299414 552454
rect 298794 552134 299414 552218
rect 298794 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 299414 552134
rect 298794 516454 299414 551898
rect 298794 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 299414 516454
rect 298794 516134 299414 516218
rect 298794 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 299414 516134
rect 298794 480454 299414 515898
rect 298794 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 299414 480454
rect 298794 480134 299414 480218
rect 298794 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 299414 480134
rect 298794 444454 299414 479898
rect 298794 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 299414 444454
rect 298794 444134 299414 444218
rect 298794 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 299414 444134
rect 298794 408454 299414 443898
rect 298794 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 299414 408454
rect 298794 408134 299414 408218
rect 298794 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 299414 408134
rect 298794 372454 299414 407898
rect 298794 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 299414 372454
rect 298794 372134 299414 372218
rect 298794 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 299414 372134
rect 298794 336454 299414 371898
rect 298794 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 299414 336454
rect 298794 336134 299414 336218
rect 298794 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 299414 336134
rect 298794 300454 299414 335898
rect 298794 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 299414 300454
rect 298794 300134 299414 300218
rect 298794 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 299414 300134
rect 298794 264454 299414 299898
rect 298794 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 299414 264454
rect 298794 264134 299414 264218
rect 298794 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 299414 264134
rect 298794 228454 299414 263898
rect 298794 228218 298826 228454
rect 299062 228218 299146 228454
rect 299382 228218 299414 228454
rect 298794 228134 299414 228218
rect 298794 227898 298826 228134
rect 299062 227898 299146 228134
rect 299382 227898 299414 228134
rect 298794 192454 299414 227898
rect 298794 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 299414 192454
rect 298794 192134 299414 192218
rect 298794 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 299414 192134
rect 298794 156454 299414 191898
rect 298794 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 299414 156454
rect 298794 156134 299414 156218
rect 298794 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 299414 156134
rect 298794 120454 299414 155898
rect 298794 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 299414 120454
rect 298794 120134 299414 120218
rect 298794 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 299414 120134
rect 298794 84454 299414 119898
rect 298794 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 299414 84454
rect 298794 84134 299414 84218
rect 298794 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 299414 84134
rect 298794 48454 299414 83898
rect 298794 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 299414 48454
rect 298794 48134 299414 48218
rect 298794 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 299414 48134
rect 298794 12454 299414 47898
rect 298794 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 299414 12454
rect 298794 12134 299414 12218
rect 298794 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 299414 12134
rect 298794 -2266 299414 11898
rect 298794 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 299414 -2266
rect 298794 -2586 299414 -2502
rect 298794 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 299414 -2586
rect 298794 -7654 299414 -2822
rect 303294 707718 303914 711590
rect 303294 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 303914 707718
rect 303294 707398 303914 707482
rect 303294 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 303914 707398
rect 303294 700954 303914 707162
rect 303294 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 303914 700954
rect 303294 700634 303914 700718
rect 303294 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 303914 700634
rect 303294 664954 303914 700398
rect 303294 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 303914 664954
rect 303294 664634 303914 664718
rect 303294 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 303914 664634
rect 303294 628954 303914 664398
rect 303294 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 303914 628954
rect 303294 628634 303914 628718
rect 303294 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 303914 628634
rect 303294 592954 303914 628398
rect 303294 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 303914 592954
rect 303294 592634 303914 592718
rect 303294 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 303914 592634
rect 303294 556954 303914 592398
rect 303294 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 303914 556954
rect 303294 556634 303914 556718
rect 303294 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 303914 556634
rect 303294 520954 303914 556398
rect 303294 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 303914 520954
rect 303294 520634 303914 520718
rect 303294 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 303914 520634
rect 303294 484954 303914 520398
rect 303294 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 303914 484954
rect 303294 484634 303914 484718
rect 303294 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 303914 484634
rect 303294 448954 303914 484398
rect 303294 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 303914 448954
rect 303294 448634 303914 448718
rect 303294 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 303914 448634
rect 303294 412954 303914 448398
rect 303294 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 303914 412954
rect 303294 412634 303914 412718
rect 303294 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 303914 412634
rect 303294 376954 303914 412398
rect 303294 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 303914 376954
rect 303294 376634 303914 376718
rect 303294 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 303914 376634
rect 303294 340954 303914 376398
rect 303294 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 303914 340954
rect 303294 340634 303914 340718
rect 303294 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 303914 340634
rect 303294 304954 303914 340398
rect 303294 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 303914 304954
rect 303294 304634 303914 304718
rect 303294 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 303914 304634
rect 303294 268954 303914 304398
rect 303294 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 303914 268954
rect 303294 268634 303914 268718
rect 303294 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 303914 268634
rect 303294 232954 303914 268398
rect 303294 232718 303326 232954
rect 303562 232718 303646 232954
rect 303882 232718 303914 232954
rect 303294 232634 303914 232718
rect 303294 232398 303326 232634
rect 303562 232398 303646 232634
rect 303882 232398 303914 232634
rect 303294 196954 303914 232398
rect 303294 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 303914 196954
rect 303294 196634 303914 196718
rect 303294 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 303914 196634
rect 303294 160954 303914 196398
rect 303294 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 303914 160954
rect 303294 160634 303914 160718
rect 303294 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 303914 160634
rect 303294 124954 303914 160398
rect 303294 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 303914 124954
rect 303294 124634 303914 124718
rect 303294 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 303914 124634
rect 303294 88954 303914 124398
rect 303294 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 303914 88954
rect 303294 88634 303914 88718
rect 303294 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 303914 88634
rect 303294 52954 303914 88398
rect 303294 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 303914 52954
rect 303294 52634 303914 52718
rect 303294 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 303914 52634
rect 303294 16954 303914 52398
rect 303294 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 303914 16954
rect 303294 16634 303914 16718
rect 303294 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 303914 16634
rect 303294 -3226 303914 16398
rect 303294 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 303914 -3226
rect 303294 -3546 303914 -3462
rect 303294 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 303914 -3546
rect 303294 -7654 303914 -3782
rect 307794 708678 308414 711590
rect 307794 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 308414 708678
rect 307794 708358 308414 708442
rect 307794 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 308414 708358
rect 307794 669454 308414 708122
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -4186 308414 20898
rect 307794 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 308414 -4186
rect 307794 -4506 308414 -4422
rect 307794 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 308414 -4506
rect 307794 -7654 308414 -4742
rect 312294 709638 312914 711590
rect 312294 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 312914 709638
rect 312294 709318 312914 709402
rect 312294 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 312914 709318
rect 312294 673954 312914 709082
rect 312294 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 312914 673954
rect 312294 673634 312914 673718
rect 312294 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 312914 673634
rect 312294 637954 312914 673398
rect 312294 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 312914 637954
rect 312294 637634 312914 637718
rect 312294 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 312914 637634
rect 312294 601954 312914 637398
rect 312294 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 312914 601954
rect 312294 601634 312914 601718
rect 312294 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 312914 601634
rect 312294 565954 312914 601398
rect 312294 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 312914 565954
rect 312294 565634 312914 565718
rect 312294 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 312914 565634
rect 312294 529954 312914 565398
rect 312294 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 312914 529954
rect 312294 529634 312914 529718
rect 312294 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 312914 529634
rect 312294 493954 312914 529398
rect 312294 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 312914 493954
rect 312294 493634 312914 493718
rect 312294 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 312914 493634
rect 312294 457954 312914 493398
rect 312294 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 312914 457954
rect 312294 457634 312914 457718
rect 312294 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 312914 457634
rect 312294 421954 312914 457398
rect 312294 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 312914 421954
rect 312294 421634 312914 421718
rect 312294 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 312914 421634
rect 312294 385954 312914 421398
rect 312294 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 312914 385954
rect 312294 385634 312914 385718
rect 312294 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 312914 385634
rect 312294 349954 312914 385398
rect 312294 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 312914 349954
rect 312294 349634 312914 349718
rect 312294 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 312914 349634
rect 312294 313954 312914 349398
rect 312294 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 312914 313954
rect 312294 313634 312914 313718
rect 312294 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 312914 313634
rect 312294 277954 312914 313398
rect 312294 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 312914 277954
rect 312294 277634 312914 277718
rect 312294 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 312914 277634
rect 312294 241954 312914 277398
rect 312294 241718 312326 241954
rect 312562 241718 312646 241954
rect 312882 241718 312914 241954
rect 312294 241634 312914 241718
rect 312294 241398 312326 241634
rect 312562 241398 312646 241634
rect 312882 241398 312914 241634
rect 312294 205954 312914 241398
rect 312294 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 312914 205954
rect 312294 205634 312914 205718
rect 312294 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 312914 205634
rect 312294 169954 312914 205398
rect 312294 169718 312326 169954
rect 312562 169718 312646 169954
rect 312882 169718 312914 169954
rect 312294 169634 312914 169718
rect 312294 169398 312326 169634
rect 312562 169398 312646 169634
rect 312882 169398 312914 169634
rect 312294 133954 312914 169398
rect 312294 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 312914 133954
rect 312294 133634 312914 133718
rect 312294 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 312914 133634
rect 312294 97954 312914 133398
rect 312294 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 312914 97954
rect 312294 97634 312914 97718
rect 312294 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 312914 97634
rect 312294 61954 312914 97398
rect 312294 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 312914 61954
rect 312294 61634 312914 61718
rect 312294 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 312914 61634
rect 312294 25954 312914 61398
rect 312294 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 312914 25954
rect 312294 25634 312914 25718
rect 312294 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 312914 25634
rect 312294 -5146 312914 25398
rect 312294 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 312914 -5146
rect 312294 -5466 312914 -5382
rect 312294 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 312914 -5466
rect 312294 -7654 312914 -5702
rect 316794 710598 317414 711590
rect 316794 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 317414 710598
rect 316794 710278 317414 710362
rect 316794 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 317414 710278
rect 316794 678454 317414 710042
rect 316794 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 317414 678454
rect 316794 678134 317414 678218
rect 316794 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 317414 678134
rect 316794 642454 317414 677898
rect 316794 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 317414 642454
rect 316794 642134 317414 642218
rect 316794 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 317414 642134
rect 316794 606454 317414 641898
rect 316794 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 317414 606454
rect 316794 606134 317414 606218
rect 316794 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 317414 606134
rect 316794 570454 317414 605898
rect 316794 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 317414 570454
rect 316794 570134 317414 570218
rect 316794 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 317414 570134
rect 316794 534454 317414 569898
rect 316794 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 317414 534454
rect 316794 534134 317414 534218
rect 316794 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 317414 534134
rect 316794 498454 317414 533898
rect 316794 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 317414 498454
rect 316794 498134 317414 498218
rect 316794 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 317414 498134
rect 316794 462454 317414 497898
rect 316794 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 317414 462454
rect 316794 462134 317414 462218
rect 316794 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 317414 462134
rect 316794 426454 317414 461898
rect 316794 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 317414 426454
rect 316794 426134 317414 426218
rect 316794 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 317414 426134
rect 316794 390454 317414 425898
rect 316794 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 317414 390454
rect 316794 390134 317414 390218
rect 316794 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 317414 390134
rect 316794 354454 317414 389898
rect 316794 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 317414 354454
rect 316794 354134 317414 354218
rect 316794 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 317414 354134
rect 316794 318454 317414 353898
rect 316794 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 317414 318454
rect 316794 318134 317414 318218
rect 316794 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 317414 318134
rect 316794 282454 317414 317898
rect 316794 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 317414 282454
rect 316794 282134 317414 282218
rect 316794 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 317414 282134
rect 316794 246454 317414 281898
rect 316794 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 317414 246454
rect 316794 246134 317414 246218
rect 316794 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 317414 246134
rect 316794 210454 317414 245898
rect 316794 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 317414 210454
rect 316794 210134 317414 210218
rect 316794 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 317414 210134
rect 316794 174454 317414 209898
rect 316794 174218 316826 174454
rect 317062 174218 317146 174454
rect 317382 174218 317414 174454
rect 316794 174134 317414 174218
rect 316794 173898 316826 174134
rect 317062 173898 317146 174134
rect 317382 173898 317414 174134
rect 316794 138454 317414 173898
rect 316794 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 317414 138454
rect 316794 138134 317414 138218
rect 316794 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 317414 138134
rect 316794 102454 317414 137898
rect 316794 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 317414 102454
rect 316794 102134 317414 102218
rect 316794 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 317414 102134
rect 316794 66454 317414 101898
rect 316794 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 317414 66454
rect 316794 66134 317414 66218
rect 316794 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 317414 66134
rect 316794 30454 317414 65898
rect 316794 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 317414 30454
rect 316794 30134 317414 30218
rect 316794 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 317414 30134
rect 316794 -6106 317414 29898
rect 316794 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 317414 -6106
rect 316794 -6426 317414 -6342
rect 316794 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 317414 -6426
rect 316794 -7654 317414 -6662
rect 321294 711558 321914 711590
rect 321294 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 321914 711558
rect 321294 711238 321914 711322
rect 321294 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 321914 711238
rect 321294 682954 321914 711002
rect 321294 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 321914 682954
rect 321294 682634 321914 682718
rect 321294 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 321914 682634
rect 321294 646954 321914 682398
rect 321294 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 321914 646954
rect 321294 646634 321914 646718
rect 321294 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 321914 646634
rect 321294 610954 321914 646398
rect 321294 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 321914 610954
rect 321294 610634 321914 610718
rect 321294 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 321914 610634
rect 321294 574954 321914 610398
rect 321294 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 321914 574954
rect 321294 574634 321914 574718
rect 321294 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 321914 574634
rect 321294 538954 321914 574398
rect 321294 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 321914 538954
rect 321294 538634 321914 538718
rect 321294 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 321914 538634
rect 321294 502954 321914 538398
rect 321294 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 321914 502954
rect 321294 502634 321914 502718
rect 321294 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 321914 502634
rect 321294 466954 321914 502398
rect 321294 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 321914 466954
rect 321294 466634 321914 466718
rect 321294 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 321914 466634
rect 321294 430954 321914 466398
rect 321294 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 321914 430954
rect 321294 430634 321914 430718
rect 321294 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 321914 430634
rect 321294 394954 321914 430398
rect 321294 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 321914 394954
rect 321294 394634 321914 394718
rect 321294 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 321914 394634
rect 321294 358954 321914 394398
rect 321294 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 321914 358954
rect 321294 358634 321914 358718
rect 321294 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 321914 358634
rect 321294 322954 321914 358398
rect 321294 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 321914 322954
rect 321294 322634 321914 322718
rect 321294 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 321914 322634
rect 321294 286954 321914 322398
rect 321294 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 321914 286954
rect 321294 286634 321914 286718
rect 321294 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 321914 286634
rect 321294 250954 321914 286398
rect 321294 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 321914 250954
rect 321294 250634 321914 250718
rect 321294 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 321914 250634
rect 321294 214954 321914 250398
rect 321294 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 321914 214954
rect 321294 214634 321914 214718
rect 321294 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 321914 214634
rect 321294 178954 321914 214398
rect 321294 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 321914 178954
rect 321294 178634 321914 178718
rect 321294 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 321914 178634
rect 321294 142954 321914 178398
rect 321294 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 321914 142954
rect 321294 142634 321914 142718
rect 321294 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 321914 142634
rect 321294 106954 321914 142398
rect 321294 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 321914 106954
rect 321294 106634 321914 106718
rect 321294 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 321914 106634
rect 321294 70954 321914 106398
rect 321294 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 321914 70954
rect 321294 70634 321914 70718
rect 321294 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 321914 70634
rect 321294 34954 321914 70398
rect 321294 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 321914 34954
rect 321294 34634 321914 34718
rect 321294 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 321914 34634
rect 321294 -7066 321914 34398
rect 321294 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 321914 -7066
rect 321294 -7386 321914 -7302
rect 321294 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 321914 -7386
rect 321294 -7654 321914 -7622
rect 325794 704838 326414 711590
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 330294 705798 330914 711590
rect 330294 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 330914 705798
rect 330294 705478 330914 705562
rect 330294 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 330914 705478
rect 330294 691954 330914 705242
rect 330294 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 330914 691954
rect 330294 691634 330914 691718
rect 330294 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 330914 691634
rect 330294 655954 330914 691398
rect 330294 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 330914 655954
rect 330294 655634 330914 655718
rect 330294 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 330914 655634
rect 330294 619954 330914 655398
rect 330294 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 330914 619954
rect 330294 619634 330914 619718
rect 330294 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 330914 619634
rect 330294 583954 330914 619398
rect 330294 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 330914 583954
rect 330294 583634 330914 583718
rect 330294 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 330914 583634
rect 330294 547954 330914 583398
rect 330294 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 330914 547954
rect 330294 547634 330914 547718
rect 330294 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 330914 547634
rect 330294 511954 330914 547398
rect 330294 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 330914 511954
rect 330294 511634 330914 511718
rect 330294 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 330914 511634
rect 330294 475954 330914 511398
rect 330294 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 330914 475954
rect 330294 475634 330914 475718
rect 330294 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 330914 475634
rect 330294 439954 330914 475398
rect 330294 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 330914 439954
rect 330294 439634 330914 439718
rect 330294 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 330914 439634
rect 330294 403954 330914 439398
rect 330294 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 330914 403954
rect 330294 403634 330914 403718
rect 330294 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 330914 403634
rect 330294 367954 330914 403398
rect 330294 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 330914 367954
rect 330294 367634 330914 367718
rect 330294 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 330914 367634
rect 330294 331954 330914 367398
rect 330294 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 330914 331954
rect 330294 331634 330914 331718
rect 330294 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 330914 331634
rect 330294 295954 330914 331398
rect 330294 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 330914 295954
rect 330294 295634 330914 295718
rect 330294 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 330914 295634
rect 330294 259954 330914 295398
rect 330294 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 330914 259954
rect 330294 259634 330914 259718
rect 330294 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 330914 259634
rect 330294 223954 330914 259398
rect 330294 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 330914 223954
rect 330294 223634 330914 223718
rect 330294 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 330914 223634
rect 330294 187954 330914 223398
rect 330294 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 330914 187954
rect 330294 187634 330914 187718
rect 330294 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 330914 187634
rect 330294 151954 330914 187398
rect 330294 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 330914 151954
rect 330294 151634 330914 151718
rect 330294 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 330914 151634
rect 330294 115954 330914 151398
rect 330294 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 330914 115954
rect 330294 115634 330914 115718
rect 330294 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 330914 115634
rect 330294 79954 330914 115398
rect 330294 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 330914 79954
rect 330294 79634 330914 79718
rect 330294 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 330914 79634
rect 330294 43954 330914 79398
rect 330294 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 330914 43954
rect 330294 43634 330914 43718
rect 330294 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 330914 43634
rect 330294 7954 330914 43398
rect 330294 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 330914 7954
rect 330294 7634 330914 7718
rect 330294 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 330914 7634
rect 330294 -1306 330914 7398
rect 330294 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 330914 -1306
rect 330294 -1626 330914 -1542
rect 330294 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 330914 -1626
rect 330294 -7654 330914 -1862
rect 334794 706758 335414 711590
rect 334794 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 335414 706758
rect 334794 706438 335414 706522
rect 334794 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 335414 706438
rect 334794 696454 335414 706202
rect 334794 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 335414 696454
rect 334794 696134 335414 696218
rect 334794 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 335414 696134
rect 334794 660454 335414 695898
rect 334794 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 335414 660454
rect 334794 660134 335414 660218
rect 334794 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 335414 660134
rect 334794 624454 335414 659898
rect 334794 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 335414 624454
rect 334794 624134 335414 624218
rect 334794 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 335414 624134
rect 334794 588454 335414 623898
rect 334794 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 335414 588454
rect 334794 588134 335414 588218
rect 334794 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 335414 588134
rect 334794 552454 335414 587898
rect 334794 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 335414 552454
rect 334794 552134 335414 552218
rect 334794 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 335414 552134
rect 334794 516454 335414 551898
rect 334794 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 335414 516454
rect 334794 516134 335414 516218
rect 334794 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 335414 516134
rect 334794 480454 335414 515898
rect 334794 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 335414 480454
rect 334794 480134 335414 480218
rect 334794 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 335414 480134
rect 334794 444454 335414 479898
rect 334794 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 335414 444454
rect 334794 444134 335414 444218
rect 334794 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 335414 444134
rect 334794 408454 335414 443898
rect 334794 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 335414 408454
rect 334794 408134 335414 408218
rect 334794 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 335414 408134
rect 334794 372454 335414 407898
rect 334794 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 335414 372454
rect 334794 372134 335414 372218
rect 334794 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 335414 372134
rect 334794 336454 335414 371898
rect 334794 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 335414 336454
rect 334794 336134 335414 336218
rect 334794 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 335414 336134
rect 334794 300454 335414 335898
rect 334794 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 335414 300454
rect 334794 300134 335414 300218
rect 334794 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 335414 300134
rect 334794 264454 335414 299898
rect 334794 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 335414 264454
rect 334794 264134 335414 264218
rect 334794 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 335414 264134
rect 334794 228454 335414 263898
rect 334794 228218 334826 228454
rect 335062 228218 335146 228454
rect 335382 228218 335414 228454
rect 334794 228134 335414 228218
rect 334794 227898 334826 228134
rect 335062 227898 335146 228134
rect 335382 227898 335414 228134
rect 334794 192454 335414 227898
rect 334794 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 335414 192454
rect 334794 192134 335414 192218
rect 334794 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 335414 192134
rect 334794 156454 335414 191898
rect 334794 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 335414 156454
rect 334794 156134 335414 156218
rect 334794 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 335414 156134
rect 334794 120454 335414 155898
rect 334794 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 335414 120454
rect 334794 120134 335414 120218
rect 334794 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 335414 120134
rect 334794 84454 335414 119898
rect 334794 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 335414 84454
rect 334794 84134 335414 84218
rect 334794 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 335414 84134
rect 334794 48454 335414 83898
rect 334794 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 335414 48454
rect 334794 48134 335414 48218
rect 334794 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 335414 48134
rect 334794 12454 335414 47898
rect 334794 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 335414 12454
rect 334794 12134 335414 12218
rect 334794 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 335414 12134
rect 334794 -2266 335414 11898
rect 334794 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 335414 -2266
rect 334794 -2586 335414 -2502
rect 334794 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 335414 -2586
rect 334794 -7654 335414 -2822
rect 339294 707718 339914 711590
rect 339294 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 339914 707718
rect 339294 707398 339914 707482
rect 339294 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 339914 707398
rect 339294 700954 339914 707162
rect 339294 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 339914 700954
rect 339294 700634 339914 700718
rect 339294 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 339914 700634
rect 339294 664954 339914 700398
rect 339294 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 339914 664954
rect 339294 664634 339914 664718
rect 339294 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 339914 664634
rect 339294 628954 339914 664398
rect 339294 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 339914 628954
rect 339294 628634 339914 628718
rect 339294 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 339914 628634
rect 339294 592954 339914 628398
rect 339294 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 339914 592954
rect 339294 592634 339914 592718
rect 339294 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 339914 592634
rect 339294 556954 339914 592398
rect 339294 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 339914 556954
rect 339294 556634 339914 556718
rect 339294 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 339914 556634
rect 339294 520954 339914 556398
rect 339294 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 339914 520954
rect 339294 520634 339914 520718
rect 339294 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 339914 520634
rect 339294 484954 339914 520398
rect 339294 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 339914 484954
rect 339294 484634 339914 484718
rect 339294 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 339914 484634
rect 339294 448954 339914 484398
rect 339294 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 339914 448954
rect 339294 448634 339914 448718
rect 339294 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 339914 448634
rect 339294 412954 339914 448398
rect 339294 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 339914 412954
rect 339294 412634 339914 412718
rect 339294 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 339914 412634
rect 339294 376954 339914 412398
rect 339294 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 339914 376954
rect 339294 376634 339914 376718
rect 339294 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 339914 376634
rect 339294 340954 339914 376398
rect 339294 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 339914 340954
rect 339294 340634 339914 340718
rect 339294 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 339914 340634
rect 339294 304954 339914 340398
rect 339294 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 339914 304954
rect 339294 304634 339914 304718
rect 339294 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 339914 304634
rect 339294 268954 339914 304398
rect 339294 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 339914 268954
rect 339294 268634 339914 268718
rect 339294 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 339914 268634
rect 339294 232954 339914 268398
rect 339294 232718 339326 232954
rect 339562 232718 339646 232954
rect 339882 232718 339914 232954
rect 339294 232634 339914 232718
rect 339294 232398 339326 232634
rect 339562 232398 339646 232634
rect 339882 232398 339914 232634
rect 339294 196954 339914 232398
rect 339294 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 339914 196954
rect 339294 196634 339914 196718
rect 339294 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 339914 196634
rect 339294 160954 339914 196398
rect 339294 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 339914 160954
rect 339294 160634 339914 160718
rect 339294 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 339914 160634
rect 339294 124954 339914 160398
rect 339294 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 339914 124954
rect 339294 124634 339914 124718
rect 339294 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 339914 124634
rect 339294 88954 339914 124398
rect 339294 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 339914 88954
rect 339294 88634 339914 88718
rect 339294 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 339914 88634
rect 339294 52954 339914 88398
rect 339294 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 339914 52954
rect 339294 52634 339914 52718
rect 339294 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 339914 52634
rect 339294 16954 339914 52398
rect 339294 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 339914 16954
rect 339294 16634 339914 16718
rect 339294 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 339914 16634
rect 339294 -3226 339914 16398
rect 339294 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 339914 -3226
rect 339294 -3546 339914 -3462
rect 339294 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 339914 -3546
rect 339294 -7654 339914 -3782
rect 343794 708678 344414 711590
rect 343794 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 344414 708678
rect 343794 708358 344414 708442
rect 343794 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 344414 708358
rect 343794 669454 344414 708122
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -4186 344414 20898
rect 343794 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 344414 -4186
rect 343794 -4506 344414 -4422
rect 343794 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 344414 -4506
rect 343794 -7654 344414 -4742
rect 348294 709638 348914 711590
rect 348294 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 348914 709638
rect 348294 709318 348914 709402
rect 348294 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 348914 709318
rect 348294 673954 348914 709082
rect 348294 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 348914 673954
rect 348294 673634 348914 673718
rect 348294 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 348914 673634
rect 348294 637954 348914 673398
rect 348294 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 348914 637954
rect 348294 637634 348914 637718
rect 348294 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 348914 637634
rect 348294 601954 348914 637398
rect 348294 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 348914 601954
rect 348294 601634 348914 601718
rect 348294 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 348914 601634
rect 348294 565954 348914 601398
rect 348294 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 348914 565954
rect 348294 565634 348914 565718
rect 348294 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 348914 565634
rect 348294 529954 348914 565398
rect 348294 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 348914 529954
rect 348294 529634 348914 529718
rect 348294 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 348914 529634
rect 348294 493954 348914 529398
rect 348294 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 348914 493954
rect 348294 493634 348914 493718
rect 348294 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 348914 493634
rect 348294 457954 348914 493398
rect 348294 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 348914 457954
rect 348294 457634 348914 457718
rect 348294 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 348914 457634
rect 348294 421954 348914 457398
rect 348294 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 348914 421954
rect 348294 421634 348914 421718
rect 348294 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 348914 421634
rect 348294 385954 348914 421398
rect 348294 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 348914 385954
rect 348294 385634 348914 385718
rect 348294 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 348914 385634
rect 348294 349954 348914 385398
rect 348294 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 348914 349954
rect 348294 349634 348914 349718
rect 348294 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 348914 349634
rect 348294 313954 348914 349398
rect 348294 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 348914 313954
rect 348294 313634 348914 313718
rect 348294 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 348914 313634
rect 348294 277954 348914 313398
rect 348294 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 348914 277954
rect 348294 277634 348914 277718
rect 348294 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 348914 277634
rect 348294 241954 348914 277398
rect 348294 241718 348326 241954
rect 348562 241718 348646 241954
rect 348882 241718 348914 241954
rect 348294 241634 348914 241718
rect 348294 241398 348326 241634
rect 348562 241398 348646 241634
rect 348882 241398 348914 241634
rect 348294 205954 348914 241398
rect 348294 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 348914 205954
rect 348294 205634 348914 205718
rect 348294 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 348914 205634
rect 348294 169954 348914 205398
rect 348294 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 348914 169954
rect 348294 169634 348914 169718
rect 348294 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 348914 169634
rect 348294 133954 348914 169398
rect 348294 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 348914 133954
rect 348294 133634 348914 133718
rect 348294 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 348914 133634
rect 348294 97954 348914 133398
rect 348294 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 348914 97954
rect 348294 97634 348914 97718
rect 348294 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 348914 97634
rect 348294 61954 348914 97398
rect 348294 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 348914 61954
rect 348294 61634 348914 61718
rect 348294 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 348914 61634
rect 348294 25954 348914 61398
rect 348294 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 348914 25954
rect 348294 25634 348914 25718
rect 348294 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 348914 25634
rect 348294 -5146 348914 25398
rect 348294 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 348914 -5146
rect 348294 -5466 348914 -5382
rect 348294 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 348914 -5466
rect 348294 -7654 348914 -5702
rect 352794 710598 353414 711590
rect 352794 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 353414 710598
rect 352794 710278 353414 710362
rect 352794 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 353414 710278
rect 352794 678454 353414 710042
rect 352794 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 353414 678454
rect 352794 678134 353414 678218
rect 352794 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 353414 678134
rect 352794 642454 353414 677898
rect 352794 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 353414 642454
rect 352794 642134 353414 642218
rect 352794 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 353414 642134
rect 352794 606454 353414 641898
rect 352794 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 353414 606454
rect 352794 606134 353414 606218
rect 352794 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 353414 606134
rect 352794 570454 353414 605898
rect 352794 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 353414 570454
rect 352794 570134 353414 570218
rect 352794 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 353414 570134
rect 352794 534454 353414 569898
rect 352794 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 353414 534454
rect 352794 534134 353414 534218
rect 352794 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 353414 534134
rect 352794 498454 353414 533898
rect 352794 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 353414 498454
rect 352794 498134 353414 498218
rect 352794 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 353414 498134
rect 352794 462454 353414 497898
rect 352794 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 353414 462454
rect 352794 462134 353414 462218
rect 352794 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 353414 462134
rect 352794 426454 353414 461898
rect 352794 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 353414 426454
rect 352794 426134 353414 426218
rect 352794 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 353414 426134
rect 352794 390454 353414 425898
rect 352794 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 353414 390454
rect 352794 390134 353414 390218
rect 352794 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 353414 390134
rect 352794 354454 353414 389898
rect 352794 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 353414 354454
rect 352794 354134 353414 354218
rect 352794 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 353414 354134
rect 352794 318454 353414 353898
rect 352794 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 353414 318454
rect 352794 318134 353414 318218
rect 352794 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 353414 318134
rect 352794 282454 353414 317898
rect 352794 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 353414 282454
rect 352794 282134 353414 282218
rect 352794 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 353414 282134
rect 352794 246454 353414 281898
rect 352794 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 353414 246454
rect 352794 246134 353414 246218
rect 352794 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 353414 246134
rect 352794 210454 353414 245898
rect 352794 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 353414 210454
rect 352794 210134 353414 210218
rect 352794 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 353414 210134
rect 352794 174454 353414 209898
rect 352794 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 353414 174454
rect 352794 174134 353414 174218
rect 352794 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 353414 174134
rect 352794 138454 353414 173898
rect 352794 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 353414 138454
rect 352794 138134 353414 138218
rect 352794 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 353414 138134
rect 352794 102454 353414 137898
rect 352794 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 353414 102454
rect 352794 102134 353414 102218
rect 352794 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 353414 102134
rect 352794 66454 353414 101898
rect 352794 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 353414 66454
rect 352794 66134 353414 66218
rect 352794 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 353414 66134
rect 352794 30454 353414 65898
rect 352794 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 353414 30454
rect 352794 30134 353414 30218
rect 352794 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 353414 30134
rect 352794 -6106 353414 29898
rect 352794 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 353414 -6106
rect 352794 -6426 353414 -6342
rect 352794 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 353414 -6426
rect 352794 -7654 353414 -6662
rect 357294 711558 357914 711590
rect 357294 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 357914 711558
rect 357294 711238 357914 711322
rect 357294 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 357914 711238
rect 357294 682954 357914 711002
rect 357294 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 357914 682954
rect 357294 682634 357914 682718
rect 357294 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 357914 682634
rect 357294 646954 357914 682398
rect 357294 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 357914 646954
rect 357294 646634 357914 646718
rect 357294 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 357914 646634
rect 357294 610954 357914 646398
rect 357294 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 357914 610954
rect 357294 610634 357914 610718
rect 357294 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 357914 610634
rect 357294 574954 357914 610398
rect 357294 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 357914 574954
rect 357294 574634 357914 574718
rect 357294 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 357914 574634
rect 357294 538954 357914 574398
rect 357294 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 357914 538954
rect 357294 538634 357914 538718
rect 357294 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 357914 538634
rect 357294 502954 357914 538398
rect 357294 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 357914 502954
rect 357294 502634 357914 502718
rect 357294 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 357914 502634
rect 357294 466954 357914 502398
rect 357294 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 357914 466954
rect 357294 466634 357914 466718
rect 357294 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 357914 466634
rect 357294 430954 357914 466398
rect 357294 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 357914 430954
rect 357294 430634 357914 430718
rect 357294 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 357914 430634
rect 357294 394954 357914 430398
rect 357294 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 357914 394954
rect 357294 394634 357914 394718
rect 357294 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 357914 394634
rect 357294 358954 357914 394398
rect 357294 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 357914 358954
rect 357294 358634 357914 358718
rect 357294 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 357914 358634
rect 357294 322954 357914 358398
rect 357294 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 357914 322954
rect 357294 322634 357914 322718
rect 357294 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 357914 322634
rect 357294 286954 357914 322398
rect 357294 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 357914 286954
rect 357294 286634 357914 286718
rect 357294 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 357914 286634
rect 357294 250954 357914 286398
rect 357294 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 357914 250954
rect 357294 250634 357914 250718
rect 357294 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 357914 250634
rect 357294 214954 357914 250398
rect 357294 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 357914 214954
rect 357294 214634 357914 214718
rect 357294 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 357914 214634
rect 357294 178954 357914 214398
rect 357294 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 357914 178954
rect 357294 178634 357914 178718
rect 357294 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 357914 178634
rect 357294 142954 357914 178398
rect 357294 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 357914 142954
rect 357294 142634 357914 142718
rect 357294 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 357914 142634
rect 357294 106954 357914 142398
rect 357294 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 357914 106954
rect 357294 106634 357914 106718
rect 357294 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 357914 106634
rect 357294 70954 357914 106398
rect 357294 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 357914 70954
rect 357294 70634 357914 70718
rect 357294 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 357914 70634
rect 357294 34954 357914 70398
rect 357294 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 357914 34954
rect 357294 34634 357914 34718
rect 357294 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 357914 34634
rect 357294 -7066 357914 34398
rect 357294 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 357914 -7066
rect 357294 -7386 357914 -7302
rect 357294 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 357914 -7386
rect 357294 -7654 357914 -7622
rect 361794 704838 362414 711590
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 366294 705798 366914 711590
rect 366294 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 366914 705798
rect 366294 705478 366914 705562
rect 366294 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 366914 705478
rect 366294 691954 366914 705242
rect 366294 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 366914 691954
rect 366294 691634 366914 691718
rect 366294 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 366914 691634
rect 366294 655954 366914 691398
rect 366294 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 366914 655954
rect 366294 655634 366914 655718
rect 366294 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 366914 655634
rect 366294 619954 366914 655398
rect 366294 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 366914 619954
rect 366294 619634 366914 619718
rect 366294 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 366914 619634
rect 366294 583954 366914 619398
rect 366294 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 366914 583954
rect 366294 583634 366914 583718
rect 366294 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 366914 583634
rect 366294 547954 366914 583398
rect 366294 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 366914 547954
rect 366294 547634 366914 547718
rect 366294 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 366914 547634
rect 366294 511954 366914 547398
rect 366294 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 366914 511954
rect 366294 511634 366914 511718
rect 366294 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 366914 511634
rect 366294 475954 366914 511398
rect 366294 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 366914 475954
rect 366294 475634 366914 475718
rect 366294 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 366914 475634
rect 366294 439954 366914 475398
rect 366294 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 366914 439954
rect 366294 439634 366914 439718
rect 366294 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 366914 439634
rect 366294 403954 366914 439398
rect 366294 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 366914 403954
rect 366294 403634 366914 403718
rect 366294 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 366914 403634
rect 366294 367954 366914 403398
rect 366294 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 366914 367954
rect 366294 367634 366914 367718
rect 366294 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 366914 367634
rect 366294 331954 366914 367398
rect 366294 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 366914 331954
rect 366294 331634 366914 331718
rect 366294 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 366914 331634
rect 366294 295954 366914 331398
rect 366294 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 366914 295954
rect 366294 295634 366914 295718
rect 366294 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 366914 295634
rect 366294 259954 366914 295398
rect 366294 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 366914 259954
rect 366294 259634 366914 259718
rect 366294 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 366914 259634
rect 366294 223954 366914 259398
rect 366294 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 366914 223954
rect 366294 223634 366914 223718
rect 366294 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 366914 223634
rect 366294 187954 366914 223398
rect 366294 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 366914 187954
rect 366294 187634 366914 187718
rect 366294 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 366914 187634
rect 366294 151954 366914 187398
rect 366294 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 366914 151954
rect 366294 151634 366914 151718
rect 366294 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 366914 151634
rect 366294 115954 366914 151398
rect 366294 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 366914 115954
rect 366294 115634 366914 115718
rect 366294 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 366914 115634
rect 366294 79954 366914 115398
rect 366294 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 366914 79954
rect 366294 79634 366914 79718
rect 366294 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 366914 79634
rect 366294 43954 366914 79398
rect 366294 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 366914 43954
rect 366294 43634 366914 43718
rect 366294 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 366914 43634
rect 366294 7954 366914 43398
rect 366294 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 366914 7954
rect 366294 7634 366914 7718
rect 366294 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 366914 7634
rect 366294 -1306 366914 7398
rect 366294 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 366914 -1306
rect 366294 -1626 366914 -1542
rect 366294 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 366914 -1626
rect 366294 -7654 366914 -1862
rect 370794 706758 371414 711590
rect 370794 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 371414 706758
rect 370794 706438 371414 706522
rect 370794 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 371414 706438
rect 370794 696454 371414 706202
rect 370794 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 371414 696454
rect 370794 696134 371414 696218
rect 370794 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 371414 696134
rect 370794 660454 371414 695898
rect 370794 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 371414 660454
rect 370794 660134 371414 660218
rect 370794 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 371414 660134
rect 370794 624454 371414 659898
rect 370794 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 371414 624454
rect 370794 624134 371414 624218
rect 370794 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 371414 624134
rect 370794 588454 371414 623898
rect 370794 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 371414 588454
rect 370794 588134 371414 588218
rect 370794 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 371414 588134
rect 370794 552454 371414 587898
rect 370794 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 371414 552454
rect 370794 552134 371414 552218
rect 370794 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 371414 552134
rect 370794 516454 371414 551898
rect 370794 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 371414 516454
rect 370794 516134 371414 516218
rect 370794 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 371414 516134
rect 370794 480454 371414 515898
rect 370794 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 371414 480454
rect 370794 480134 371414 480218
rect 370794 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 371414 480134
rect 370794 444454 371414 479898
rect 370794 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 371414 444454
rect 370794 444134 371414 444218
rect 370794 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 371414 444134
rect 370794 408454 371414 443898
rect 370794 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 371414 408454
rect 370794 408134 371414 408218
rect 370794 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 371414 408134
rect 370794 372454 371414 407898
rect 370794 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 371414 372454
rect 370794 372134 371414 372218
rect 370794 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 371414 372134
rect 370794 336454 371414 371898
rect 370794 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 371414 336454
rect 370794 336134 371414 336218
rect 370794 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 371414 336134
rect 370794 300454 371414 335898
rect 370794 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 371414 300454
rect 370794 300134 371414 300218
rect 370794 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 371414 300134
rect 370794 264454 371414 299898
rect 370794 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 371414 264454
rect 370794 264134 371414 264218
rect 370794 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 371414 264134
rect 370794 228454 371414 263898
rect 370794 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 371414 228454
rect 370794 228134 371414 228218
rect 370794 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 371414 228134
rect 370794 192454 371414 227898
rect 370794 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 371414 192454
rect 370794 192134 371414 192218
rect 370794 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 371414 192134
rect 370794 156454 371414 191898
rect 370794 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 371414 156454
rect 370794 156134 371414 156218
rect 370794 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 371414 156134
rect 370794 120454 371414 155898
rect 370794 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 371414 120454
rect 370794 120134 371414 120218
rect 370794 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 371414 120134
rect 370794 84454 371414 119898
rect 370794 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 371414 84454
rect 370794 84134 371414 84218
rect 370794 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 371414 84134
rect 370794 48454 371414 83898
rect 370794 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 371414 48454
rect 370794 48134 371414 48218
rect 370794 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 371414 48134
rect 370794 12454 371414 47898
rect 370794 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 371414 12454
rect 370794 12134 371414 12218
rect 370794 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 371414 12134
rect 370794 -2266 371414 11898
rect 370794 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 371414 -2266
rect 370794 -2586 371414 -2502
rect 370794 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 371414 -2586
rect 370794 -7654 371414 -2822
rect 375294 707718 375914 711590
rect 375294 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 375914 707718
rect 375294 707398 375914 707482
rect 375294 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 375914 707398
rect 375294 700954 375914 707162
rect 375294 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 375914 700954
rect 375294 700634 375914 700718
rect 375294 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 375914 700634
rect 375294 664954 375914 700398
rect 375294 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 375914 664954
rect 375294 664634 375914 664718
rect 375294 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 375914 664634
rect 375294 628954 375914 664398
rect 375294 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 375914 628954
rect 375294 628634 375914 628718
rect 375294 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 375914 628634
rect 375294 592954 375914 628398
rect 375294 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 375914 592954
rect 375294 592634 375914 592718
rect 375294 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 375914 592634
rect 375294 556954 375914 592398
rect 375294 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 375914 556954
rect 375294 556634 375914 556718
rect 375294 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 375914 556634
rect 375294 520954 375914 556398
rect 375294 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 375914 520954
rect 375294 520634 375914 520718
rect 375294 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 375914 520634
rect 375294 484954 375914 520398
rect 375294 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 375914 484954
rect 375294 484634 375914 484718
rect 375294 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 375914 484634
rect 375294 448954 375914 484398
rect 375294 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 375914 448954
rect 375294 448634 375914 448718
rect 375294 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 375914 448634
rect 375294 412954 375914 448398
rect 375294 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 375914 412954
rect 375294 412634 375914 412718
rect 375294 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 375914 412634
rect 375294 376954 375914 412398
rect 375294 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 375914 376954
rect 375294 376634 375914 376718
rect 375294 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 375914 376634
rect 375294 340954 375914 376398
rect 375294 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 375914 340954
rect 375294 340634 375914 340718
rect 375294 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 375914 340634
rect 375294 304954 375914 340398
rect 375294 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 375914 304954
rect 375294 304634 375914 304718
rect 375294 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 375914 304634
rect 375294 268954 375914 304398
rect 375294 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 375914 268954
rect 375294 268634 375914 268718
rect 375294 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 375914 268634
rect 375294 232954 375914 268398
rect 375294 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 375914 232954
rect 375294 232634 375914 232718
rect 375294 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 375914 232634
rect 375294 196954 375914 232398
rect 375294 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 375914 196954
rect 375294 196634 375914 196718
rect 375294 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 375914 196634
rect 375294 160954 375914 196398
rect 375294 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 375914 160954
rect 375294 160634 375914 160718
rect 375294 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 375914 160634
rect 375294 124954 375914 160398
rect 375294 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 375914 124954
rect 375294 124634 375914 124718
rect 375294 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 375914 124634
rect 375294 88954 375914 124398
rect 375294 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 375914 88954
rect 375294 88634 375914 88718
rect 375294 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 375914 88634
rect 375294 52954 375914 88398
rect 375294 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 375914 52954
rect 375294 52634 375914 52718
rect 375294 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 375914 52634
rect 375294 16954 375914 52398
rect 375294 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 375914 16954
rect 375294 16634 375914 16718
rect 375294 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 375914 16634
rect 375294 -3226 375914 16398
rect 375294 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 375914 -3226
rect 375294 -3546 375914 -3462
rect 375294 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 375914 -3546
rect 375294 -7654 375914 -3782
rect 379794 708678 380414 711590
rect 379794 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 380414 708678
rect 379794 708358 380414 708442
rect 379794 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 380414 708358
rect 379794 669454 380414 708122
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -4186 380414 20898
rect 379794 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 380414 -4186
rect 379794 -4506 380414 -4422
rect 379794 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 380414 -4506
rect 379794 -7654 380414 -4742
rect 384294 709638 384914 711590
rect 384294 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 384914 709638
rect 384294 709318 384914 709402
rect 384294 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 384914 709318
rect 384294 673954 384914 709082
rect 384294 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 384914 673954
rect 384294 673634 384914 673718
rect 384294 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 384914 673634
rect 384294 637954 384914 673398
rect 384294 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 384914 637954
rect 384294 637634 384914 637718
rect 384294 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 384914 637634
rect 384294 601954 384914 637398
rect 384294 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 384914 601954
rect 384294 601634 384914 601718
rect 384294 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 384914 601634
rect 384294 565954 384914 601398
rect 384294 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 384914 565954
rect 384294 565634 384914 565718
rect 384294 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 384914 565634
rect 384294 529954 384914 565398
rect 384294 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 384914 529954
rect 384294 529634 384914 529718
rect 384294 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 384914 529634
rect 384294 493954 384914 529398
rect 384294 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 384914 493954
rect 384294 493634 384914 493718
rect 384294 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 384914 493634
rect 384294 457954 384914 493398
rect 384294 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 384914 457954
rect 384294 457634 384914 457718
rect 384294 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 384914 457634
rect 384294 421954 384914 457398
rect 384294 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 384914 421954
rect 384294 421634 384914 421718
rect 384294 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 384914 421634
rect 384294 385954 384914 421398
rect 384294 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 384914 385954
rect 384294 385634 384914 385718
rect 384294 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 384914 385634
rect 384294 349954 384914 385398
rect 384294 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 384914 349954
rect 384294 349634 384914 349718
rect 384294 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 384914 349634
rect 384294 313954 384914 349398
rect 384294 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 384914 313954
rect 384294 313634 384914 313718
rect 384294 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 384914 313634
rect 384294 277954 384914 313398
rect 384294 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 384914 277954
rect 384294 277634 384914 277718
rect 384294 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 384914 277634
rect 384294 241954 384914 277398
rect 384294 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 384914 241954
rect 384294 241634 384914 241718
rect 384294 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 384914 241634
rect 384294 205954 384914 241398
rect 384294 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 384914 205954
rect 384294 205634 384914 205718
rect 384294 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 384914 205634
rect 384294 169954 384914 205398
rect 384294 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 384914 169954
rect 384294 169634 384914 169718
rect 384294 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 384914 169634
rect 384294 133954 384914 169398
rect 384294 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 384914 133954
rect 384294 133634 384914 133718
rect 384294 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 384914 133634
rect 384294 97954 384914 133398
rect 384294 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 384914 97954
rect 384294 97634 384914 97718
rect 384294 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 384914 97634
rect 384294 61954 384914 97398
rect 384294 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 384914 61954
rect 384294 61634 384914 61718
rect 384294 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 384914 61634
rect 384294 25954 384914 61398
rect 384294 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 384914 25954
rect 384294 25634 384914 25718
rect 384294 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 384914 25634
rect 384294 -5146 384914 25398
rect 384294 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 384914 -5146
rect 384294 -5466 384914 -5382
rect 384294 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 384914 -5466
rect 384294 -7654 384914 -5702
rect 388794 710598 389414 711590
rect 388794 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 389414 710598
rect 388794 710278 389414 710362
rect 388794 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 389414 710278
rect 388794 678454 389414 710042
rect 388794 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 389414 678454
rect 388794 678134 389414 678218
rect 388794 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 389414 678134
rect 388794 642454 389414 677898
rect 388794 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 389414 642454
rect 388794 642134 389414 642218
rect 388794 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 389414 642134
rect 388794 606454 389414 641898
rect 388794 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 389414 606454
rect 388794 606134 389414 606218
rect 388794 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 389414 606134
rect 388794 570454 389414 605898
rect 388794 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 389414 570454
rect 388794 570134 389414 570218
rect 388794 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 389414 570134
rect 388794 534454 389414 569898
rect 388794 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 389414 534454
rect 388794 534134 389414 534218
rect 388794 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 389414 534134
rect 388794 498454 389414 533898
rect 388794 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 389414 498454
rect 388794 498134 389414 498218
rect 388794 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 389414 498134
rect 388794 462454 389414 497898
rect 388794 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 389414 462454
rect 388794 462134 389414 462218
rect 388794 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 389414 462134
rect 388794 426454 389414 461898
rect 388794 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 389414 426454
rect 388794 426134 389414 426218
rect 388794 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 389414 426134
rect 388794 390454 389414 425898
rect 388794 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 389414 390454
rect 388794 390134 389414 390218
rect 388794 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 389414 390134
rect 388794 354454 389414 389898
rect 388794 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 389414 354454
rect 388794 354134 389414 354218
rect 388794 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 389414 354134
rect 388794 318454 389414 353898
rect 388794 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 389414 318454
rect 388794 318134 389414 318218
rect 388794 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 389414 318134
rect 388794 282454 389414 317898
rect 388794 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 389414 282454
rect 388794 282134 389414 282218
rect 388794 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 389414 282134
rect 388794 246454 389414 281898
rect 388794 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 389414 246454
rect 388794 246134 389414 246218
rect 388794 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 389414 246134
rect 388794 210454 389414 245898
rect 388794 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 389414 210454
rect 388794 210134 389414 210218
rect 388794 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 389414 210134
rect 388794 174454 389414 209898
rect 388794 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 389414 174454
rect 388794 174134 389414 174218
rect 388794 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 389414 174134
rect 388794 138454 389414 173898
rect 388794 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 389414 138454
rect 388794 138134 389414 138218
rect 388794 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 389414 138134
rect 388794 102454 389414 137898
rect 388794 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 389414 102454
rect 388794 102134 389414 102218
rect 388794 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 389414 102134
rect 388794 66454 389414 101898
rect 388794 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 389414 66454
rect 388794 66134 389414 66218
rect 388794 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 389414 66134
rect 388794 30454 389414 65898
rect 388794 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 389414 30454
rect 388794 30134 389414 30218
rect 388794 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 389414 30134
rect 388794 -6106 389414 29898
rect 388794 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 389414 -6106
rect 388794 -6426 389414 -6342
rect 388794 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 389414 -6426
rect 388794 -7654 389414 -6662
rect 393294 711558 393914 711590
rect 393294 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 393914 711558
rect 393294 711238 393914 711322
rect 393294 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 393914 711238
rect 393294 682954 393914 711002
rect 393294 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 393914 682954
rect 393294 682634 393914 682718
rect 393294 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 393914 682634
rect 393294 646954 393914 682398
rect 393294 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 393914 646954
rect 393294 646634 393914 646718
rect 393294 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 393914 646634
rect 393294 610954 393914 646398
rect 393294 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 393914 610954
rect 393294 610634 393914 610718
rect 393294 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 393914 610634
rect 393294 574954 393914 610398
rect 393294 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 393914 574954
rect 393294 574634 393914 574718
rect 393294 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 393914 574634
rect 393294 538954 393914 574398
rect 393294 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 393914 538954
rect 393294 538634 393914 538718
rect 393294 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 393914 538634
rect 393294 502954 393914 538398
rect 393294 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 393914 502954
rect 393294 502634 393914 502718
rect 393294 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 393914 502634
rect 393294 466954 393914 502398
rect 393294 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 393914 466954
rect 393294 466634 393914 466718
rect 393294 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 393914 466634
rect 393294 430954 393914 466398
rect 393294 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 393914 430954
rect 393294 430634 393914 430718
rect 393294 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 393914 430634
rect 393294 394954 393914 430398
rect 393294 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 393914 394954
rect 393294 394634 393914 394718
rect 393294 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 393914 394634
rect 393294 358954 393914 394398
rect 393294 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 393914 358954
rect 393294 358634 393914 358718
rect 393294 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 393914 358634
rect 393294 322954 393914 358398
rect 393294 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 393914 322954
rect 393294 322634 393914 322718
rect 393294 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 393914 322634
rect 393294 286954 393914 322398
rect 393294 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 393914 286954
rect 393294 286634 393914 286718
rect 393294 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 393914 286634
rect 393294 250954 393914 286398
rect 393294 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 393914 250954
rect 393294 250634 393914 250718
rect 393294 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 393914 250634
rect 393294 214954 393914 250398
rect 393294 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 393914 214954
rect 393294 214634 393914 214718
rect 393294 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 393914 214634
rect 393294 178954 393914 214398
rect 393294 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 393914 178954
rect 393294 178634 393914 178718
rect 393294 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 393914 178634
rect 393294 142954 393914 178398
rect 393294 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 393914 142954
rect 393294 142634 393914 142718
rect 393294 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 393914 142634
rect 393294 106954 393914 142398
rect 393294 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 393914 106954
rect 393294 106634 393914 106718
rect 393294 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 393914 106634
rect 393294 70954 393914 106398
rect 393294 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 393914 70954
rect 393294 70634 393914 70718
rect 393294 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 393914 70634
rect 393294 34954 393914 70398
rect 393294 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 393914 34954
rect 393294 34634 393914 34718
rect 393294 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 393914 34634
rect 393294 -7066 393914 34398
rect 393294 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 393914 -7066
rect 393294 -7386 393914 -7302
rect 393294 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 393914 -7386
rect 393294 -7654 393914 -7622
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 402294 705798 402914 711590
rect 402294 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 402914 705798
rect 402294 705478 402914 705562
rect 402294 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 402914 705478
rect 402294 691954 402914 705242
rect 402294 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 402914 691954
rect 402294 691634 402914 691718
rect 402294 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 402914 691634
rect 402294 655954 402914 691398
rect 402294 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 402914 655954
rect 402294 655634 402914 655718
rect 402294 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 402914 655634
rect 402294 619954 402914 655398
rect 402294 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 402914 619954
rect 402294 619634 402914 619718
rect 402294 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 402914 619634
rect 402294 583954 402914 619398
rect 402294 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 402914 583954
rect 402294 583634 402914 583718
rect 402294 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 402914 583634
rect 402294 547954 402914 583398
rect 402294 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 402914 547954
rect 402294 547634 402914 547718
rect 402294 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 402914 547634
rect 402294 511954 402914 547398
rect 402294 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 402914 511954
rect 402294 511634 402914 511718
rect 402294 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 402914 511634
rect 402294 475954 402914 511398
rect 402294 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 402914 475954
rect 402294 475634 402914 475718
rect 402294 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 402914 475634
rect 402294 439954 402914 475398
rect 402294 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 402914 439954
rect 402294 439634 402914 439718
rect 402294 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 402914 439634
rect 402294 403954 402914 439398
rect 402294 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 402914 403954
rect 402294 403634 402914 403718
rect 402294 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 402914 403634
rect 402294 367954 402914 403398
rect 402294 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 402914 367954
rect 402294 367634 402914 367718
rect 402294 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 402914 367634
rect 402294 331954 402914 367398
rect 402294 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 402914 331954
rect 402294 331634 402914 331718
rect 402294 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 402914 331634
rect 402294 295954 402914 331398
rect 402294 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 402914 295954
rect 402294 295634 402914 295718
rect 402294 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 402914 295634
rect 402294 259954 402914 295398
rect 402294 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 402914 259954
rect 402294 259634 402914 259718
rect 402294 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 402914 259634
rect 402294 223954 402914 259398
rect 402294 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 402914 223954
rect 402294 223634 402914 223718
rect 402294 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 402914 223634
rect 402294 187954 402914 223398
rect 402294 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 402914 187954
rect 402294 187634 402914 187718
rect 402294 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 402914 187634
rect 402294 151954 402914 187398
rect 402294 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 402914 151954
rect 402294 151634 402914 151718
rect 402294 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 402914 151634
rect 402294 115954 402914 151398
rect 402294 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 402914 115954
rect 402294 115634 402914 115718
rect 402294 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 402914 115634
rect 402294 79954 402914 115398
rect 402294 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 402914 79954
rect 402294 79634 402914 79718
rect 402294 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 402914 79634
rect 402294 43954 402914 79398
rect 402294 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 402914 43954
rect 402294 43634 402914 43718
rect 402294 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 402914 43634
rect 402294 7954 402914 43398
rect 402294 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 402914 7954
rect 402294 7634 402914 7718
rect 402294 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 402914 7634
rect 402294 -1306 402914 7398
rect 402294 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 402914 -1306
rect 402294 -1626 402914 -1542
rect 402294 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 402914 -1626
rect 402294 -7654 402914 -1862
rect 406794 706758 407414 711590
rect 406794 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 407414 706758
rect 406794 706438 407414 706522
rect 406794 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 407414 706438
rect 406794 696454 407414 706202
rect 406794 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 407414 696454
rect 406794 696134 407414 696218
rect 406794 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 407414 696134
rect 406794 660454 407414 695898
rect 406794 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 407414 660454
rect 406794 660134 407414 660218
rect 406794 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 407414 660134
rect 406794 624454 407414 659898
rect 406794 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 407414 624454
rect 406794 624134 407414 624218
rect 406794 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 407414 624134
rect 406794 588454 407414 623898
rect 406794 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 407414 588454
rect 406794 588134 407414 588218
rect 406794 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 407414 588134
rect 406794 552454 407414 587898
rect 406794 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 407414 552454
rect 406794 552134 407414 552218
rect 406794 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 407414 552134
rect 406794 516454 407414 551898
rect 406794 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 407414 516454
rect 406794 516134 407414 516218
rect 406794 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 407414 516134
rect 406794 480454 407414 515898
rect 406794 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 407414 480454
rect 406794 480134 407414 480218
rect 406794 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 407414 480134
rect 406794 444454 407414 479898
rect 406794 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 407414 444454
rect 406794 444134 407414 444218
rect 406794 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 407414 444134
rect 406794 408454 407414 443898
rect 406794 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 407414 408454
rect 406794 408134 407414 408218
rect 406794 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 407414 408134
rect 406794 372454 407414 407898
rect 406794 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 407414 372454
rect 406794 372134 407414 372218
rect 406794 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 407414 372134
rect 406794 336454 407414 371898
rect 406794 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 407414 336454
rect 406794 336134 407414 336218
rect 406794 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 407414 336134
rect 406794 300454 407414 335898
rect 406794 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 407414 300454
rect 406794 300134 407414 300218
rect 406794 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 407414 300134
rect 406794 264454 407414 299898
rect 406794 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 407414 264454
rect 406794 264134 407414 264218
rect 406794 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 407414 264134
rect 406794 228454 407414 263898
rect 406794 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 407414 228454
rect 406794 228134 407414 228218
rect 406794 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 407414 228134
rect 406794 192454 407414 227898
rect 406794 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 407414 192454
rect 406794 192134 407414 192218
rect 406794 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 407414 192134
rect 406794 156454 407414 191898
rect 406794 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 407414 156454
rect 406794 156134 407414 156218
rect 406794 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 407414 156134
rect 406794 120454 407414 155898
rect 406794 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 407414 120454
rect 406794 120134 407414 120218
rect 406794 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 407414 120134
rect 406794 84454 407414 119898
rect 406794 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 407414 84454
rect 406794 84134 407414 84218
rect 406794 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 407414 84134
rect 406794 48454 407414 83898
rect 406794 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 407414 48454
rect 406794 48134 407414 48218
rect 406794 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 407414 48134
rect 406794 12454 407414 47898
rect 406794 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 407414 12454
rect 406794 12134 407414 12218
rect 406794 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 407414 12134
rect 406794 -2266 407414 11898
rect 406794 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 407414 -2266
rect 406794 -2586 407414 -2502
rect 406794 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 407414 -2586
rect 406794 -7654 407414 -2822
rect 411294 707718 411914 711590
rect 411294 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 411914 707718
rect 411294 707398 411914 707482
rect 411294 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 411914 707398
rect 411294 700954 411914 707162
rect 411294 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 411914 700954
rect 411294 700634 411914 700718
rect 411294 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 411914 700634
rect 411294 664954 411914 700398
rect 411294 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 411914 664954
rect 411294 664634 411914 664718
rect 411294 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 411914 664634
rect 411294 628954 411914 664398
rect 411294 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 411914 628954
rect 411294 628634 411914 628718
rect 411294 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 411914 628634
rect 411294 592954 411914 628398
rect 411294 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 411914 592954
rect 411294 592634 411914 592718
rect 411294 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 411914 592634
rect 411294 556954 411914 592398
rect 411294 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 411914 556954
rect 411294 556634 411914 556718
rect 411294 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 411914 556634
rect 411294 520954 411914 556398
rect 411294 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 411914 520954
rect 411294 520634 411914 520718
rect 411294 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 411914 520634
rect 411294 484954 411914 520398
rect 411294 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 411914 484954
rect 411294 484634 411914 484718
rect 411294 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 411914 484634
rect 411294 448954 411914 484398
rect 411294 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 411914 448954
rect 411294 448634 411914 448718
rect 411294 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 411914 448634
rect 411294 412954 411914 448398
rect 411294 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 411914 412954
rect 411294 412634 411914 412718
rect 411294 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 411914 412634
rect 411294 376954 411914 412398
rect 411294 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 411914 376954
rect 411294 376634 411914 376718
rect 411294 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 411914 376634
rect 411294 340954 411914 376398
rect 411294 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 411914 340954
rect 411294 340634 411914 340718
rect 411294 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 411914 340634
rect 411294 304954 411914 340398
rect 411294 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 411914 304954
rect 411294 304634 411914 304718
rect 411294 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 411914 304634
rect 411294 268954 411914 304398
rect 411294 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 411914 268954
rect 411294 268634 411914 268718
rect 411294 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 411914 268634
rect 411294 232954 411914 268398
rect 411294 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 411914 232954
rect 411294 232634 411914 232718
rect 411294 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 411914 232634
rect 411294 196954 411914 232398
rect 411294 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 411914 196954
rect 411294 196634 411914 196718
rect 411294 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 411914 196634
rect 411294 160954 411914 196398
rect 411294 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 411914 160954
rect 411294 160634 411914 160718
rect 411294 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 411914 160634
rect 411294 124954 411914 160398
rect 411294 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 411914 124954
rect 411294 124634 411914 124718
rect 411294 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 411914 124634
rect 411294 88954 411914 124398
rect 411294 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 411914 88954
rect 411294 88634 411914 88718
rect 411294 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 411914 88634
rect 411294 52954 411914 88398
rect 411294 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 411914 52954
rect 411294 52634 411914 52718
rect 411294 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 411914 52634
rect 411294 16954 411914 52398
rect 411294 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 411914 16954
rect 411294 16634 411914 16718
rect 411294 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 411914 16634
rect 411294 -3226 411914 16398
rect 411294 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 411914 -3226
rect 411294 -3546 411914 -3462
rect 411294 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 411914 -3546
rect 411294 -7654 411914 -3782
rect 415794 708678 416414 711590
rect 415794 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 416414 708678
rect 415794 708358 416414 708442
rect 415794 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 416414 708358
rect 415794 669454 416414 708122
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -4186 416414 20898
rect 415794 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 416414 -4186
rect 415794 -4506 416414 -4422
rect 415794 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 416414 -4506
rect 415794 -7654 416414 -4742
rect 420294 709638 420914 711590
rect 420294 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 420914 709638
rect 420294 709318 420914 709402
rect 420294 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 420914 709318
rect 420294 673954 420914 709082
rect 420294 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 420914 673954
rect 420294 673634 420914 673718
rect 420294 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 420914 673634
rect 420294 637954 420914 673398
rect 420294 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 420914 637954
rect 420294 637634 420914 637718
rect 420294 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 420914 637634
rect 420294 601954 420914 637398
rect 420294 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 420914 601954
rect 420294 601634 420914 601718
rect 420294 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 420914 601634
rect 420294 565954 420914 601398
rect 420294 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 420914 565954
rect 420294 565634 420914 565718
rect 420294 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 420914 565634
rect 420294 529954 420914 565398
rect 420294 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 420914 529954
rect 420294 529634 420914 529718
rect 420294 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 420914 529634
rect 420294 493954 420914 529398
rect 420294 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 420914 493954
rect 420294 493634 420914 493718
rect 420294 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 420914 493634
rect 420294 457954 420914 493398
rect 420294 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 420914 457954
rect 420294 457634 420914 457718
rect 420294 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 420914 457634
rect 420294 421954 420914 457398
rect 420294 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 420914 421954
rect 420294 421634 420914 421718
rect 420294 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 420914 421634
rect 420294 385954 420914 421398
rect 420294 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 420914 385954
rect 420294 385634 420914 385718
rect 420294 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 420914 385634
rect 420294 349954 420914 385398
rect 420294 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 420914 349954
rect 420294 349634 420914 349718
rect 420294 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 420914 349634
rect 420294 313954 420914 349398
rect 420294 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 420914 313954
rect 420294 313634 420914 313718
rect 420294 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 420914 313634
rect 420294 277954 420914 313398
rect 420294 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 420914 277954
rect 420294 277634 420914 277718
rect 420294 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 420914 277634
rect 420294 241954 420914 277398
rect 420294 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 420914 241954
rect 420294 241634 420914 241718
rect 420294 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 420914 241634
rect 420294 205954 420914 241398
rect 420294 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 420914 205954
rect 420294 205634 420914 205718
rect 420294 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 420914 205634
rect 420294 169954 420914 205398
rect 420294 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 420914 169954
rect 420294 169634 420914 169718
rect 420294 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 420914 169634
rect 420294 133954 420914 169398
rect 420294 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 420914 133954
rect 420294 133634 420914 133718
rect 420294 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 420914 133634
rect 420294 97954 420914 133398
rect 420294 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 420914 97954
rect 420294 97634 420914 97718
rect 420294 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 420914 97634
rect 420294 61954 420914 97398
rect 420294 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 420914 61954
rect 420294 61634 420914 61718
rect 420294 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 420914 61634
rect 420294 25954 420914 61398
rect 420294 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 420914 25954
rect 420294 25634 420914 25718
rect 420294 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 420914 25634
rect 420294 -5146 420914 25398
rect 420294 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 420914 -5146
rect 420294 -5466 420914 -5382
rect 420294 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 420914 -5466
rect 420294 -7654 420914 -5702
rect 424794 710598 425414 711590
rect 424794 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 425414 710598
rect 424794 710278 425414 710362
rect 424794 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 425414 710278
rect 424794 678454 425414 710042
rect 424794 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 425414 678454
rect 424794 678134 425414 678218
rect 424794 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 425414 678134
rect 424794 642454 425414 677898
rect 424794 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 425414 642454
rect 424794 642134 425414 642218
rect 424794 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 425414 642134
rect 424794 606454 425414 641898
rect 424794 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 425414 606454
rect 424794 606134 425414 606218
rect 424794 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 425414 606134
rect 424794 570454 425414 605898
rect 424794 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 425414 570454
rect 424794 570134 425414 570218
rect 424794 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 425414 570134
rect 424794 534454 425414 569898
rect 424794 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 425414 534454
rect 424794 534134 425414 534218
rect 424794 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 425414 534134
rect 424794 498454 425414 533898
rect 424794 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 425414 498454
rect 424794 498134 425414 498218
rect 424794 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 425414 498134
rect 424794 462454 425414 497898
rect 424794 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 425414 462454
rect 424794 462134 425414 462218
rect 424794 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 425414 462134
rect 424794 426454 425414 461898
rect 424794 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 425414 426454
rect 424794 426134 425414 426218
rect 424794 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 425414 426134
rect 424794 390454 425414 425898
rect 424794 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 425414 390454
rect 424794 390134 425414 390218
rect 424794 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 425414 390134
rect 424794 354454 425414 389898
rect 424794 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 425414 354454
rect 424794 354134 425414 354218
rect 424794 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 425414 354134
rect 424794 318454 425414 353898
rect 424794 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 425414 318454
rect 424794 318134 425414 318218
rect 424794 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 425414 318134
rect 424794 282454 425414 317898
rect 424794 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 425414 282454
rect 424794 282134 425414 282218
rect 424794 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 425414 282134
rect 424794 246454 425414 281898
rect 424794 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 425414 246454
rect 424794 246134 425414 246218
rect 424794 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 425414 246134
rect 424794 210454 425414 245898
rect 424794 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 425414 210454
rect 424794 210134 425414 210218
rect 424794 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 425414 210134
rect 424794 174454 425414 209898
rect 424794 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 425414 174454
rect 424794 174134 425414 174218
rect 424794 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 425414 174134
rect 424794 138454 425414 173898
rect 424794 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 425414 138454
rect 424794 138134 425414 138218
rect 424794 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 425414 138134
rect 424794 102454 425414 137898
rect 424794 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 425414 102454
rect 424794 102134 425414 102218
rect 424794 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 425414 102134
rect 424794 66454 425414 101898
rect 424794 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 425414 66454
rect 424794 66134 425414 66218
rect 424794 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 425414 66134
rect 424794 30454 425414 65898
rect 424794 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 425414 30454
rect 424794 30134 425414 30218
rect 424794 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 425414 30134
rect 424794 -6106 425414 29898
rect 424794 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 425414 -6106
rect 424794 -6426 425414 -6342
rect 424794 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 425414 -6426
rect 424794 -7654 425414 -6662
rect 429294 711558 429914 711590
rect 429294 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 429914 711558
rect 429294 711238 429914 711322
rect 429294 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 429914 711238
rect 429294 682954 429914 711002
rect 429294 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 429914 682954
rect 429294 682634 429914 682718
rect 429294 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 429914 682634
rect 429294 646954 429914 682398
rect 429294 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 429914 646954
rect 429294 646634 429914 646718
rect 429294 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 429914 646634
rect 429294 610954 429914 646398
rect 429294 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 429914 610954
rect 429294 610634 429914 610718
rect 429294 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 429914 610634
rect 429294 574954 429914 610398
rect 429294 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 429914 574954
rect 429294 574634 429914 574718
rect 429294 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 429914 574634
rect 429294 538954 429914 574398
rect 429294 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 429914 538954
rect 429294 538634 429914 538718
rect 429294 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 429914 538634
rect 429294 502954 429914 538398
rect 429294 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 429914 502954
rect 429294 502634 429914 502718
rect 429294 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 429914 502634
rect 429294 466954 429914 502398
rect 429294 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 429914 466954
rect 429294 466634 429914 466718
rect 429294 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 429914 466634
rect 429294 430954 429914 466398
rect 429294 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 429914 430954
rect 429294 430634 429914 430718
rect 429294 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 429914 430634
rect 429294 394954 429914 430398
rect 429294 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 429914 394954
rect 429294 394634 429914 394718
rect 429294 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 429914 394634
rect 429294 358954 429914 394398
rect 429294 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 429914 358954
rect 429294 358634 429914 358718
rect 429294 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 429914 358634
rect 429294 322954 429914 358398
rect 429294 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 429914 322954
rect 429294 322634 429914 322718
rect 429294 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 429914 322634
rect 429294 286954 429914 322398
rect 429294 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 429914 286954
rect 429294 286634 429914 286718
rect 429294 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 429914 286634
rect 429294 250954 429914 286398
rect 429294 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 429914 250954
rect 429294 250634 429914 250718
rect 429294 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 429914 250634
rect 429294 214954 429914 250398
rect 429294 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 429914 214954
rect 429294 214634 429914 214718
rect 429294 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 429914 214634
rect 429294 178954 429914 214398
rect 429294 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 429914 178954
rect 429294 178634 429914 178718
rect 429294 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 429914 178634
rect 429294 142954 429914 178398
rect 429294 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 429914 142954
rect 429294 142634 429914 142718
rect 429294 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 429914 142634
rect 429294 106954 429914 142398
rect 429294 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 429914 106954
rect 429294 106634 429914 106718
rect 429294 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 429914 106634
rect 429294 70954 429914 106398
rect 429294 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 429914 70954
rect 429294 70634 429914 70718
rect 429294 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 429914 70634
rect 429294 34954 429914 70398
rect 429294 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 429914 34954
rect 429294 34634 429914 34718
rect 429294 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 429914 34634
rect 429294 -7066 429914 34398
rect 429294 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 429914 -7066
rect 429294 -7386 429914 -7302
rect 429294 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 429914 -7386
rect 429294 -7654 429914 -7622
rect 433794 704838 434414 711590
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 438294 705798 438914 711590
rect 438294 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 438914 705798
rect 438294 705478 438914 705562
rect 438294 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 438914 705478
rect 438294 691954 438914 705242
rect 438294 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 438914 691954
rect 438294 691634 438914 691718
rect 438294 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 438914 691634
rect 438294 655954 438914 691398
rect 438294 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 438914 655954
rect 438294 655634 438914 655718
rect 438294 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 438914 655634
rect 438294 619954 438914 655398
rect 438294 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 438914 619954
rect 438294 619634 438914 619718
rect 438294 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 438914 619634
rect 438294 583954 438914 619398
rect 438294 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 438914 583954
rect 438294 583634 438914 583718
rect 438294 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 438914 583634
rect 438294 547954 438914 583398
rect 438294 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 438914 547954
rect 438294 547634 438914 547718
rect 438294 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 438914 547634
rect 438294 511954 438914 547398
rect 438294 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 438914 511954
rect 438294 511634 438914 511718
rect 438294 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 438914 511634
rect 438294 475954 438914 511398
rect 438294 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 438914 475954
rect 438294 475634 438914 475718
rect 438294 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 438914 475634
rect 438294 439954 438914 475398
rect 438294 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 438914 439954
rect 438294 439634 438914 439718
rect 438294 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 438914 439634
rect 438294 403954 438914 439398
rect 438294 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 438914 403954
rect 438294 403634 438914 403718
rect 438294 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 438914 403634
rect 438294 367954 438914 403398
rect 438294 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 438914 367954
rect 438294 367634 438914 367718
rect 438294 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 438914 367634
rect 438294 331954 438914 367398
rect 438294 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 438914 331954
rect 438294 331634 438914 331718
rect 438294 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 438914 331634
rect 438294 295954 438914 331398
rect 438294 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 438914 295954
rect 438294 295634 438914 295718
rect 438294 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 438914 295634
rect 438294 259954 438914 295398
rect 438294 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 438914 259954
rect 438294 259634 438914 259718
rect 438294 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 438914 259634
rect 438294 223954 438914 259398
rect 438294 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 438914 223954
rect 438294 223634 438914 223718
rect 438294 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 438914 223634
rect 438294 187954 438914 223398
rect 438294 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 438914 187954
rect 438294 187634 438914 187718
rect 438294 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 438914 187634
rect 438294 151954 438914 187398
rect 438294 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 438914 151954
rect 438294 151634 438914 151718
rect 438294 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 438914 151634
rect 438294 115954 438914 151398
rect 438294 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 438914 115954
rect 438294 115634 438914 115718
rect 438294 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 438914 115634
rect 438294 79954 438914 115398
rect 438294 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 438914 79954
rect 438294 79634 438914 79718
rect 438294 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 438914 79634
rect 438294 43954 438914 79398
rect 438294 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 438914 43954
rect 438294 43634 438914 43718
rect 438294 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 438914 43634
rect 438294 7954 438914 43398
rect 438294 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 438914 7954
rect 438294 7634 438914 7718
rect 438294 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 438914 7634
rect 438294 -1306 438914 7398
rect 438294 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 438914 -1306
rect 438294 -1626 438914 -1542
rect 438294 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 438914 -1626
rect 438294 -7654 438914 -1862
rect 442794 706758 443414 711590
rect 442794 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 443414 706758
rect 442794 706438 443414 706522
rect 442794 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 443414 706438
rect 442794 696454 443414 706202
rect 442794 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 443414 696454
rect 442794 696134 443414 696218
rect 442794 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 443414 696134
rect 442794 660454 443414 695898
rect 442794 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 443414 660454
rect 442794 660134 443414 660218
rect 442794 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 443414 660134
rect 442794 624454 443414 659898
rect 442794 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 443414 624454
rect 442794 624134 443414 624218
rect 442794 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 443414 624134
rect 442794 588454 443414 623898
rect 442794 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 443414 588454
rect 442794 588134 443414 588218
rect 442794 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 443414 588134
rect 442794 552454 443414 587898
rect 442794 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 443414 552454
rect 442794 552134 443414 552218
rect 442794 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 443414 552134
rect 442794 516454 443414 551898
rect 442794 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 443414 516454
rect 442794 516134 443414 516218
rect 442794 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 443414 516134
rect 442794 480454 443414 515898
rect 442794 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 443414 480454
rect 442794 480134 443414 480218
rect 442794 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 443414 480134
rect 442794 444454 443414 479898
rect 442794 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 443414 444454
rect 442794 444134 443414 444218
rect 442794 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 443414 444134
rect 442794 408454 443414 443898
rect 442794 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 443414 408454
rect 442794 408134 443414 408218
rect 442794 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 443414 408134
rect 442794 372454 443414 407898
rect 442794 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 443414 372454
rect 442794 372134 443414 372218
rect 442794 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 443414 372134
rect 442794 336454 443414 371898
rect 442794 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 443414 336454
rect 442794 336134 443414 336218
rect 442794 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 443414 336134
rect 442794 300454 443414 335898
rect 442794 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 443414 300454
rect 442794 300134 443414 300218
rect 442794 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 443414 300134
rect 442794 264454 443414 299898
rect 442794 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 443414 264454
rect 442794 264134 443414 264218
rect 442794 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 443414 264134
rect 442794 228454 443414 263898
rect 442794 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 443414 228454
rect 442794 228134 443414 228218
rect 442794 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 443414 228134
rect 442794 192454 443414 227898
rect 442794 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 443414 192454
rect 442794 192134 443414 192218
rect 442794 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 443414 192134
rect 442794 156454 443414 191898
rect 442794 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 443414 156454
rect 442794 156134 443414 156218
rect 442794 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 443414 156134
rect 442794 120454 443414 155898
rect 442794 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 443414 120454
rect 442794 120134 443414 120218
rect 442794 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 443414 120134
rect 442794 84454 443414 119898
rect 442794 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 443414 84454
rect 442794 84134 443414 84218
rect 442794 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 443414 84134
rect 442794 48454 443414 83898
rect 442794 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 443414 48454
rect 442794 48134 443414 48218
rect 442794 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 443414 48134
rect 442794 12454 443414 47898
rect 442794 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 443414 12454
rect 442794 12134 443414 12218
rect 442794 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 443414 12134
rect 442794 -2266 443414 11898
rect 442794 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 443414 -2266
rect 442794 -2586 443414 -2502
rect 442794 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 443414 -2586
rect 442794 -7654 443414 -2822
rect 447294 707718 447914 711590
rect 447294 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 447914 707718
rect 447294 707398 447914 707482
rect 447294 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 447914 707398
rect 447294 700954 447914 707162
rect 447294 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 447914 700954
rect 447294 700634 447914 700718
rect 447294 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 447914 700634
rect 447294 664954 447914 700398
rect 447294 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 447914 664954
rect 447294 664634 447914 664718
rect 447294 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 447914 664634
rect 447294 628954 447914 664398
rect 447294 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 447914 628954
rect 447294 628634 447914 628718
rect 447294 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 447914 628634
rect 447294 592954 447914 628398
rect 447294 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 447914 592954
rect 447294 592634 447914 592718
rect 447294 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 447914 592634
rect 447294 556954 447914 592398
rect 447294 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 447914 556954
rect 447294 556634 447914 556718
rect 447294 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 447914 556634
rect 447294 520954 447914 556398
rect 447294 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 447914 520954
rect 447294 520634 447914 520718
rect 447294 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 447914 520634
rect 447294 484954 447914 520398
rect 447294 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 447914 484954
rect 447294 484634 447914 484718
rect 447294 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 447914 484634
rect 447294 448954 447914 484398
rect 447294 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 447914 448954
rect 447294 448634 447914 448718
rect 447294 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 447914 448634
rect 447294 412954 447914 448398
rect 447294 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 447914 412954
rect 447294 412634 447914 412718
rect 447294 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 447914 412634
rect 447294 376954 447914 412398
rect 447294 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 447914 376954
rect 447294 376634 447914 376718
rect 447294 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 447914 376634
rect 447294 340954 447914 376398
rect 447294 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 447914 340954
rect 447294 340634 447914 340718
rect 447294 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 447914 340634
rect 447294 304954 447914 340398
rect 447294 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 447914 304954
rect 447294 304634 447914 304718
rect 447294 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 447914 304634
rect 447294 268954 447914 304398
rect 447294 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 447914 268954
rect 447294 268634 447914 268718
rect 447294 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 447914 268634
rect 447294 232954 447914 268398
rect 447294 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 447914 232954
rect 447294 232634 447914 232718
rect 447294 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 447914 232634
rect 447294 196954 447914 232398
rect 447294 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 447914 196954
rect 447294 196634 447914 196718
rect 447294 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 447914 196634
rect 447294 160954 447914 196398
rect 447294 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 447914 160954
rect 447294 160634 447914 160718
rect 447294 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 447914 160634
rect 447294 124954 447914 160398
rect 447294 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 447914 124954
rect 447294 124634 447914 124718
rect 447294 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 447914 124634
rect 447294 88954 447914 124398
rect 447294 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 447914 88954
rect 447294 88634 447914 88718
rect 447294 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 447914 88634
rect 447294 52954 447914 88398
rect 447294 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 447914 52954
rect 447294 52634 447914 52718
rect 447294 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 447914 52634
rect 447294 16954 447914 52398
rect 447294 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 447914 16954
rect 447294 16634 447914 16718
rect 447294 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 447914 16634
rect 447294 -3226 447914 16398
rect 447294 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 447914 -3226
rect 447294 -3546 447914 -3462
rect 447294 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 447914 -3546
rect 447294 -7654 447914 -3782
rect 451794 708678 452414 711590
rect 451794 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 452414 708678
rect 451794 708358 452414 708442
rect 451794 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 452414 708358
rect 451794 669454 452414 708122
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -4186 452414 20898
rect 451794 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 452414 -4186
rect 451794 -4506 452414 -4422
rect 451794 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 452414 -4506
rect 451794 -7654 452414 -4742
rect 456294 709638 456914 711590
rect 456294 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 456914 709638
rect 456294 709318 456914 709402
rect 456294 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 456914 709318
rect 456294 673954 456914 709082
rect 456294 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 456914 673954
rect 456294 673634 456914 673718
rect 456294 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 456914 673634
rect 456294 637954 456914 673398
rect 456294 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 456914 637954
rect 456294 637634 456914 637718
rect 456294 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 456914 637634
rect 456294 601954 456914 637398
rect 456294 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 456914 601954
rect 456294 601634 456914 601718
rect 456294 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 456914 601634
rect 456294 565954 456914 601398
rect 456294 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 456914 565954
rect 456294 565634 456914 565718
rect 456294 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 456914 565634
rect 456294 529954 456914 565398
rect 456294 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 456914 529954
rect 456294 529634 456914 529718
rect 456294 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 456914 529634
rect 456294 493954 456914 529398
rect 456294 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 456914 493954
rect 456294 493634 456914 493718
rect 456294 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 456914 493634
rect 456294 457954 456914 493398
rect 456294 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 456914 457954
rect 456294 457634 456914 457718
rect 456294 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 456914 457634
rect 456294 421954 456914 457398
rect 456294 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 456914 421954
rect 456294 421634 456914 421718
rect 456294 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 456914 421634
rect 456294 385954 456914 421398
rect 456294 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 456914 385954
rect 456294 385634 456914 385718
rect 456294 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 456914 385634
rect 456294 349954 456914 385398
rect 456294 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 456914 349954
rect 456294 349634 456914 349718
rect 456294 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 456914 349634
rect 456294 313954 456914 349398
rect 456294 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 456914 313954
rect 456294 313634 456914 313718
rect 456294 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 456914 313634
rect 456294 277954 456914 313398
rect 456294 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 456914 277954
rect 456294 277634 456914 277718
rect 456294 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 456914 277634
rect 456294 241954 456914 277398
rect 456294 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 456914 241954
rect 456294 241634 456914 241718
rect 456294 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 456914 241634
rect 456294 205954 456914 241398
rect 456294 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 456914 205954
rect 456294 205634 456914 205718
rect 456294 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 456914 205634
rect 456294 169954 456914 205398
rect 456294 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 456914 169954
rect 456294 169634 456914 169718
rect 456294 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 456914 169634
rect 456294 133954 456914 169398
rect 456294 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 456914 133954
rect 456294 133634 456914 133718
rect 456294 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 456914 133634
rect 456294 97954 456914 133398
rect 456294 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 456914 97954
rect 456294 97634 456914 97718
rect 456294 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 456914 97634
rect 456294 61954 456914 97398
rect 456294 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 456914 61954
rect 456294 61634 456914 61718
rect 456294 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 456914 61634
rect 456294 25954 456914 61398
rect 456294 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 456914 25954
rect 456294 25634 456914 25718
rect 456294 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 456914 25634
rect 456294 -5146 456914 25398
rect 456294 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 456914 -5146
rect 456294 -5466 456914 -5382
rect 456294 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 456914 -5466
rect 456294 -7654 456914 -5702
rect 460794 710598 461414 711590
rect 460794 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 461414 710598
rect 460794 710278 461414 710362
rect 460794 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 461414 710278
rect 460794 678454 461414 710042
rect 460794 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 461414 678454
rect 460794 678134 461414 678218
rect 460794 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 461414 678134
rect 460794 642454 461414 677898
rect 460794 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 461414 642454
rect 460794 642134 461414 642218
rect 460794 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 461414 642134
rect 460794 606454 461414 641898
rect 460794 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 461414 606454
rect 460794 606134 461414 606218
rect 460794 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 461414 606134
rect 460794 570454 461414 605898
rect 460794 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 461414 570454
rect 460794 570134 461414 570218
rect 460794 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 461414 570134
rect 460794 534454 461414 569898
rect 460794 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 461414 534454
rect 460794 534134 461414 534218
rect 460794 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 461414 534134
rect 460794 498454 461414 533898
rect 460794 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 461414 498454
rect 460794 498134 461414 498218
rect 460794 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 461414 498134
rect 460794 462454 461414 497898
rect 460794 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 461414 462454
rect 460794 462134 461414 462218
rect 460794 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 461414 462134
rect 460794 426454 461414 461898
rect 460794 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 461414 426454
rect 460794 426134 461414 426218
rect 460794 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 461414 426134
rect 460794 390454 461414 425898
rect 460794 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 461414 390454
rect 460794 390134 461414 390218
rect 460794 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 461414 390134
rect 460794 354454 461414 389898
rect 460794 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 461414 354454
rect 460794 354134 461414 354218
rect 460794 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 461414 354134
rect 460794 318454 461414 353898
rect 460794 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 461414 318454
rect 460794 318134 461414 318218
rect 460794 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 461414 318134
rect 460794 282454 461414 317898
rect 460794 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 461414 282454
rect 460794 282134 461414 282218
rect 460794 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 461414 282134
rect 460794 246454 461414 281898
rect 460794 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 461414 246454
rect 460794 246134 461414 246218
rect 460794 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 461414 246134
rect 460794 210454 461414 245898
rect 460794 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 461414 210454
rect 460794 210134 461414 210218
rect 460794 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 461414 210134
rect 460794 174454 461414 209898
rect 460794 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 461414 174454
rect 460794 174134 461414 174218
rect 460794 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 461414 174134
rect 460794 138454 461414 173898
rect 460794 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 461414 138454
rect 460794 138134 461414 138218
rect 460794 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 461414 138134
rect 460794 102454 461414 137898
rect 460794 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 461414 102454
rect 460794 102134 461414 102218
rect 460794 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 461414 102134
rect 460794 66454 461414 101898
rect 460794 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 461414 66454
rect 460794 66134 461414 66218
rect 460794 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 461414 66134
rect 460794 30454 461414 65898
rect 460794 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 461414 30454
rect 460794 30134 461414 30218
rect 460794 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 461414 30134
rect 460794 -6106 461414 29898
rect 460794 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 461414 -6106
rect 460794 -6426 461414 -6342
rect 460794 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 461414 -6426
rect 460794 -7654 461414 -6662
rect 465294 711558 465914 711590
rect 465294 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 465914 711558
rect 465294 711238 465914 711322
rect 465294 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 465914 711238
rect 465294 682954 465914 711002
rect 465294 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 465914 682954
rect 465294 682634 465914 682718
rect 465294 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 465914 682634
rect 465294 646954 465914 682398
rect 465294 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 465914 646954
rect 465294 646634 465914 646718
rect 465294 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 465914 646634
rect 465294 610954 465914 646398
rect 465294 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 465914 610954
rect 465294 610634 465914 610718
rect 465294 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 465914 610634
rect 465294 574954 465914 610398
rect 465294 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 465914 574954
rect 465294 574634 465914 574718
rect 465294 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 465914 574634
rect 465294 538954 465914 574398
rect 465294 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 465914 538954
rect 465294 538634 465914 538718
rect 465294 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 465914 538634
rect 465294 502954 465914 538398
rect 465294 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 465914 502954
rect 465294 502634 465914 502718
rect 465294 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 465914 502634
rect 465294 466954 465914 502398
rect 465294 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 465914 466954
rect 465294 466634 465914 466718
rect 465294 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 465914 466634
rect 465294 430954 465914 466398
rect 465294 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 465914 430954
rect 465294 430634 465914 430718
rect 465294 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 465914 430634
rect 465294 394954 465914 430398
rect 465294 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 465914 394954
rect 465294 394634 465914 394718
rect 465294 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 465914 394634
rect 465294 358954 465914 394398
rect 465294 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 465914 358954
rect 465294 358634 465914 358718
rect 465294 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 465914 358634
rect 465294 322954 465914 358398
rect 465294 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 465914 322954
rect 465294 322634 465914 322718
rect 465294 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 465914 322634
rect 465294 286954 465914 322398
rect 465294 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 465914 286954
rect 465294 286634 465914 286718
rect 465294 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 465914 286634
rect 465294 250954 465914 286398
rect 465294 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 465914 250954
rect 465294 250634 465914 250718
rect 465294 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 465914 250634
rect 465294 214954 465914 250398
rect 465294 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 465914 214954
rect 465294 214634 465914 214718
rect 465294 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 465914 214634
rect 465294 178954 465914 214398
rect 465294 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 465914 178954
rect 465294 178634 465914 178718
rect 465294 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 465914 178634
rect 465294 142954 465914 178398
rect 465294 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 465914 142954
rect 465294 142634 465914 142718
rect 465294 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 465914 142634
rect 465294 106954 465914 142398
rect 465294 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 465914 106954
rect 465294 106634 465914 106718
rect 465294 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 465914 106634
rect 465294 70954 465914 106398
rect 465294 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 465914 70954
rect 465294 70634 465914 70718
rect 465294 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 465914 70634
rect 465294 34954 465914 70398
rect 465294 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 465914 34954
rect 465294 34634 465914 34718
rect 465294 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 465914 34634
rect 465294 -7066 465914 34398
rect 465294 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 465914 -7066
rect 465294 -7386 465914 -7302
rect 465294 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 465914 -7386
rect 465294 -7654 465914 -7622
rect 469794 704838 470414 711590
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 474294 705798 474914 711590
rect 474294 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 474914 705798
rect 474294 705478 474914 705562
rect 474294 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 474914 705478
rect 474294 691954 474914 705242
rect 474294 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 474914 691954
rect 474294 691634 474914 691718
rect 474294 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 474914 691634
rect 474294 655954 474914 691398
rect 474294 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 474914 655954
rect 474294 655634 474914 655718
rect 474294 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 474914 655634
rect 474294 619954 474914 655398
rect 474294 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 474914 619954
rect 474294 619634 474914 619718
rect 474294 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 474914 619634
rect 474294 583954 474914 619398
rect 474294 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 474914 583954
rect 474294 583634 474914 583718
rect 474294 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 474914 583634
rect 474294 547954 474914 583398
rect 474294 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 474914 547954
rect 474294 547634 474914 547718
rect 474294 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 474914 547634
rect 474294 511954 474914 547398
rect 474294 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 474914 511954
rect 474294 511634 474914 511718
rect 474294 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 474914 511634
rect 474294 475954 474914 511398
rect 474294 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 474914 475954
rect 474294 475634 474914 475718
rect 474294 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 474914 475634
rect 474294 439954 474914 475398
rect 474294 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 474914 439954
rect 474294 439634 474914 439718
rect 474294 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 474914 439634
rect 474294 403954 474914 439398
rect 474294 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 474914 403954
rect 474294 403634 474914 403718
rect 474294 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 474914 403634
rect 474294 367954 474914 403398
rect 474294 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 474914 367954
rect 474294 367634 474914 367718
rect 474294 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 474914 367634
rect 474294 331954 474914 367398
rect 474294 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 474914 331954
rect 474294 331634 474914 331718
rect 474294 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 474914 331634
rect 474294 295954 474914 331398
rect 474294 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 474914 295954
rect 474294 295634 474914 295718
rect 474294 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 474914 295634
rect 474294 259954 474914 295398
rect 474294 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 474914 259954
rect 474294 259634 474914 259718
rect 474294 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 474914 259634
rect 474294 223954 474914 259398
rect 474294 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 474914 223954
rect 474294 223634 474914 223718
rect 474294 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 474914 223634
rect 474294 187954 474914 223398
rect 474294 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 474914 187954
rect 474294 187634 474914 187718
rect 474294 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 474914 187634
rect 474294 151954 474914 187398
rect 474294 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 474914 151954
rect 474294 151634 474914 151718
rect 474294 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 474914 151634
rect 474294 115954 474914 151398
rect 474294 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 474914 115954
rect 474294 115634 474914 115718
rect 474294 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 474914 115634
rect 474294 79954 474914 115398
rect 474294 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 474914 79954
rect 474294 79634 474914 79718
rect 474294 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 474914 79634
rect 474294 43954 474914 79398
rect 474294 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 474914 43954
rect 474294 43634 474914 43718
rect 474294 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 474914 43634
rect 474294 7954 474914 43398
rect 474294 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 474914 7954
rect 474294 7634 474914 7718
rect 474294 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 474914 7634
rect 474294 -1306 474914 7398
rect 474294 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 474914 -1306
rect 474294 -1626 474914 -1542
rect 474294 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 474914 -1626
rect 474294 -7654 474914 -1862
rect 478794 706758 479414 711590
rect 478794 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 479414 706758
rect 478794 706438 479414 706522
rect 478794 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 479414 706438
rect 478794 696454 479414 706202
rect 478794 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 479414 696454
rect 478794 696134 479414 696218
rect 478794 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 479414 696134
rect 478794 660454 479414 695898
rect 478794 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 479414 660454
rect 478794 660134 479414 660218
rect 478794 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 479414 660134
rect 478794 624454 479414 659898
rect 478794 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 479414 624454
rect 478794 624134 479414 624218
rect 478794 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 479414 624134
rect 478794 588454 479414 623898
rect 478794 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 479414 588454
rect 478794 588134 479414 588218
rect 478794 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 479414 588134
rect 478794 552454 479414 587898
rect 478794 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 479414 552454
rect 478794 552134 479414 552218
rect 478794 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 479414 552134
rect 478794 516454 479414 551898
rect 478794 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 479414 516454
rect 478794 516134 479414 516218
rect 478794 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 479414 516134
rect 478794 480454 479414 515898
rect 478794 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 479414 480454
rect 478794 480134 479414 480218
rect 478794 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 479414 480134
rect 478794 444454 479414 479898
rect 478794 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 479414 444454
rect 478794 444134 479414 444218
rect 478794 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 479414 444134
rect 478794 408454 479414 443898
rect 478794 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 479414 408454
rect 478794 408134 479414 408218
rect 478794 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 479414 408134
rect 478794 372454 479414 407898
rect 478794 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 479414 372454
rect 478794 372134 479414 372218
rect 478794 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 479414 372134
rect 478794 336454 479414 371898
rect 478794 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 479414 336454
rect 478794 336134 479414 336218
rect 478794 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 479414 336134
rect 478794 300454 479414 335898
rect 478794 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 479414 300454
rect 478794 300134 479414 300218
rect 478794 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 479414 300134
rect 478794 264454 479414 299898
rect 478794 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 479414 264454
rect 478794 264134 479414 264218
rect 478794 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 479414 264134
rect 478794 228454 479414 263898
rect 478794 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 479414 228454
rect 478794 228134 479414 228218
rect 478794 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 479414 228134
rect 478794 192454 479414 227898
rect 478794 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 479414 192454
rect 478794 192134 479414 192218
rect 478794 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 479414 192134
rect 478794 156454 479414 191898
rect 478794 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 479414 156454
rect 478794 156134 479414 156218
rect 478794 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 479414 156134
rect 478794 120454 479414 155898
rect 478794 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 479414 120454
rect 478794 120134 479414 120218
rect 478794 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 479414 120134
rect 478794 84454 479414 119898
rect 478794 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 479414 84454
rect 478794 84134 479414 84218
rect 478794 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 479414 84134
rect 478794 48454 479414 83898
rect 478794 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 479414 48454
rect 478794 48134 479414 48218
rect 478794 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 479414 48134
rect 478794 12454 479414 47898
rect 478794 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 479414 12454
rect 478794 12134 479414 12218
rect 478794 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 479414 12134
rect 478794 -2266 479414 11898
rect 478794 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 479414 -2266
rect 478794 -2586 479414 -2502
rect 478794 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 479414 -2586
rect 478794 -7654 479414 -2822
rect 483294 707718 483914 711590
rect 483294 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 483914 707718
rect 483294 707398 483914 707482
rect 483294 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 483914 707398
rect 483294 700954 483914 707162
rect 483294 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 483914 700954
rect 483294 700634 483914 700718
rect 483294 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 483914 700634
rect 483294 664954 483914 700398
rect 483294 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 483914 664954
rect 483294 664634 483914 664718
rect 483294 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 483914 664634
rect 483294 628954 483914 664398
rect 483294 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 483914 628954
rect 483294 628634 483914 628718
rect 483294 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 483914 628634
rect 483294 592954 483914 628398
rect 483294 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 483914 592954
rect 483294 592634 483914 592718
rect 483294 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 483914 592634
rect 483294 556954 483914 592398
rect 483294 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 483914 556954
rect 483294 556634 483914 556718
rect 483294 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 483914 556634
rect 483294 520954 483914 556398
rect 483294 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 483914 520954
rect 483294 520634 483914 520718
rect 483294 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 483914 520634
rect 483294 484954 483914 520398
rect 483294 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 483914 484954
rect 483294 484634 483914 484718
rect 483294 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 483914 484634
rect 483294 448954 483914 484398
rect 483294 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 483914 448954
rect 483294 448634 483914 448718
rect 483294 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 483914 448634
rect 483294 412954 483914 448398
rect 483294 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 483914 412954
rect 483294 412634 483914 412718
rect 483294 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 483914 412634
rect 483294 376954 483914 412398
rect 483294 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 483914 376954
rect 483294 376634 483914 376718
rect 483294 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 483914 376634
rect 483294 340954 483914 376398
rect 483294 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 483914 340954
rect 483294 340634 483914 340718
rect 483294 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 483914 340634
rect 483294 304954 483914 340398
rect 483294 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 483914 304954
rect 483294 304634 483914 304718
rect 483294 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 483914 304634
rect 483294 268954 483914 304398
rect 483294 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 483914 268954
rect 483294 268634 483914 268718
rect 483294 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 483914 268634
rect 483294 232954 483914 268398
rect 483294 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 483914 232954
rect 483294 232634 483914 232718
rect 483294 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 483914 232634
rect 483294 196954 483914 232398
rect 483294 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 483914 196954
rect 483294 196634 483914 196718
rect 483294 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 483914 196634
rect 483294 160954 483914 196398
rect 483294 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 483914 160954
rect 483294 160634 483914 160718
rect 483294 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 483914 160634
rect 483294 124954 483914 160398
rect 483294 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 483914 124954
rect 483294 124634 483914 124718
rect 483294 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 483914 124634
rect 483294 88954 483914 124398
rect 483294 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 483914 88954
rect 483294 88634 483914 88718
rect 483294 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 483914 88634
rect 483294 52954 483914 88398
rect 483294 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 483914 52954
rect 483294 52634 483914 52718
rect 483294 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 483914 52634
rect 483294 16954 483914 52398
rect 483294 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 483914 16954
rect 483294 16634 483914 16718
rect 483294 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 483914 16634
rect 483294 -3226 483914 16398
rect 483294 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 483914 -3226
rect 483294 -3546 483914 -3462
rect 483294 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 483914 -3546
rect 483294 -7654 483914 -3782
rect 487794 708678 488414 711590
rect 487794 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 488414 708678
rect 487794 708358 488414 708442
rect 487794 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 488414 708358
rect 487794 669454 488414 708122
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -4186 488414 20898
rect 487794 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 488414 -4186
rect 487794 -4506 488414 -4422
rect 487794 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 488414 -4506
rect 487794 -7654 488414 -4742
rect 492294 709638 492914 711590
rect 492294 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 492914 709638
rect 492294 709318 492914 709402
rect 492294 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 492914 709318
rect 492294 673954 492914 709082
rect 492294 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 492914 673954
rect 492294 673634 492914 673718
rect 492294 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 492914 673634
rect 492294 637954 492914 673398
rect 492294 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 492914 637954
rect 492294 637634 492914 637718
rect 492294 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 492914 637634
rect 492294 601954 492914 637398
rect 492294 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 492914 601954
rect 492294 601634 492914 601718
rect 492294 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 492914 601634
rect 492294 565954 492914 601398
rect 492294 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 492914 565954
rect 492294 565634 492914 565718
rect 492294 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 492914 565634
rect 492294 529954 492914 565398
rect 492294 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 492914 529954
rect 492294 529634 492914 529718
rect 492294 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 492914 529634
rect 492294 493954 492914 529398
rect 492294 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 492914 493954
rect 492294 493634 492914 493718
rect 492294 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 492914 493634
rect 492294 457954 492914 493398
rect 492294 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 492914 457954
rect 492294 457634 492914 457718
rect 492294 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 492914 457634
rect 492294 421954 492914 457398
rect 492294 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 492914 421954
rect 492294 421634 492914 421718
rect 492294 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 492914 421634
rect 492294 385954 492914 421398
rect 492294 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 492914 385954
rect 492294 385634 492914 385718
rect 492294 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 492914 385634
rect 492294 349954 492914 385398
rect 492294 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 492914 349954
rect 492294 349634 492914 349718
rect 492294 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 492914 349634
rect 492294 313954 492914 349398
rect 492294 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 492914 313954
rect 492294 313634 492914 313718
rect 492294 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 492914 313634
rect 492294 277954 492914 313398
rect 492294 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 492914 277954
rect 492294 277634 492914 277718
rect 492294 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 492914 277634
rect 492294 241954 492914 277398
rect 492294 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 492914 241954
rect 492294 241634 492914 241718
rect 492294 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 492914 241634
rect 492294 205954 492914 241398
rect 492294 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 492914 205954
rect 492294 205634 492914 205718
rect 492294 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 492914 205634
rect 492294 169954 492914 205398
rect 492294 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 492914 169954
rect 492294 169634 492914 169718
rect 492294 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 492914 169634
rect 492294 133954 492914 169398
rect 492294 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 492914 133954
rect 492294 133634 492914 133718
rect 492294 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 492914 133634
rect 492294 97954 492914 133398
rect 492294 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 492914 97954
rect 492294 97634 492914 97718
rect 492294 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 492914 97634
rect 492294 61954 492914 97398
rect 492294 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 492914 61954
rect 492294 61634 492914 61718
rect 492294 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 492914 61634
rect 492294 25954 492914 61398
rect 492294 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 492914 25954
rect 492294 25634 492914 25718
rect 492294 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 492914 25634
rect 492294 -5146 492914 25398
rect 492294 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 492914 -5146
rect 492294 -5466 492914 -5382
rect 492294 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 492914 -5466
rect 492294 -7654 492914 -5702
rect 496794 710598 497414 711590
rect 496794 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 497414 710598
rect 496794 710278 497414 710362
rect 496794 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 497414 710278
rect 496794 678454 497414 710042
rect 496794 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 497414 678454
rect 496794 678134 497414 678218
rect 496794 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 497414 678134
rect 496794 642454 497414 677898
rect 496794 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 497414 642454
rect 496794 642134 497414 642218
rect 496794 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 497414 642134
rect 496794 606454 497414 641898
rect 496794 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 497414 606454
rect 496794 606134 497414 606218
rect 496794 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 497414 606134
rect 496794 570454 497414 605898
rect 496794 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 497414 570454
rect 496794 570134 497414 570218
rect 496794 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 497414 570134
rect 496794 534454 497414 569898
rect 496794 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 497414 534454
rect 496794 534134 497414 534218
rect 496794 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 497414 534134
rect 496794 498454 497414 533898
rect 496794 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 497414 498454
rect 496794 498134 497414 498218
rect 496794 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 497414 498134
rect 496794 462454 497414 497898
rect 496794 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 497414 462454
rect 496794 462134 497414 462218
rect 496794 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 497414 462134
rect 496794 426454 497414 461898
rect 496794 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 497414 426454
rect 496794 426134 497414 426218
rect 496794 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 497414 426134
rect 496794 390454 497414 425898
rect 496794 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 497414 390454
rect 496794 390134 497414 390218
rect 496794 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 497414 390134
rect 496794 354454 497414 389898
rect 496794 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 497414 354454
rect 496794 354134 497414 354218
rect 496794 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 497414 354134
rect 496794 318454 497414 353898
rect 496794 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 497414 318454
rect 496794 318134 497414 318218
rect 496794 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 497414 318134
rect 496794 282454 497414 317898
rect 496794 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 497414 282454
rect 496794 282134 497414 282218
rect 496794 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 497414 282134
rect 496794 246454 497414 281898
rect 496794 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 497414 246454
rect 496794 246134 497414 246218
rect 496794 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 497414 246134
rect 496794 210454 497414 245898
rect 496794 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 497414 210454
rect 496794 210134 497414 210218
rect 496794 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 497414 210134
rect 496794 174454 497414 209898
rect 496794 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 497414 174454
rect 496794 174134 497414 174218
rect 496794 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 497414 174134
rect 496794 138454 497414 173898
rect 496794 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 497414 138454
rect 496794 138134 497414 138218
rect 496794 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 497414 138134
rect 496794 102454 497414 137898
rect 496794 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 497414 102454
rect 496794 102134 497414 102218
rect 496794 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 497414 102134
rect 496794 66454 497414 101898
rect 496794 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 497414 66454
rect 496794 66134 497414 66218
rect 496794 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 497414 66134
rect 496794 30454 497414 65898
rect 496794 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 497414 30454
rect 496794 30134 497414 30218
rect 496794 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 497414 30134
rect 496794 -6106 497414 29898
rect 496794 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 497414 -6106
rect 496794 -6426 497414 -6342
rect 496794 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 497414 -6426
rect 496794 -7654 497414 -6662
rect 501294 711558 501914 711590
rect 501294 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 501914 711558
rect 501294 711238 501914 711322
rect 501294 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 501914 711238
rect 501294 682954 501914 711002
rect 501294 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 501914 682954
rect 501294 682634 501914 682718
rect 501294 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 501914 682634
rect 501294 646954 501914 682398
rect 501294 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 501914 646954
rect 501294 646634 501914 646718
rect 501294 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 501914 646634
rect 501294 610954 501914 646398
rect 501294 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 501914 610954
rect 501294 610634 501914 610718
rect 501294 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 501914 610634
rect 501294 574954 501914 610398
rect 501294 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 501914 574954
rect 501294 574634 501914 574718
rect 501294 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 501914 574634
rect 501294 538954 501914 574398
rect 501294 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 501914 538954
rect 501294 538634 501914 538718
rect 501294 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 501914 538634
rect 501294 502954 501914 538398
rect 501294 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 501914 502954
rect 501294 502634 501914 502718
rect 501294 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 501914 502634
rect 501294 466954 501914 502398
rect 501294 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 501914 466954
rect 501294 466634 501914 466718
rect 501294 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 501914 466634
rect 501294 430954 501914 466398
rect 501294 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 501914 430954
rect 501294 430634 501914 430718
rect 501294 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 501914 430634
rect 501294 394954 501914 430398
rect 501294 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 501914 394954
rect 501294 394634 501914 394718
rect 501294 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 501914 394634
rect 501294 358954 501914 394398
rect 501294 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 501914 358954
rect 501294 358634 501914 358718
rect 501294 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 501914 358634
rect 501294 322954 501914 358398
rect 501294 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 501914 322954
rect 501294 322634 501914 322718
rect 501294 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 501914 322634
rect 501294 286954 501914 322398
rect 501294 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 501914 286954
rect 501294 286634 501914 286718
rect 501294 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 501914 286634
rect 501294 250954 501914 286398
rect 501294 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 501914 250954
rect 501294 250634 501914 250718
rect 501294 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 501914 250634
rect 501294 214954 501914 250398
rect 501294 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 501914 214954
rect 501294 214634 501914 214718
rect 501294 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 501914 214634
rect 501294 178954 501914 214398
rect 501294 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 501914 178954
rect 501294 178634 501914 178718
rect 501294 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 501914 178634
rect 501294 142954 501914 178398
rect 501294 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 501914 142954
rect 501294 142634 501914 142718
rect 501294 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 501914 142634
rect 501294 106954 501914 142398
rect 501294 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 501914 106954
rect 501294 106634 501914 106718
rect 501294 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 501914 106634
rect 501294 70954 501914 106398
rect 501294 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 501914 70954
rect 501294 70634 501914 70718
rect 501294 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 501914 70634
rect 501294 34954 501914 70398
rect 501294 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 501914 34954
rect 501294 34634 501914 34718
rect 501294 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 501914 34634
rect 501294 -7066 501914 34398
rect 501294 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 501914 -7066
rect 501294 -7386 501914 -7302
rect 501294 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 501914 -7386
rect 501294 -7654 501914 -7622
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 510294 705798 510914 711590
rect 510294 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 510914 705798
rect 510294 705478 510914 705562
rect 510294 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 510914 705478
rect 510294 691954 510914 705242
rect 510294 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 510914 691954
rect 510294 691634 510914 691718
rect 510294 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 510914 691634
rect 510294 655954 510914 691398
rect 510294 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 510914 655954
rect 510294 655634 510914 655718
rect 510294 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 510914 655634
rect 510294 619954 510914 655398
rect 510294 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 510914 619954
rect 510294 619634 510914 619718
rect 510294 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 510914 619634
rect 510294 583954 510914 619398
rect 510294 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 510914 583954
rect 510294 583634 510914 583718
rect 510294 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 510914 583634
rect 510294 547954 510914 583398
rect 510294 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 510914 547954
rect 510294 547634 510914 547718
rect 510294 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 510914 547634
rect 510294 511954 510914 547398
rect 510294 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 510914 511954
rect 510294 511634 510914 511718
rect 510294 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 510914 511634
rect 510294 475954 510914 511398
rect 510294 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 510914 475954
rect 510294 475634 510914 475718
rect 510294 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 510914 475634
rect 510294 439954 510914 475398
rect 510294 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 510914 439954
rect 510294 439634 510914 439718
rect 510294 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 510914 439634
rect 510294 403954 510914 439398
rect 510294 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 510914 403954
rect 510294 403634 510914 403718
rect 510294 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 510914 403634
rect 510294 367954 510914 403398
rect 510294 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 510914 367954
rect 510294 367634 510914 367718
rect 510294 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 510914 367634
rect 510294 331954 510914 367398
rect 510294 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 510914 331954
rect 510294 331634 510914 331718
rect 510294 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 510914 331634
rect 510294 295954 510914 331398
rect 510294 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 510914 295954
rect 510294 295634 510914 295718
rect 510294 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 510914 295634
rect 510294 259954 510914 295398
rect 510294 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 510914 259954
rect 510294 259634 510914 259718
rect 510294 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 510914 259634
rect 510294 223954 510914 259398
rect 510294 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 510914 223954
rect 510294 223634 510914 223718
rect 510294 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 510914 223634
rect 510294 187954 510914 223398
rect 510294 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 510914 187954
rect 510294 187634 510914 187718
rect 510294 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 510914 187634
rect 510294 151954 510914 187398
rect 510294 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 510914 151954
rect 510294 151634 510914 151718
rect 510294 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 510914 151634
rect 510294 115954 510914 151398
rect 510294 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 510914 115954
rect 510294 115634 510914 115718
rect 510294 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 510914 115634
rect 510294 79954 510914 115398
rect 510294 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 510914 79954
rect 510294 79634 510914 79718
rect 510294 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 510914 79634
rect 510294 43954 510914 79398
rect 510294 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 510914 43954
rect 510294 43634 510914 43718
rect 510294 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 510914 43634
rect 510294 7954 510914 43398
rect 510294 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 510914 7954
rect 510294 7634 510914 7718
rect 510294 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 510914 7634
rect 510294 -1306 510914 7398
rect 510294 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 510914 -1306
rect 510294 -1626 510914 -1542
rect 510294 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 510914 -1626
rect 510294 -7654 510914 -1862
rect 514794 706758 515414 711590
rect 514794 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 515414 706758
rect 514794 706438 515414 706522
rect 514794 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 515414 706438
rect 514794 696454 515414 706202
rect 514794 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 515414 696454
rect 514794 696134 515414 696218
rect 514794 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 515414 696134
rect 514794 660454 515414 695898
rect 514794 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 515414 660454
rect 514794 660134 515414 660218
rect 514794 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 515414 660134
rect 514794 624454 515414 659898
rect 514794 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 515414 624454
rect 514794 624134 515414 624218
rect 514794 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 515414 624134
rect 514794 588454 515414 623898
rect 514794 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 515414 588454
rect 514794 588134 515414 588218
rect 514794 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 515414 588134
rect 514794 552454 515414 587898
rect 514794 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 515414 552454
rect 514794 552134 515414 552218
rect 514794 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 515414 552134
rect 514794 516454 515414 551898
rect 514794 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 515414 516454
rect 514794 516134 515414 516218
rect 514794 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 515414 516134
rect 514794 480454 515414 515898
rect 514794 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 515414 480454
rect 514794 480134 515414 480218
rect 514794 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 515414 480134
rect 514794 444454 515414 479898
rect 514794 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 515414 444454
rect 514794 444134 515414 444218
rect 514794 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 515414 444134
rect 514794 408454 515414 443898
rect 514794 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 515414 408454
rect 514794 408134 515414 408218
rect 514794 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 515414 408134
rect 514794 372454 515414 407898
rect 514794 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 515414 372454
rect 514794 372134 515414 372218
rect 514794 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 515414 372134
rect 514794 336454 515414 371898
rect 514794 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 515414 336454
rect 514794 336134 515414 336218
rect 514794 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 515414 336134
rect 514794 300454 515414 335898
rect 514794 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 515414 300454
rect 514794 300134 515414 300218
rect 514794 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 515414 300134
rect 514794 264454 515414 299898
rect 514794 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 515414 264454
rect 514794 264134 515414 264218
rect 514794 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 515414 264134
rect 514794 228454 515414 263898
rect 514794 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 515414 228454
rect 514794 228134 515414 228218
rect 514794 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 515414 228134
rect 514794 192454 515414 227898
rect 514794 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 515414 192454
rect 514794 192134 515414 192218
rect 514794 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 515414 192134
rect 514794 156454 515414 191898
rect 514794 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 515414 156454
rect 514794 156134 515414 156218
rect 514794 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 515414 156134
rect 514794 120454 515414 155898
rect 514794 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 515414 120454
rect 514794 120134 515414 120218
rect 514794 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 515414 120134
rect 514794 84454 515414 119898
rect 514794 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 515414 84454
rect 514794 84134 515414 84218
rect 514794 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 515414 84134
rect 514794 48454 515414 83898
rect 514794 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 515414 48454
rect 514794 48134 515414 48218
rect 514794 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 515414 48134
rect 514794 12454 515414 47898
rect 514794 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 515414 12454
rect 514794 12134 515414 12218
rect 514794 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 515414 12134
rect 514794 -2266 515414 11898
rect 514794 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 515414 -2266
rect 514794 -2586 515414 -2502
rect 514794 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 515414 -2586
rect 514794 -7654 515414 -2822
rect 519294 707718 519914 711590
rect 519294 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 519914 707718
rect 519294 707398 519914 707482
rect 519294 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 519914 707398
rect 519294 700954 519914 707162
rect 519294 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 519914 700954
rect 519294 700634 519914 700718
rect 519294 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 519914 700634
rect 519294 664954 519914 700398
rect 519294 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 519914 664954
rect 519294 664634 519914 664718
rect 519294 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 519914 664634
rect 519294 628954 519914 664398
rect 519294 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 519914 628954
rect 519294 628634 519914 628718
rect 519294 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 519914 628634
rect 519294 592954 519914 628398
rect 519294 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 519914 592954
rect 519294 592634 519914 592718
rect 519294 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 519914 592634
rect 519294 556954 519914 592398
rect 519294 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 519914 556954
rect 519294 556634 519914 556718
rect 519294 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 519914 556634
rect 519294 520954 519914 556398
rect 519294 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 519914 520954
rect 519294 520634 519914 520718
rect 519294 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 519914 520634
rect 519294 484954 519914 520398
rect 519294 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 519914 484954
rect 519294 484634 519914 484718
rect 519294 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 519914 484634
rect 519294 448954 519914 484398
rect 519294 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 519914 448954
rect 519294 448634 519914 448718
rect 519294 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 519914 448634
rect 519294 412954 519914 448398
rect 519294 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 519914 412954
rect 519294 412634 519914 412718
rect 519294 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 519914 412634
rect 519294 376954 519914 412398
rect 519294 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 519914 376954
rect 519294 376634 519914 376718
rect 519294 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 519914 376634
rect 519294 340954 519914 376398
rect 519294 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 519914 340954
rect 519294 340634 519914 340718
rect 519294 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 519914 340634
rect 519294 304954 519914 340398
rect 519294 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 519914 304954
rect 519294 304634 519914 304718
rect 519294 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 519914 304634
rect 519294 268954 519914 304398
rect 519294 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 519914 268954
rect 519294 268634 519914 268718
rect 519294 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 519914 268634
rect 519294 232954 519914 268398
rect 519294 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 519914 232954
rect 519294 232634 519914 232718
rect 519294 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 519914 232634
rect 519294 196954 519914 232398
rect 519294 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 519914 196954
rect 519294 196634 519914 196718
rect 519294 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 519914 196634
rect 519294 160954 519914 196398
rect 519294 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 519914 160954
rect 519294 160634 519914 160718
rect 519294 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 519914 160634
rect 519294 124954 519914 160398
rect 519294 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 519914 124954
rect 519294 124634 519914 124718
rect 519294 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 519914 124634
rect 519294 88954 519914 124398
rect 519294 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 519914 88954
rect 519294 88634 519914 88718
rect 519294 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 519914 88634
rect 519294 52954 519914 88398
rect 519294 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 519914 52954
rect 519294 52634 519914 52718
rect 519294 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 519914 52634
rect 519294 16954 519914 52398
rect 519294 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 519914 16954
rect 519294 16634 519914 16718
rect 519294 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 519914 16634
rect 519294 -3226 519914 16398
rect 519294 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 519914 -3226
rect 519294 -3546 519914 -3462
rect 519294 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 519914 -3546
rect 519294 -7654 519914 -3782
rect 523794 708678 524414 711590
rect 523794 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 524414 708678
rect 523794 708358 524414 708442
rect 523794 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 524414 708358
rect 523794 669454 524414 708122
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -4186 524414 20898
rect 523794 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 524414 -4186
rect 523794 -4506 524414 -4422
rect 523794 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 524414 -4506
rect 523794 -7654 524414 -4742
rect 528294 709638 528914 711590
rect 528294 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 528914 709638
rect 528294 709318 528914 709402
rect 528294 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 528914 709318
rect 528294 673954 528914 709082
rect 528294 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 528914 673954
rect 528294 673634 528914 673718
rect 528294 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 528914 673634
rect 528294 637954 528914 673398
rect 528294 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 528914 637954
rect 528294 637634 528914 637718
rect 528294 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 528914 637634
rect 528294 601954 528914 637398
rect 528294 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 528914 601954
rect 528294 601634 528914 601718
rect 528294 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 528914 601634
rect 528294 565954 528914 601398
rect 528294 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 528914 565954
rect 528294 565634 528914 565718
rect 528294 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 528914 565634
rect 528294 529954 528914 565398
rect 528294 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 528914 529954
rect 528294 529634 528914 529718
rect 528294 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 528914 529634
rect 528294 493954 528914 529398
rect 528294 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 528914 493954
rect 528294 493634 528914 493718
rect 528294 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 528914 493634
rect 528294 457954 528914 493398
rect 528294 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 528914 457954
rect 528294 457634 528914 457718
rect 528294 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 528914 457634
rect 528294 421954 528914 457398
rect 528294 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 528914 421954
rect 528294 421634 528914 421718
rect 528294 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 528914 421634
rect 528294 385954 528914 421398
rect 528294 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 528914 385954
rect 528294 385634 528914 385718
rect 528294 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 528914 385634
rect 528294 349954 528914 385398
rect 528294 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 528914 349954
rect 528294 349634 528914 349718
rect 528294 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 528914 349634
rect 528294 313954 528914 349398
rect 528294 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 528914 313954
rect 528294 313634 528914 313718
rect 528294 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 528914 313634
rect 528294 277954 528914 313398
rect 528294 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 528914 277954
rect 528294 277634 528914 277718
rect 528294 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 528914 277634
rect 528294 241954 528914 277398
rect 528294 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 528914 241954
rect 528294 241634 528914 241718
rect 528294 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 528914 241634
rect 528294 205954 528914 241398
rect 528294 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 528914 205954
rect 528294 205634 528914 205718
rect 528294 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 528914 205634
rect 528294 169954 528914 205398
rect 528294 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 528914 169954
rect 528294 169634 528914 169718
rect 528294 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 528914 169634
rect 528294 133954 528914 169398
rect 528294 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 528914 133954
rect 528294 133634 528914 133718
rect 528294 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 528914 133634
rect 528294 97954 528914 133398
rect 528294 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 528914 97954
rect 528294 97634 528914 97718
rect 528294 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 528914 97634
rect 528294 61954 528914 97398
rect 528294 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 528914 61954
rect 528294 61634 528914 61718
rect 528294 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 528914 61634
rect 528294 25954 528914 61398
rect 528294 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 528914 25954
rect 528294 25634 528914 25718
rect 528294 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 528914 25634
rect 528294 -5146 528914 25398
rect 528294 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 528914 -5146
rect 528294 -5466 528914 -5382
rect 528294 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 528914 -5466
rect 528294 -7654 528914 -5702
rect 532794 710598 533414 711590
rect 532794 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 533414 710598
rect 532794 710278 533414 710362
rect 532794 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 533414 710278
rect 532794 678454 533414 710042
rect 532794 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 533414 678454
rect 532794 678134 533414 678218
rect 532794 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 533414 678134
rect 532794 642454 533414 677898
rect 532794 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 533414 642454
rect 532794 642134 533414 642218
rect 532794 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 533414 642134
rect 532794 606454 533414 641898
rect 532794 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 533414 606454
rect 532794 606134 533414 606218
rect 532794 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 533414 606134
rect 532794 570454 533414 605898
rect 532794 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 533414 570454
rect 532794 570134 533414 570218
rect 532794 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 533414 570134
rect 532794 534454 533414 569898
rect 532794 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 533414 534454
rect 532794 534134 533414 534218
rect 532794 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 533414 534134
rect 532794 498454 533414 533898
rect 532794 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 533414 498454
rect 532794 498134 533414 498218
rect 532794 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 533414 498134
rect 532794 462454 533414 497898
rect 532794 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 533414 462454
rect 532794 462134 533414 462218
rect 532794 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 533414 462134
rect 532794 426454 533414 461898
rect 532794 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 533414 426454
rect 532794 426134 533414 426218
rect 532794 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 533414 426134
rect 532794 390454 533414 425898
rect 532794 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 533414 390454
rect 532794 390134 533414 390218
rect 532794 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 533414 390134
rect 532794 354454 533414 389898
rect 532794 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 533414 354454
rect 532794 354134 533414 354218
rect 532794 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 533414 354134
rect 532794 318454 533414 353898
rect 532794 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 533414 318454
rect 532794 318134 533414 318218
rect 532794 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 533414 318134
rect 532794 282454 533414 317898
rect 532794 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 533414 282454
rect 532794 282134 533414 282218
rect 532794 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 533414 282134
rect 532794 246454 533414 281898
rect 532794 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 533414 246454
rect 532794 246134 533414 246218
rect 532794 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 533414 246134
rect 532794 210454 533414 245898
rect 532794 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 533414 210454
rect 532794 210134 533414 210218
rect 532794 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 533414 210134
rect 532794 174454 533414 209898
rect 532794 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 533414 174454
rect 532794 174134 533414 174218
rect 532794 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 533414 174134
rect 532794 138454 533414 173898
rect 532794 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 533414 138454
rect 532794 138134 533414 138218
rect 532794 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 533414 138134
rect 532794 102454 533414 137898
rect 532794 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 533414 102454
rect 532794 102134 533414 102218
rect 532794 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 533414 102134
rect 532794 66454 533414 101898
rect 532794 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 533414 66454
rect 532794 66134 533414 66218
rect 532794 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 533414 66134
rect 532794 30454 533414 65898
rect 532794 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 533414 30454
rect 532794 30134 533414 30218
rect 532794 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 533414 30134
rect 532794 -6106 533414 29898
rect 532794 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 533414 -6106
rect 532794 -6426 533414 -6342
rect 532794 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 533414 -6426
rect 532794 -7654 533414 -6662
rect 537294 711558 537914 711590
rect 537294 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 537914 711558
rect 537294 711238 537914 711322
rect 537294 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 537914 711238
rect 537294 682954 537914 711002
rect 537294 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 537914 682954
rect 537294 682634 537914 682718
rect 537294 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 537914 682634
rect 537294 646954 537914 682398
rect 537294 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 537914 646954
rect 537294 646634 537914 646718
rect 537294 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 537914 646634
rect 537294 610954 537914 646398
rect 537294 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 537914 610954
rect 537294 610634 537914 610718
rect 537294 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 537914 610634
rect 537294 574954 537914 610398
rect 537294 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 537914 574954
rect 537294 574634 537914 574718
rect 537294 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 537914 574634
rect 537294 538954 537914 574398
rect 537294 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 537914 538954
rect 537294 538634 537914 538718
rect 537294 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 537914 538634
rect 537294 502954 537914 538398
rect 537294 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 537914 502954
rect 537294 502634 537914 502718
rect 537294 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 537914 502634
rect 537294 466954 537914 502398
rect 537294 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 537914 466954
rect 537294 466634 537914 466718
rect 537294 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 537914 466634
rect 537294 430954 537914 466398
rect 537294 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 537914 430954
rect 537294 430634 537914 430718
rect 537294 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 537914 430634
rect 537294 394954 537914 430398
rect 537294 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 537914 394954
rect 537294 394634 537914 394718
rect 537294 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 537914 394634
rect 537294 358954 537914 394398
rect 537294 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 537914 358954
rect 537294 358634 537914 358718
rect 537294 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 537914 358634
rect 537294 322954 537914 358398
rect 537294 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 537914 322954
rect 537294 322634 537914 322718
rect 537294 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 537914 322634
rect 537294 286954 537914 322398
rect 537294 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 537914 286954
rect 537294 286634 537914 286718
rect 537294 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 537914 286634
rect 537294 250954 537914 286398
rect 537294 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 537914 250954
rect 537294 250634 537914 250718
rect 537294 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 537914 250634
rect 537294 214954 537914 250398
rect 537294 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 537914 214954
rect 537294 214634 537914 214718
rect 537294 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 537914 214634
rect 537294 178954 537914 214398
rect 537294 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 537914 178954
rect 537294 178634 537914 178718
rect 537294 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 537914 178634
rect 537294 142954 537914 178398
rect 537294 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 537914 142954
rect 537294 142634 537914 142718
rect 537294 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 537914 142634
rect 537294 106954 537914 142398
rect 537294 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 537914 106954
rect 537294 106634 537914 106718
rect 537294 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 537914 106634
rect 537294 70954 537914 106398
rect 537294 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 537914 70954
rect 537294 70634 537914 70718
rect 537294 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 537914 70634
rect 537294 34954 537914 70398
rect 537294 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 537914 34954
rect 537294 34634 537914 34718
rect 537294 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 537914 34634
rect 537294 -7066 537914 34398
rect 537294 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 537914 -7066
rect 537294 -7386 537914 -7302
rect 537294 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 537914 -7386
rect 537294 -7654 537914 -7622
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 546294 705798 546914 711590
rect 546294 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 546914 705798
rect 546294 705478 546914 705562
rect 546294 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 546914 705478
rect 546294 691954 546914 705242
rect 546294 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 546914 691954
rect 546294 691634 546914 691718
rect 546294 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 546914 691634
rect 546294 655954 546914 691398
rect 546294 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 546914 655954
rect 546294 655634 546914 655718
rect 546294 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 546914 655634
rect 546294 619954 546914 655398
rect 546294 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 546914 619954
rect 546294 619634 546914 619718
rect 546294 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 546914 619634
rect 546294 583954 546914 619398
rect 546294 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 546914 583954
rect 546294 583634 546914 583718
rect 546294 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 546914 583634
rect 546294 547954 546914 583398
rect 546294 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 546914 547954
rect 546294 547634 546914 547718
rect 546294 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 546914 547634
rect 546294 511954 546914 547398
rect 546294 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 546914 511954
rect 546294 511634 546914 511718
rect 546294 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 546914 511634
rect 546294 475954 546914 511398
rect 546294 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 546914 475954
rect 546294 475634 546914 475718
rect 546294 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 546914 475634
rect 546294 439954 546914 475398
rect 546294 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 546914 439954
rect 546294 439634 546914 439718
rect 546294 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 546914 439634
rect 546294 403954 546914 439398
rect 546294 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 546914 403954
rect 546294 403634 546914 403718
rect 546294 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 546914 403634
rect 546294 367954 546914 403398
rect 546294 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 546914 367954
rect 546294 367634 546914 367718
rect 546294 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 546914 367634
rect 546294 331954 546914 367398
rect 546294 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 546914 331954
rect 546294 331634 546914 331718
rect 546294 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 546914 331634
rect 546294 295954 546914 331398
rect 546294 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 546914 295954
rect 546294 295634 546914 295718
rect 546294 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 546914 295634
rect 546294 259954 546914 295398
rect 546294 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 546914 259954
rect 546294 259634 546914 259718
rect 546294 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 546914 259634
rect 546294 223954 546914 259398
rect 546294 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 546914 223954
rect 546294 223634 546914 223718
rect 546294 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 546914 223634
rect 546294 187954 546914 223398
rect 546294 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 546914 187954
rect 546294 187634 546914 187718
rect 546294 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 546914 187634
rect 546294 151954 546914 187398
rect 546294 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 546914 151954
rect 546294 151634 546914 151718
rect 546294 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 546914 151634
rect 546294 115954 546914 151398
rect 546294 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 546914 115954
rect 546294 115634 546914 115718
rect 546294 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 546914 115634
rect 546294 79954 546914 115398
rect 546294 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 546914 79954
rect 546294 79634 546914 79718
rect 546294 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 546914 79634
rect 546294 43954 546914 79398
rect 546294 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 546914 43954
rect 546294 43634 546914 43718
rect 546294 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 546914 43634
rect 546294 7954 546914 43398
rect 546294 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 546914 7954
rect 546294 7634 546914 7718
rect 546294 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 546914 7634
rect 546294 -1306 546914 7398
rect 546294 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 546914 -1306
rect 546294 -1626 546914 -1542
rect 546294 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 546914 -1626
rect 546294 -7654 546914 -1862
rect 550794 706758 551414 711590
rect 550794 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 551414 706758
rect 550794 706438 551414 706522
rect 550794 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 551414 706438
rect 550794 696454 551414 706202
rect 550794 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 551414 696454
rect 550794 696134 551414 696218
rect 550794 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 551414 696134
rect 550794 660454 551414 695898
rect 550794 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 551414 660454
rect 550794 660134 551414 660218
rect 550794 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 551414 660134
rect 550794 624454 551414 659898
rect 550794 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 551414 624454
rect 550794 624134 551414 624218
rect 550794 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 551414 624134
rect 550794 588454 551414 623898
rect 550794 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 551414 588454
rect 550794 588134 551414 588218
rect 550794 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 551414 588134
rect 550794 552454 551414 587898
rect 550794 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 551414 552454
rect 550794 552134 551414 552218
rect 550794 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 551414 552134
rect 550794 516454 551414 551898
rect 550794 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 551414 516454
rect 550794 516134 551414 516218
rect 550794 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 551414 516134
rect 550794 480454 551414 515898
rect 550794 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 551414 480454
rect 550794 480134 551414 480218
rect 550794 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 551414 480134
rect 550794 444454 551414 479898
rect 550794 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 551414 444454
rect 550794 444134 551414 444218
rect 550794 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 551414 444134
rect 550794 408454 551414 443898
rect 550794 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 551414 408454
rect 550794 408134 551414 408218
rect 550794 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 551414 408134
rect 550794 372454 551414 407898
rect 550794 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 551414 372454
rect 550794 372134 551414 372218
rect 550794 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 551414 372134
rect 550794 336454 551414 371898
rect 550794 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 551414 336454
rect 550794 336134 551414 336218
rect 550794 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 551414 336134
rect 550794 300454 551414 335898
rect 550794 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 551414 300454
rect 550794 300134 551414 300218
rect 550794 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 551414 300134
rect 550794 264454 551414 299898
rect 550794 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 551414 264454
rect 550794 264134 551414 264218
rect 550794 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 551414 264134
rect 550794 228454 551414 263898
rect 550794 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 551414 228454
rect 550794 228134 551414 228218
rect 550794 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 551414 228134
rect 550794 192454 551414 227898
rect 550794 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 551414 192454
rect 550794 192134 551414 192218
rect 550794 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 551414 192134
rect 550794 156454 551414 191898
rect 550794 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 551414 156454
rect 550794 156134 551414 156218
rect 550794 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 551414 156134
rect 550794 120454 551414 155898
rect 550794 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 551414 120454
rect 550794 120134 551414 120218
rect 550794 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 551414 120134
rect 550794 84454 551414 119898
rect 550794 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 551414 84454
rect 550794 84134 551414 84218
rect 550794 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 551414 84134
rect 550794 48454 551414 83898
rect 550794 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 551414 48454
rect 550794 48134 551414 48218
rect 550794 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 551414 48134
rect 550794 12454 551414 47898
rect 550794 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 551414 12454
rect 550794 12134 551414 12218
rect 550794 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 551414 12134
rect 550794 -2266 551414 11898
rect 550794 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 551414 -2266
rect 550794 -2586 551414 -2502
rect 550794 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 551414 -2586
rect 550794 -7654 551414 -2822
rect 555294 707718 555914 711590
rect 555294 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 555914 707718
rect 555294 707398 555914 707482
rect 555294 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 555914 707398
rect 555294 700954 555914 707162
rect 555294 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 555914 700954
rect 555294 700634 555914 700718
rect 555294 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 555914 700634
rect 555294 664954 555914 700398
rect 555294 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 555914 664954
rect 555294 664634 555914 664718
rect 555294 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 555914 664634
rect 555294 628954 555914 664398
rect 555294 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 555914 628954
rect 555294 628634 555914 628718
rect 555294 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 555914 628634
rect 555294 592954 555914 628398
rect 555294 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 555914 592954
rect 555294 592634 555914 592718
rect 555294 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 555914 592634
rect 555294 556954 555914 592398
rect 555294 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 555914 556954
rect 555294 556634 555914 556718
rect 555294 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 555914 556634
rect 555294 520954 555914 556398
rect 555294 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 555914 520954
rect 555294 520634 555914 520718
rect 555294 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 555914 520634
rect 555294 484954 555914 520398
rect 555294 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 555914 484954
rect 555294 484634 555914 484718
rect 555294 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 555914 484634
rect 555294 448954 555914 484398
rect 555294 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 555914 448954
rect 555294 448634 555914 448718
rect 555294 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 555914 448634
rect 555294 412954 555914 448398
rect 555294 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 555914 412954
rect 555294 412634 555914 412718
rect 555294 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 555914 412634
rect 555294 376954 555914 412398
rect 555294 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 555914 376954
rect 555294 376634 555914 376718
rect 555294 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 555914 376634
rect 555294 340954 555914 376398
rect 555294 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 555914 340954
rect 555294 340634 555914 340718
rect 555294 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 555914 340634
rect 555294 304954 555914 340398
rect 555294 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 555914 304954
rect 555294 304634 555914 304718
rect 555294 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 555914 304634
rect 555294 268954 555914 304398
rect 555294 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 555914 268954
rect 555294 268634 555914 268718
rect 555294 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 555914 268634
rect 555294 232954 555914 268398
rect 555294 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 555914 232954
rect 555294 232634 555914 232718
rect 555294 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 555914 232634
rect 555294 196954 555914 232398
rect 555294 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 555914 196954
rect 555294 196634 555914 196718
rect 555294 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 555914 196634
rect 555294 160954 555914 196398
rect 555294 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 555914 160954
rect 555294 160634 555914 160718
rect 555294 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 555914 160634
rect 555294 124954 555914 160398
rect 555294 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 555914 124954
rect 555294 124634 555914 124718
rect 555294 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 555914 124634
rect 555294 88954 555914 124398
rect 555294 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 555914 88954
rect 555294 88634 555914 88718
rect 555294 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 555914 88634
rect 555294 52954 555914 88398
rect 555294 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 555914 52954
rect 555294 52634 555914 52718
rect 555294 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 555914 52634
rect 555294 16954 555914 52398
rect 555294 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 555914 16954
rect 555294 16634 555914 16718
rect 555294 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 555914 16634
rect 555294 -3226 555914 16398
rect 555294 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 555914 -3226
rect 555294 -3546 555914 -3462
rect 555294 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 555914 -3546
rect 555294 -7654 555914 -3782
rect 559794 708678 560414 711590
rect 559794 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 560414 708678
rect 559794 708358 560414 708442
rect 559794 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 560414 708358
rect 559794 669454 560414 708122
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -4186 560414 20898
rect 559794 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 560414 -4186
rect 559794 -4506 560414 -4422
rect 559794 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 560414 -4506
rect 559794 -7654 560414 -4742
rect 564294 709638 564914 711590
rect 564294 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 564914 709638
rect 564294 709318 564914 709402
rect 564294 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 564914 709318
rect 564294 673954 564914 709082
rect 564294 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 564914 673954
rect 564294 673634 564914 673718
rect 564294 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 564914 673634
rect 564294 637954 564914 673398
rect 564294 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 564914 637954
rect 564294 637634 564914 637718
rect 564294 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 564914 637634
rect 564294 601954 564914 637398
rect 564294 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 564914 601954
rect 564294 601634 564914 601718
rect 564294 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 564914 601634
rect 564294 565954 564914 601398
rect 564294 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 564914 565954
rect 564294 565634 564914 565718
rect 564294 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 564914 565634
rect 564294 529954 564914 565398
rect 564294 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 564914 529954
rect 564294 529634 564914 529718
rect 564294 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 564914 529634
rect 564294 493954 564914 529398
rect 564294 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 564914 493954
rect 564294 493634 564914 493718
rect 564294 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 564914 493634
rect 564294 457954 564914 493398
rect 564294 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 564914 457954
rect 564294 457634 564914 457718
rect 564294 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 564914 457634
rect 564294 421954 564914 457398
rect 564294 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 564914 421954
rect 564294 421634 564914 421718
rect 564294 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 564914 421634
rect 564294 385954 564914 421398
rect 564294 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 564914 385954
rect 564294 385634 564914 385718
rect 564294 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 564914 385634
rect 564294 349954 564914 385398
rect 564294 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 564914 349954
rect 564294 349634 564914 349718
rect 564294 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 564914 349634
rect 564294 313954 564914 349398
rect 564294 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 564914 313954
rect 564294 313634 564914 313718
rect 564294 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 564914 313634
rect 564294 277954 564914 313398
rect 564294 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 564914 277954
rect 564294 277634 564914 277718
rect 564294 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 564914 277634
rect 564294 241954 564914 277398
rect 564294 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 564914 241954
rect 564294 241634 564914 241718
rect 564294 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 564914 241634
rect 564294 205954 564914 241398
rect 564294 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 564914 205954
rect 564294 205634 564914 205718
rect 564294 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 564914 205634
rect 564294 169954 564914 205398
rect 564294 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 564914 169954
rect 564294 169634 564914 169718
rect 564294 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 564914 169634
rect 564294 133954 564914 169398
rect 564294 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 564914 133954
rect 564294 133634 564914 133718
rect 564294 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 564914 133634
rect 564294 97954 564914 133398
rect 564294 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 564914 97954
rect 564294 97634 564914 97718
rect 564294 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 564914 97634
rect 564294 61954 564914 97398
rect 564294 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 564914 61954
rect 564294 61634 564914 61718
rect 564294 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 564914 61634
rect 564294 25954 564914 61398
rect 564294 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 564914 25954
rect 564294 25634 564914 25718
rect 564294 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 564914 25634
rect 564294 -5146 564914 25398
rect 564294 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 564914 -5146
rect 564294 -5466 564914 -5382
rect 564294 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 564914 -5466
rect 564294 -7654 564914 -5702
rect 568794 710598 569414 711590
rect 568794 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 569414 710598
rect 568794 710278 569414 710362
rect 568794 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 569414 710278
rect 568794 678454 569414 710042
rect 568794 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 569414 678454
rect 568794 678134 569414 678218
rect 568794 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 569414 678134
rect 568794 642454 569414 677898
rect 568794 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 569414 642454
rect 568794 642134 569414 642218
rect 568794 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 569414 642134
rect 568794 606454 569414 641898
rect 568794 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 569414 606454
rect 568794 606134 569414 606218
rect 568794 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 569414 606134
rect 568794 570454 569414 605898
rect 568794 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 569414 570454
rect 568794 570134 569414 570218
rect 568794 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 569414 570134
rect 568794 534454 569414 569898
rect 568794 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 569414 534454
rect 568794 534134 569414 534218
rect 568794 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 569414 534134
rect 568794 498454 569414 533898
rect 568794 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 569414 498454
rect 568794 498134 569414 498218
rect 568794 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 569414 498134
rect 568794 462454 569414 497898
rect 568794 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 569414 462454
rect 568794 462134 569414 462218
rect 568794 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 569414 462134
rect 568794 426454 569414 461898
rect 568794 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 569414 426454
rect 568794 426134 569414 426218
rect 568794 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 569414 426134
rect 568794 390454 569414 425898
rect 568794 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 569414 390454
rect 568794 390134 569414 390218
rect 568794 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 569414 390134
rect 568794 354454 569414 389898
rect 568794 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 569414 354454
rect 568794 354134 569414 354218
rect 568794 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 569414 354134
rect 568794 318454 569414 353898
rect 568794 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 569414 318454
rect 568794 318134 569414 318218
rect 568794 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 569414 318134
rect 568794 282454 569414 317898
rect 568794 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 569414 282454
rect 568794 282134 569414 282218
rect 568794 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 569414 282134
rect 568794 246454 569414 281898
rect 568794 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 569414 246454
rect 568794 246134 569414 246218
rect 568794 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 569414 246134
rect 568794 210454 569414 245898
rect 568794 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 569414 210454
rect 568794 210134 569414 210218
rect 568794 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 569414 210134
rect 568794 174454 569414 209898
rect 568794 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 569414 174454
rect 568794 174134 569414 174218
rect 568794 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 569414 174134
rect 568794 138454 569414 173898
rect 568794 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 569414 138454
rect 568794 138134 569414 138218
rect 568794 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 569414 138134
rect 568794 102454 569414 137898
rect 568794 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 569414 102454
rect 568794 102134 569414 102218
rect 568794 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 569414 102134
rect 568794 66454 569414 101898
rect 568794 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 569414 66454
rect 568794 66134 569414 66218
rect 568794 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 569414 66134
rect 568794 30454 569414 65898
rect 568794 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 569414 30454
rect 568794 30134 569414 30218
rect 568794 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 569414 30134
rect 568794 -6106 569414 29898
rect 568794 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 569414 -6106
rect 568794 -6426 569414 -6342
rect 568794 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 569414 -6426
rect 568794 -7654 569414 -6662
rect 573294 711558 573914 711590
rect 573294 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 573914 711558
rect 573294 711238 573914 711322
rect 573294 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 573914 711238
rect 573294 682954 573914 711002
rect 573294 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 573914 682954
rect 573294 682634 573914 682718
rect 573294 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 573914 682634
rect 573294 646954 573914 682398
rect 573294 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 573914 646954
rect 573294 646634 573914 646718
rect 573294 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 573914 646634
rect 573294 610954 573914 646398
rect 573294 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 573914 610954
rect 573294 610634 573914 610718
rect 573294 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 573914 610634
rect 573294 574954 573914 610398
rect 573294 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 573914 574954
rect 573294 574634 573914 574718
rect 573294 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 573914 574634
rect 573294 538954 573914 574398
rect 573294 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 573914 538954
rect 573294 538634 573914 538718
rect 573294 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 573914 538634
rect 573294 502954 573914 538398
rect 573294 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 573914 502954
rect 573294 502634 573914 502718
rect 573294 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 573914 502634
rect 573294 466954 573914 502398
rect 573294 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 573914 466954
rect 573294 466634 573914 466718
rect 573294 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 573914 466634
rect 573294 430954 573914 466398
rect 573294 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 573914 430954
rect 573294 430634 573914 430718
rect 573294 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 573914 430634
rect 573294 394954 573914 430398
rect 573294 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 573914 394954
rect 573294 394634 573914 394718
rect 573294 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 573914 394634
rect 573294 358954 573914 394398
rect 573294 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 573914 358954
rect 573294 358634 573914 358718
rect 573294 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 573914 358634
rect 573294 322954 573914 358398
rect 573294 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 573914 322954
rect 573294 322634 573914 322718
rect 573294 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 573914 322634
rect 573294 286954 573914 322398
rect 573294 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 573914 286954
rect 573294 286634 573914 286718
rect 573294 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 573914 286634
rect 573294 250954 573914 286398
rect 573294 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 573914 250954
rect 573294 250634 573914 250718
rect 573294 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 573914 250634
rect 573294 214954 573914 250398
rect 573294 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 573914 214954
rect 573294 214634 573914 214718
rect 573294 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 573914 214634
rect 573294 178954 573914 214398
rect 573294 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 573914 178954
rect 573294 178634 573914 178718
rect 573294 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 573914 178634
rect 573294 142954 573914 178398
rect 573294 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 573914 142954
rect 573294 142634 573914 142718
rect 573294 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 573914 142634
rect 573294 106954 573914 142398
rect 573294 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 573914 106954
rect 573294 106634 573914 106718
rect 573294 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 573914 106634
rect 573294 70954 573914 106398
rect 573294 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 573914 70954
rect 573294 70634 573914 70718
rect 573294 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 573914 70634
rect 573294 34954 573914 70398
rect 573294 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 573914 34954
rect 573294 34634 573914 34718
rect 573294 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 573914 34634
rect 573294 -7066 573914 34398
rect 573294 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 573914 -7066
rect 573294 -7386 573914 -7302
rect 573294 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 573914 -7386
rect 573294 -7654 573914 -7622
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 582294 705798 582914 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 582294 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 582914 705798
rect 582294 705478 582914 705562
rect 582294 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 582914 705478
rect 582294 691954 582914 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 582294 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 582914 691954
rect 582294 691634 582914 691718
rect 582294 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 582914 691634
rect 582294 655954 582914 691398
rect 582294 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 582914 655954
rect 582294 655634 582914 655718
rect 582294 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 582914 655634
rect 582294 619954 582914 655398
rect 582294 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 582914 619954
rect 582294 619634 582914 619718
rect 582294 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 582914 619634
rect 582294 583954 582914 619398
rect 582294 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 582914 583954
rect 582294 583634 582914 583718
rect 582294 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 582914 583634
rect 582294 547954 582914 583398
rect 582294 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 582914 547954
rect 582294 547634 582914 547718
rect 582294 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 582914 547634
rect 582294 511954 582914 547398
rect 582294 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 582914 511954
rect 582294 511634 582914 511718
rect 582294 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 582914 511634
rect 582294 475954 582914 511398
rect 582294 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 582914 475954
rect 582294 475634 582914 475718
rect 582294 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 582914 475634
rect 582294 439954 582914 475398
rect 582294 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 582914 439954
rect 582294 439634 582914 439718
rect 582294 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 582914 439634
rect 582294 403954 582914 439398
rect 582294 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 582914 403954
rect 582294 403634 582914 403718
rect 582294 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 582914 403634
rect 582294 367954 582914 403398
rect 582294 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 582914 367954
rect 582294 367634 582914 367718
rect 582294 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 582914 367634
rect 582294 331954 582914 367398
rect 582294 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 582914 331954
rect 582294 331634 582914 331718
rect 582294 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 582914 331634
rect 582294 295954 582914 331398
rect 582294 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 582914 295954
rect 582294 295634 582914 295718
rect 582294 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 582914 295634
rect 582294 259954 582914 295398
rect 582294 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 582914 259954
rect 582294 259634 582914 259718
rect 582294 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 582914 259634
rect 582294 223954 582914 259398
rect 582294 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 582914 223954
rect 582294 223634 582914 223718
rect 582294 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 582914 223634
rect 582294 187954 582914 223398
rect 582294 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 582914 187954
rect 582294 187634 582914 187718
rect 582294 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 582914 187634
rect 582294 151954 582914 187398
rect 582294 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 582914 151954
rect 582294 151634 582914 151718
rect 582294 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 582914 151634
rect 582294 115954 582914 151398
rect 582294 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 582914 115954
rect 582294 115634 582914 115718
rect 582294 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 582914 115634
rect 582294 79954 582914 115398
rect 582294 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 582914 79954
rect 582294 79634 582914 79718
rect 582294 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 582914 79634
rect 582294 43954 582914 79398
rect 582294 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 582914 43954
rect 582294 43634 582914 43718
rect 582294 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 582914 43634
rect 582294 7954 582914 43398
rect 582294 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 582914 7954
rect 582294 7634 582914 7718
rect 582294 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 582914 7634
rect 582294 -1306 582914 7398
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691954 586890 705242
rect 586270 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 586890 691954
rect 586270 691634 586890 691718
rect 586270 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 586890 691634
rect 586270 655954 586890 691398
rect 586270 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 586890 655954
rect 586270 655634 586890 655718
rect 586270 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 586890 655634
rect 586270 619954 586890 655398
rect 586270 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 586890 619954
rect 586270 619634 586890 619718
rect 586270 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 586890 619634
rect 586270 583954 586890 619398
rect 586270 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 586890 583954
rect 586270 583634 586890 583718
rect 586270 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 586890 583634
rect 586270 547954 586890 583398
rect 586270 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 586890 547954
rect 586270 547634 586890 547718
rect 586270 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 586890 547634
rect 586270 511954 586890 547398
rect 586270 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 586890 511954
rect 586270 511634 586890 511718
rect 586270 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 586890 511634
rect 586270 475954 586890 511398
rect 586270 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 586890 475954
rect 586270 475634 586890 475718
rect 586270 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 586890 475634
rect 586270 439954 586890 475398
rect 586270 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 586890 439954
rect 586270 439634 586890 439718
rect 586270 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 586890 439634
rect 586270 403954 586890 439398
rect 586270 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 586890 403954
rect 586270 403634 586890 403718
rect 586270 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 586890 403634
rect 586270 367954 586890 403398
rect 586270 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 586890 367954
rect 586270 367634 586890 367718
rect 586270 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 586890 367634
rect 586270 331954 586890 367398
rect 586270 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 586890 331954
rect 586270 331634 586890 331718
rect 586270 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 586890 331634
rect 586270 295954 586890 331398
rect 586270 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 586890 295954
rect 586270 295634 586890 295718
rect 586270 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 586890 295634
rect 586270 259954 586890 295398
rect 586270 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 586890 259954
rect 586270 259634 586890 259718
rect 586270 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 586890 259634
rect 586270 223954 586890 259398
rect 586270 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 586890 223954
rect 586270 223634 586890 223718
rect 586270 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 586890 223634
rect 586270 187954 586890 223398
rect 586270 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 586890 187954
rect 586270 187634 586890 187718
rect 586270 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 586890 187634
rect 586270 151954 586890 187398
rect 586270 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 586890 151954
rect 586270 151634 586890 151718
rect 586270 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 586890 151634
rect 586270 115954 586890 151398
rect 586270 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 586890 115954
rect 586270 115634 586890 115718
rect 586270 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 586890 115634
rect 586270 79954 586890 115398
rect 586270 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 586890 79954
rect 586270 79634 586890 79718
rect 586270 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 586890 79634
rect 586270 43954 586890 79398
rect 586270 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 586890 43954
rect 586270 43634 586890 43718
rect 586270 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 586890 43634
rect 586270 7954 586890 43398
rect 586270 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 586890 7954
rect 586270 7634 586890 7718
rect 586270 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 586890 7634
rect 582294 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 582914 -1306
rect 582294 -1626 582914 -1542
rect 582294 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 582914 -1626
rect 582294 -7654 582914 -1862
rect 586270 -1306 586890 7398
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 696454 587850 706202
rect 587230 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 587850 696454
rect 587230 696134 587850 696218
rect 587230 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 587850 696134
rect 587230 660454 587850 695898
rect 587230 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 587850 660454
rect 587230 660134 587850 660218
rect 587230 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 587850 660134
rect 587230 624454 587850 659898
rect 587230 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 587850 624454
rect 587230 624134 587850 624218
rect 587230 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 587850 624134
rect 587230 588454 587850 623898
rect 587230 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 587850 588454
rect 587230 588134 587850 588218
rect 587230 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 587850 588134
rect 587230 552454 587850 587898
rect 587230 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 587850 552454
rect 587230 552134 587850 552218
rect 587230 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 587850 552134
rect 587230 516454 587850 551898
rect 587230 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 587850 516454
rect 587230 516134 587850 516218
rect 587230 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 587850 516134
rect 587230 480454 587850 515898
rect 587230 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 587850 480454
rect 587230 480134 587850 480218
rect 587230 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 587850 480134
rect 587230 444454 587850 479898
rect 587230 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 587850 444454
rect 587230 444134 587850 444218
rect 587230 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 587850 444134
rect 587230 408454 587850 443898
rect 587230 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 587850 408454
rect 587230 408134 587850 408218
rect 587230 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 587850 408134
rect 587230 372454 587850 407898
rect 587230 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 587850 372454
rect 587230 372134 587850 372218
rect 587230 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 587850 372134
rect 587230 336454 587850 371898
rect 587230 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 587850 336454
rect 587230 336134 587850 336218
rect 587230 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 587850 336134
rect 587230 300454 587850 335898
rect 587230 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 587850 300454
rect 587230 300134 587850 300218
rect 587230 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 587850 300134
rect 587230 264454 587850 299898
rect 587230 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 587850 264454
rect 587230 264134 587850 264218
rect 587230 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 587850 264134
rect 587230 228454 587850 263898
rect 587230 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 587850 228454
rect 587230 228134 587850 228218
rect 587230 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 587850 228134
rect 587230 192454 587850 227898
rect 587230 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 587850 192454
rect 587230 192134 587850 192218
rect 587230 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 587850 192134
rect 587230 156454 587850 191898
rect 587230 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 587850 156454
rect 587230 156134 587850 156218
rect 587230 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 587850 156134
rect 587230 120454 587850 155898
rect 587230 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 587850 120454
rect 587230 120134 587850 120218
rect 587230 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 587850 120134
rect 587230 84454 587850 119898
rect 587230 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 587850 84454
rect 587230 84134 587850 84218
rect 587230 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 587850 84134
rect 587230 48454 587850 83898
rect 587230 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 587850 48454
rect 587230 48134 587850 48218
rect 587230 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 587850 48134
rect 587230 12454 587850 47898
rect 587230 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 587850 12454
rect 587230 12134 587850 12218
rect 587230 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 587850 12134
rect 587230 -2266 587850 11898
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 700954 588810 707162
rect 588190 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 588810 700954
rect 588190 700634 588810 700718
rect 588190 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 588810 700634
rect 588190 664954 588810 700398
rect 588190 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 588810 664954
rect 588190 664634 588810 664718
rect 588190 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 588810 664634
rect 588190 628954 588810 664398
rect 588190 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 588810 628954
rect 588190 628634 588810 628718
rect 588190 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 588810 628634
rect 588190 592954 588810 628398
rect 588190 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 588810 592954
rect 588190 592634 588810 592718
rect 588190 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 588810 592634
rect 588190 556954 588810 592398
rect 588190 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 588810 556954
rect 588190 556634 588810 556718
rect 588190 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 588810 556634
rect 588190 520954 588810 556398
rect 588190 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 588810 520954
rect 588190 520634 588810 520718
rect 588190 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 588810 520634
rect 588190 484954 588810 520398
rect 588190 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 588810 484954
rect 588190 484634 588810 484718
rect 588190 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 588810 484634
rect 588190 448954 588810 484398
rect 588190 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 588810 448954
rect 588190 448634 588810 448718
rect 588190 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 588810 448634
rect 588190 412954 588810 448398
rect 588190 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 588810 412954
rect 588190 412634 588810 412718
rect 588190 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 588810 412634
rect 588190 376954 588810 412398
rect 588190 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 588810 376954
rect 588190 376634 588810 376718
rect 588190 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 588810 376634
rect 588190 340954 588810 376398
rect 588190 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 588810 340954
rect 588190 340634 588810 340718
rect 588190 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 588810 340634
rect 588190 304954 588810 340398
rect 588190 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 588810 304954
rect 588190 304634 588810 304718
rect 588190 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 588810 304634
rect 588190 268954 588810 304398
rect 588190 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 588810 268954
rect 588190 268634 588810 268718
rect 588190 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 588810 268634
rect 588190 232954 588810 268398
rect 588190 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 588810 232954
rect 588190 232634 588810 232718
rect 588190 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 588810 232634
rect 588190 196954 588810 232398
rect 588190 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 588810 196954
rect 588190 196634 588810 196718
rect 588190 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 588810 196634
rect 588190 160954 588810 196398
rect 588190 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 588810 160954
rect 588190 160634 588810 160718
rect 588190 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 588810 160634
rect 588190 124954 588810 160398
rect 588190 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 588810 124954
rect 588190 124634 588810 124718
rect 588190 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 588810 124634
rect 588190 88954 588810 124398
rect 588190 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 588810 88954
rect 588190 88634 588810 88718
rect 588190 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 588810 88634
rect 588190 52954 588810 88398
rect 588190 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 588810 52954
rect 588190 52634 588810 52718
rect 588190 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 588810 52634
rect 588190 16954 588810 52398
rect 588190 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 588810 16954
rect 588190 16634 588810 16718
rect 588190 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 588810 16634
rect 588190 -3226 588810 16398
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 669454 589770 708122
rect 589150 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 589770 669454
rect 589150 669134 589770 669218
rect 589150 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 589770 669134
rect 589150 633454 589770 668898
rect 589150 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 589770 633454
rect 589150 633134 589770 633218
rect 589150 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 589770 633134
rect 589150 597454 589770 632898
rect 589150 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 589770 597454
rect 589150 597134 589770 597218
rect 589150 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 589770 597134
rect 589150 561454 589770 596898
rect 589150 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 589770 561454
rect 589150 561134 589770 561218
rect 589150 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 589770 561134
rect 589150 525454 589770 560898
rect 589150 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 589770 525454
rect 589150 525134 589770 525218
rect 589150 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 589770 525134
rect 589150 489454 589770 524898
rect 589150 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 589770 489454
rect 589150 489134 589770 489218
rect 589150 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 589770 489134
rect 589150 453454 589770 488898
rect 589150 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 589770 453454
rect 589150 453134 589770 453218
rect 589150 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 589770 453134
rect 589150 417454 589770 452898
rect 589150 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 589770 417454
rect 589150 417134 589770 417218
rect 589150 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 589770 417134
rect 589150 381454 589770 416898
rect 589150 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 589770 381454
rect 589150 381134 589770 381218
rect 589150 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 589770 381134
rect 589150 345454 589770 380898
rect 589150 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 589770 345454
rect 589150 345134 589770 345218
rect 589150 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 589770 345134
rect 589150 309454 589770 344898
rect 589150 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 589770 309454
rect 589150 309134 589770 309218
rect 589150 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 589770 309134
rect 589150 273454 589770 308898
rect 589150 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 589770 273454
rect 589150 273134 589770 273218
rect 589150 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 589770 273134
rect 589150 237454 589770 272898
rect 589150 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 589770 237454
rect 589150 237134 589770 237218
rect 589150 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 589770 237134
rect 589150 201454 589770 236898
rect 589150 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 589770 201454
rect 589150 201134 589770 201218
rect 589150 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 589770 201134
rect 589150 165454 589770 200898
rect 589150 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 589770 165454
rect 589150 165134 589770 165218
rect 589150 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 589770 165134
rect 589150 129454 589770 164898
rect 589150 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 589770 129454
rect 589150 129134 589770 129218
rect 589150 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 589770 129134
rect 589150 93454 589770 128898
rect 589150 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 589770 93454
rect 589150 93134 589770 93218
rect 589150 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 589770 93134
rect 589150 57454 589770 92898
rect 589150 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 589770 57454
rect 589150 57134 589770 57218
rect 589150 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 589770 57134
rect 589150 21454 589770 56898
rect 589150 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 589770 21454
rect 589150 21134 589770 21218
rect 589150 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 589770 21134
rect 589150 -4186 589770 20898
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 673954 590730 709082
rect 590110 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 590730 673954
rect 590110 673634 590730 673718
rect 590110 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 590730 673634
rect 590110 637954 590730 673398
rect 590110 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 590730 637954
rect 590110 637634 590730 637718
rect 590110 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 590730 637634
rect 590110 601954 590730 637398
rect 590110 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 590730 601954
rect 590110 601634 590730 601718
rect 590110 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 590730 601634
rect 590110 565954 590730 601398
rect 590110 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 590730 565954
rect 590110 565634 590730 565718
rect 590110 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 590730 565634
rect 590110 529954 590730 565398
rect 590110 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 590730 529954
rect 590110 529634 590730 529718
rect 590110 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 590730 529634
rect 590110 493954 590730 529398
rect 590110 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 590730 493954
rect 590110 493634 590730 493718
rect 590110 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 590730 493634
rect 590110 457954 590730 493398
rect 590110 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 590730 457954
rect 590110 457634 590730 457718
rect 590110 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 590730 457634
rect 590110 421954 590730 457398
rect 590110 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 590730 421954
rect 590110 421634 590730 421718
rect 590110 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 590730 421634
rect 590110 385954 590730 421398
rect 590110 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 590730 385954
rect 590110 385634 590730 385718
rect 590110 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 590730 385634
rect 590110 349954 590730 385398
rect 590110 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 590730 349954
rect 590110 349634 590730 349718
rect 590110 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 590730 349634
rect 590110 313954 590730 349398
rect 590110 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 590730 313954
rect 590110 313634 590730 313718
rect 590110 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 590730 313634
rect 590110 277954 590730 313398
rect 590110 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 590730 277954
rect 590110 277634 590730 277718
rect 590110 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 590730 277634
rect 590110 241954 590730 277398
rect 590110 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 590730 241954
rect 590110 241634 590730 241718
rect 590110 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 590730 241634
rect 590110 205954 590730 241398
rect 590110 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 590730 205954
rect 590110 205634 590730 205718
rect 590110 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 590730 205634
rect 590110 169954 590730 205398
rect 590110 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 590730 169954
rect 590110 169634 590730 169718
rect 590110 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 590730 169634
rect 590110 133954 590730 169398
rect 590110 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 590730 133954
rect 590110 133634 590730 133718
rect 590110 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 590730 133634
rect 590110 97954 590730 133398
rect 590110 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 590730 97954
rect 590110 97634 590730 97718
rect 590110 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 590730 97634
rect 590110 61954 590730 97398
rect 590110 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 590730 61954
rect 590110 61634 590730 61718
rect 590110 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 590730 61634
rect 590110 25954 590730 61398
rect 590110 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 590730 25954
rect 590110 25634 590730 25718
rect 590110 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 590730 25634
rect 590110 -5146 590730 25398
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 678454 591690 710042
rect 591070 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 591690 678454
rect 591070 678134 591690 678218
rect 591070 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 591690 678134
rect 591070 642454 591690 677898
rect 591070 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 591690 642454
rect 591070 642134 591690 642218
rect 591070 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 591690 642134
rect 591070 606454 591690 641898
rect 591070 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 591690 606454
rect 591070 606134 591690 606218
rect 591070 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 591690 606134
rect 591070 570454 591690 605898
rect 591070 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 591690 570454
rect 591070 570134 591690 570218
rect 591070 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 591690 570134
rect 591070 534454 591690 569898
rect 591070 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 591690 534454
rect 591070 534134 591690 534218
rect 591070 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 591690 534134
rect 591070 498454 591690 533898
rect 591070 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 591690 498454
rect 591070 498134 591690 498218
rect 591070 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 591690 498134
rect 591070 462454 591690 497898
rect 591070 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 591690 462454
rect 591070 462134 591690 462218
rect 591070 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 591690 462134
rect 591070 426454 591690 461898
rect 591070 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 591690 426454
rect 591070 426134 591690 426218
rect 591070 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 591690 426134
rect 591070 390454 591690 425898
rect 591070 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 591690 390454
rect 591070 390134 591690 390218
rect 591070 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 591690 390134
rect 591070 354454 591690 389898
rect 591070 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 591690 354454
rect 591070 354134 591690 354218
rect 591070 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 591690 354134
rect 591070 318454 591690 353898
rect 591070 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 591690 318454
rect 591070 318134 591690 318218
rect 591070 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 591690 318134
rect 591070 282454 591690 317898
rect 591070 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 591690 282454
rect 591070 282134 591690 282218
rect 591070 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 591690 282134
rect 591070 246454 591690 281898
rect 591070 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 591690 246454
rect 591070 246134 591690 246218
rect 591070 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 591690 246134
rect 591070 210454 591690 245898
rect 591070 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 591690 210454
rect 591070 210134 591690 210218
rect 591070 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 591690 210134
rect 591070 174454 591690 209898
rect 591070 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 591690 174454
rect 591070 174134 591690 174218
rect 591070 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 591690 174134
rect 591070 138454 591690 173898
rect 591070 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 591690 138454
rect 591070 138134 591690 138218
rect 591070 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 591690 138134
rect 591070 102454 591690 137898
rect 591070 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 591690 102454
rect 591070 102134 591690 102218
rect 591070 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 591690 102134
rect 591070 66454 591690 101898
rect 591070 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 591690 66454
rect 591070 66134 591690 66218
rect 591070 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 591690 66134
rect 591070 30454 591690 65898
rect 591070 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 591690 30454
rect 591070 30134 591690 30218
rect 591070 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 591690 30134
rect 591070 -6106 591690 29898
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 682954 592650 711002
rect 592030 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect 592030 682634 592650 682718
rect 592030 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect 592030 646954 592650 682398
rect 592030 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect 592030 646634 592650 646718
rect 592030 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect 592030 610954 592650 646398
rect 592030 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect 592030 610634 592650 610718
rect 592030 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect 592030 574954 592650 610398
rect 592030 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect 592030 574634 592650 574718
rect 592030 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect 592030 538954 592650 574398
rect 592030 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect 592030 538634 592650 538718
rect 592030 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect 592030 502954 592650 538398
rect 592030 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect 592030 502634 592650 502718
rect 592030 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect 592030 466954 592650 502398
rect 592030 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect 592030 466634 592650 466718
rect 592030 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect 592030 430954 592650 466398
rect 592030 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect 592030 430634 592650 430718
rect 592030 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect 592030 394954 592650 430398
rect 592030 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect 592030 394634 592650 394718
rect 592030 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect 592030 358954 592650 394398
rect 592030 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect 592030 358634 592650 358718
rect 592030 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect 592030 322954 592650 358398
rect 592030 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect 592030 322634 592650 322718
rect 592030 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect 592030 286954 592650 322398
rect 592030 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect 592030 286634 592650 286718
rect 592030 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect 592030 250954 592650 286398
rect 592030 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect 592030 250634 592650 250718
rect 592030 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect 592030 214954 592650 250398
rect 592030 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect 592030 214634 592650 214718
rect 592030 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect 592030 178954 592650 214398
rect 592030 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect 592030 178634 592650 178718
rect 592030 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect 592030 142954 592650 178398
rect 592030 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect 592030 142634 592650 142718
rect 592030 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect 592030 106954 592650 142398
rect 592030 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect 592030 106634 592650 106718
rect 592030 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect 592030 70954 592650 106398
rect 592030 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect 592030 70634 592650 70718
rect 592030 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect 592030 34954 592650 70398
rect 592030 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect 592030 34634 592650 34718
rect 592030 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect 592030 -7066 592650 34398
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 682718 -8458 682954
rect -8374 682718 -8138 682954
rect -8694 682398 -8458 682634
rect -8374 682398 -8138 682634
rect -8694 646718 -8458 646954
rect -8374 646718 -8138 646954
rect -8694 646398 -8458 646634
rect -8374 646398 -8138 646634
rect -8694 610718 -8458 610954
rect -8374 610718 -8138 610954
rect -8694 610398 -8458 610634
rect -8374 610398 -8138 610634
rect -8694 574718 -8458 574954
rect -8374 574718 -8138 574954
rect -8694 574398 -8458 574634
rect -8374 574398 -8138 574634
rect -8694 538718 -8458 538954
rect -8374 538718 -8138 538954
rect -8694 538398 -8458 538634
rect -8374 538398 -8138 538634
rect -8694 502718 -8458 502954
rect -8374 502718 -8138 502954
rect -8694 502398 -8458 502634
rect -8374 502398 -8138 502634
rect -8694 466718 -8458 466954
rect -8374 466718 -8138 466954
rect -8694 466398 -8458 466634
rect -8374 466398 -8138 466634
rect -8694 430718 -8458 430954
rect -8374 430718 -8138 430954
rect -8694 430398 -8458 430634
rect -8374 430398 -8138 430634
rect -8694 394718 -8458 394954
rect -8374 394718 -8138 394954
rect -8694 394398 -8458 394634
rect -8374 394398 -8138 394634
rect -8694 358718 -8458 358954
rect -8374 358718 -8138 358954
rect -8694 358398 -8458 358634
rect -8374 358398 -8138 358634
rect -8694 322718 -8458 322954
rect -8374 322718 -8138 322954
rect -8694 322398 -8458 322634
rect -8374 322398 -8138 322634
rect -8694 286718 -8458 286954
rect -8374 286718 -8138 286954
rect -8694 286398 -8458 286634
rect -8374 286398 -8138 286634
rect -8694 250718 -8458 250954
rect -8374 250718 -8138 250954
rect -8694 250398 -8458 250634
rect -8374 250398 -8138 250634
rect -8694 214718 -8458 214954
rect -8374 214718 -8138 214954
rect -8694 214398 -8458 214634
rect -8374 214398 -8138 214634
rect -8694 178718 -8458 178954
rect -8374 178718 -8138 178954
rect -8694 178398 -8458 178634
rect -8374 178398 -8138 178634
rect -8694 142718 -8458 142954
rect -8374 142718 -8138 142954
rect -8694 142398 -8458 142634
rect -8374 142398 -8138 142634
rect -8694 106718 -8458 106954
rect -8374 106718 -8138 106954
rect -8694 106398 -8458 106634
rect -8374 106398 -8138 106634
rect -8694 70718 -8458 70954
rect -8374 70718 -8138 70954
rect -8694 70398 -8458 70634
rect -8374 70398 -8138 70634
rect -8694 34718 -8458 34954
rect -8374 34718 -8138 34954
rect -8694 34398 -8458 34634
rect -8374 34398 -8138 34634
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 678218 -7498 678454
rect -7414 678218 -7178 678454
rect -7734 677898 -7498 678134
rect -7414 677898 -7178 678134
rect -7734 642218 -7498 642454
rect -7414 642218 -7178 642454
rect -7734 641898 -7498 642134
rect -7414 641898 -7178 642134
rect -7734 606218 -7498 606454
rect -7414 606218 -7178 606454
rect -7734 605898 -7498 606134
rect -7414 605898 -7178 606134
rect -7734 570218 -7498 570454
rect -7414 570218 -7178 570454
rect -7734 569898 -7498 570134
rect -7414 569898 -7178 570134
rect -7734 534218 -7498 534454
rect -7414 534218 -7178 534454
rect -7734 533898 -7498 534134
rect -7414 533898 -7178 534134
rect -7734 498218 -7498 498454
rect -7414 498218 -7178 498454
rect -7734 497898 -7498 498134
rect -7414 497898 -7178 498134
rect -7734 462218 -7498 462454
rect -7414 462218 -7178 462454
rect -7734 461898 -7498 462134
rect -7414 461898 -7178 462134
rect -7734 426218 -7498 426454
rect -7414 426218 -7178 426454
rect -7734 425898 -7498 426134
rect -7414 425898 -7178 426134
rect -7734 390218 -7498 390454
rect -7414 390218 -7178 390454
rect -7734 389898 -7498 390134
rect -7414 389898 -7178 390134
rect -7734 354218 -7498 354454
rect -7414 354218 -7178 354454
rect -7734 353898 -7498 354134
rect -7414 353898 -7178 354134
rect -7734 318218 -7498 318454
rect -7414 318218 -7178 318454
rect -7734 317898 -7498 318134
rect -7414 317898 -7178 318134
rect -7734 282218 -7498 282454
rect -7414 282218 -7178 282454
rect -7734 281898 -7498 282134
rect -7414 281898 -7178 282134
rect -7734 246218 -7498 246454
rect -7414 246218 -7178 246454
rect -7734 245898 -7498 246134
rect -7414 245898 -7178 246134
rect -7734 210218 -7498 210454
rect -7414 210218 -7178 210454
rect -7734 209898 -7498 210134
rect -7414 209898 -7178 210134
rect -7734 174218 -7498 174454
rect -7414 174218 -7178 174454
rect -7734 173898 -7498 174134
rect -7414 173898 -7178 174134
rect -7734 138218 -7498 138454
rect -7414 138218 -7178 138454
rect -7734 137898 -7498 138134
rect -7414 137898 -7178 138134
rect -7734 102218 -7498 102454
rect -7414 102218 -7178 102454
rect -7734 101898 -7498 102134
rect -7414 101898 -7178 102134
rect -7734 66218 -7498 66454
rect -7414 66218 -7178 66454
rect -7734 65898 -7498 66134
rect -7414 65898 -7178 66134
rect -7734 30218 -7498 30454
rect -7414 30218 -7178 30454
rect -7734 29898 -7498 30134
rect -7414 29898 -7178 30134
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 673718 -6538 673954
rect -6454 673718 -6218 673954
rect -6774 673398 -6538 673634
rect -6454 673398 -6218 673634
rect -6774 637718 -6538 637954
rect -6454 637718 -6218 637954
rect -6774 637398 -6538 637634
rect -6454 637398 -6218 637634
rect -6774 601718 -6538 601954
rect -6454 601718 -6218 601954
rect -6774 601398 -6538 601634
rect -6454 601398 -6218 601634
rect -6774 565718 -6538 565954
rect -6454 565718 -6218 565954
rect -6774 565398 -6538 565634
rect -6454 565398 -6218 565634
rect -6774 529718 -6538 529954
rect -6454 529718 -6218 529954
rect -6774 529398 -6538 529634
rect -6454 529398 -6218 529634
rect -6774 493718 -6538 493954
rect -6454 493718 -6218 493954
rect -6774 493398 -6538 493634
rect -6454 493398 -6218 493634
rect -6774 457718 -6538 457954
rect -6454 457718 -6218 457954
rect -6774 457398 -6538 457634
rect -6454 457398 -6218 457634
rect -6774 421718 -6538 421954
rect -6454 421718 -6218 421954
rect -6774 421398 -6538 421634
rect -6454 421398 -6218 421634
rect -6774 385718 -6538 385954
rect -6454 385718 -6218 385954
rect -6774 385398 -6538 385634
rect -6454 385398 -6218 385634
rect -6774 349718 -6538 349954
rect -6454 349718 -6218 349954
rect -6774 349398 -6538 349634
rect -6454 349398 -6218 349634
rect -6774 313718 -6538 313954
rect -6454 313718 -6218 313954
rect -6774 313398 -6538 313634
rect -6454 313398 -6218 313634
rect -6774 277718 -6538 277954
rect -6454 277718 -6218 277954
rect -6774 277398 -6538 277634
rect -6454 277398 -6218 277634
rect -6774 241718 -6538 241954
rect -6454 241718 -6218 241954
rect -6774 241398 -6538 241634
rect -6454 241398 -6218 241634
rect -6774 205718 -6538 205954
rect -6454 205718 -6218 205954
rect -6774 205398 -6538 205634
rect -6454 205398 -6218 205634
rect -6774 169718 -6538 169954
rect -6454 169718 -6218 169954
rect -6774 169398 -6538 169634
rect -6454 169398 -6218 169634
rect -6774 133718 -6538 133954
rect -6454 133718 -6218 133954
rect -6774 133398 -6538 133634
rect -6454 133398 -6218 133634
rect -6774 97718 -6538 97954
rect -6454 97718 -6218 97954
rect -6774 97398 -6538 97634
rect -6454 97398 -6218 97634
rect -6774 61718 -6538 61954
rect -6454 61718 -6218 61954
rect -6774 61398 -6538 61634
rect -6454 61398 -6218 61634
rect -6774 25718 -6538 25954
rect -6454 25718 -6218 25954
rect -6774 25398 -6538 25634
rect -6454 25398 -6218 25634
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 669218 -5578 669454
rect -5494 669218 -5258 669454
rect -5814 668898 -5578 669134
rect -5494 668898 -5258 669134
rect -5814 633218 -5578 633454
rect -5494 633218 -5258 633454
rect -5814 632898 -5578 633134
rect -5494 632898 -5258 633134
rect -5814 597218 -5578 597454
rect -5494 597218 -5258 597454
rect -5814 596898 -5578 597134
rect -5494 596898 -5258 597134
rect -5814 561218 -5578 561454
rect -5494 561218 -5258 561454
rect -5814 560898 -5578 561134
rect -5494 560898 -5258 561134
rect -5814 525218 -5578 525454
rect -5494 525218 -5258 525454
rect -5814 524898 -5578 525134
rect -5494 524898 -5258 525134
rect -5814 489218 -5578 489454
rect -5494 489218 -5258 489454
rect -5814 488898 -5578 489134
rect -5494 488898 -5258 489134
rect -5814 453218 -5578 453454
rect -5494 453218 -5258 453454
rect -5814 452898 -5578 453134
rect -5494 452898 -5258 453134
rect -5814 417218 -5578 417454
rect -5494 417218 -5258 417454
rect -5814 416898 -5578 417134
rect -5494 416898 -5258 417134
rect -5814 381218 -5578 381454
rect -5494 381218 -5258 381454
rect -5814 380898 -5578 381134
rect -5494 380898 -5258 381134
rect -5814 345218 -5578 345454
rect -5494 345218 -5258 345454
rect -5814 344898 -5578 345134
rect -5494 344898 -5258 345134
rect -5814 309218 -5578 309454
rect -5494 309218 -5258 309454
rect -5814 308898 -5578 309134
rect -5494 308898 -5258 309134
rect -5814 273218 -5578 273454
rect -5494 273218 -5258 273454
rect -5814 272898 -5578 273134
rect -5494 272898 -5258 273134
rect -5814 237218 -5578 237454
rect -5494 237218 -5258 237454
rect -5814 236898 -5578 237134
rect -5494 236898 -5258 237134
rect -5814 201218 -5578 201454
rect -5494 201218 -5258 201454
rect -5814 200898 -5578 201134
rect -5494 200898 -5258 201134
rect -5814 165218 -5578 165454
rect -5494 165218 -5258 165454
rect -5814 164898 -5578 165134
rect -5494 164898 -5258 165134
rect -5814 129218 -5578 129454
rect -5494 129218 -5258 129454
rect -5814 128898 -5578 129134
rect -5494 128898 -5258 129134
rect -5814 93218 -5578 93454
rect -5494 93218 -5258 93454
rect -5814 92898 -5578 93134
rect -5494 92898 -5258 93134
rect -5814 57218 -5578 57454
rect -5494 57218 -5258 57454
rect -5814 56898 -5578 57134
rect -5494 56898 -5258 57134
rect -5814 21218 -5578 21454
rect -5494 21218 -5258 21454
rect -5814 20898 -5578 21134
rect -5494 20898 -5258 21134
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 700718 -4618 700954
rect -4534 700718 -4298 700954
rect -4854 700398 -4618 700634
rect -4534 700398 -4298 700634
rect -4854 664718 -4618 664954
rect -4534 664718 -4298 664954
rect -4854 664398 -4618 664634
rect -4534 664398 -4298 664634
rect -4854 628718 -4618 628954
rect -4534 628718 -4298 628954
rect -4854 628398 -4618 628634
rect -4534 628398 -4298 628634
rect -4854 592718 -4618 592954
rect -4534 592718 -4298 592954
rect -4854 592398 -4618 592634
rect -4534 592398 -4298 592634
rect -4854 556718 -4618 556954
rect -4534 556718 -4298 556954
rect -4854 556398 -4618 556634
rect -4534 556398 -4298 556634
rect -4854 520718 -4618 520954
rect -4534 520718 -4298 520954
rect -4854 520398 -4618 520634
rect -4534 520398 -4298 520634
rect -4854 484718 -4618 484954
rect -4534 484718 -4298 484954
rect -4854 484398 -4618 484634
rect -4534 484398 -4298 484634
rect -4854 448718 -4618 448954
rect -4534 448718 -4298 448954
rect -4854 448398 -4618 448634
rect -4534 448398 -4298 448634
rect -4854 412718 -4618 412954
rect -4534 412718 -4298 412954
rect -4854 412398 -4618 412634
rect -4534 412398 -4298 412634
rect -4854 376718 -4618 376954
rect -4534 376718 -4298 376954
rect -4854 376398 -4618 376634
rect -4534 376398 -4298 376634
rect -4854 340718 -4618 340954
rect -4534 340718 -4298 340954
rect -4854 340398 -4618 340634
rect -4534 340398 -4298 340634
rect -4854 304718 -4618 304954
rect -4534 304718 -4298 304954
rect -4854 304398 -4618 304634
rect -4534 304398 -4298 304634
rect -4854 268718 -4618 268954
rect -4534 268718 -4298 268954
rect -4854 268398 -4618 268634
rect -4534 268398 -4298 268634
rect -4854 232718 -4618 232954
rect -4534 232718 -4298 232954
rect -4854 232398 -4618 232634
rect -4534 232398 -4298 232634
rect -4854 196718 -4618 196954
rect -4534 196718 -4298 196954
rect -4854 196398 -4618 196634
rect -4534 196398 -4298 196634
rect -4854 160718 -4618 160954
rect -4534 160718 -4298 160954
rect -4854 160398 -4618 160634
rect -4534 160398 -4298 160634
rect -4854 124718 -4618 124954
rect -4534 124718 -4298 124954
rect -4854 124398 -4618 124634
rect -4534 124398 -4298 124634
rect -4854 88718 -4618 88954
rect -4534 88718 -4298 88954
rect -4854 88398 -4618 88634
rect -4534 88398 -4298 88634
rect -4854 52718 -4618 52954
rect -4534 52718 -4298 52954
rect -4854 52398 -4618 52634
rect -4534 52398 -4298 52634
rect -4854 16718 -4618 16954
rect -4534 16718 -4298 16954
rect -4854 16398 -4618 16634
rect -4534 16398 -4298 16634
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 696218 -3658 696454
rect -3574 696218 -3338 696454
rect -3894 695898 -3658 696134
rect -3574 695898 -3338 696134
rect -3894 660218 -3658 660454
rect -3574 660218 -3338 660454
rect -3894 659898 -3658 660134
rect -3574 659898 -3338 660134
rect -3894 624218 -3658 624454
rect -3574 624218 -3338 624454
rect -3894 623898 -3658 624134
rect -3574 623898 -3338 624134
rect -3894 588218 -3658 588454
rect -3574 588218 -3338 588454
rect -3894 587898 -3658 588134
rect -3574 587898 -3338 588134
rect -3894 552218 -3658 552454
rect -3574 552218 -3338 552454
rect -3894 551898 -3658 552134
rect -3574 551898 -3338 552134
rect -3894 516218 -3658 516454
rect -3574 516218 -3338 516454
rect -3894 515898 -3658 516134
rect -3574 515898 -3338 516134
rect -3894 480218 -3658 480454
rect -3574 480218 -3338 480454
rect -3894 479898 -3658 480134
rect -3574 479898 -3338 480134
rect -3894 444218 -3658 444454
rect -3574 444218 -3338 444454
rect -3894 443898 -3658 444134
rect -3574 443898 -3338 444134
rect -3894 408218 -3658 408454
rect -3574 408218 -3338 408454
rect -3894 407898 -3658 408134
rect -3574 407898 -3338 408134
rect -3894 372218 -3658 372454
rect -3574 372218 -3338 372454
rect -3894 371898 -3658 372134
rect -3574 371898 -3338 372134
rect -3894 336218 -3658 336454
rect -3574 336218 -3338 336454
rect -3894 335898 -3658 336134
rect -3574 335898 -3338 336134
rect -3894 300218 -3658 300454
rect -3574 300218 -3338 300454
rect -3894 299898 -3658 300134
rect -3574 299898 -3338 300134
rect -3894 264218 -3658 264454
rect -3574 264218 -3338 264454
rect -3894 263898 -3658 264134
rect -3574 263898 -3338 264134
rect -3894 228218 -3658 228454
rect -3574 228218 -3338 228454
rect -3894 227898 -3658 228134
rect -3574 227898 -3338 228134
rect -3894 192218 -3658 192454
rect -3574 192218 -3338 192454
rect -3894 191898 -3658 192134
rect -3574 191898 -3338 192134
rect -3894 156218 -3658 156454
rect -3574 156218 -3338 156454
rect -3894 155898 -3658 156134
rect -3574 155898 -3338 156134
rect -3894 120218 -3658 120454
rect -3574 120218 -3338 120454
rect -3894 119898 -3658 120134
rect -3574 119898 -3338 120134
rect -3894 84218 -3658 84454
rect -3574 84218 -3338 84454
rect -3894 83898 -3658 84134
rect -3574 83898 -3338 84134
rect -3894 48218 -3658 48454
rect -3574 48218 -3338 48454
rect -3894 47898 -3658 48134
rect -3574 47898 -3338 48134
rect -3894 12218 -3658 12454
rect -3574 12218 -3338 12454
rect -3894 11898 -3658 12134
rect -3574 11898 -3338 12134
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 691718 -2698 691954
rect -2614 691718 -2378 691954
rect -2934 691398 -2698 691634
rect -2614 691398 -2378 691634
rect -2934 655718 -2698 655954
rect -2614 655718 -2378 655954
rect -2934 655398 -2698 655634
rect -2614 655398 -2378 655634
rect -2934 619718 -2698 619954
rect -2614 619718 -2378 619954
rect -2934 619398 -2698 619634
rect -2614 619398 -2378 619634
rect -2934 583718 -2698 583954
rect -2614 583718 -2378 583954
rect -2934 583398 -2698 583634
rect -2614 583398 -2378 583634
rect -2934 547718 -2698 547954
rect -2614 547718 -2378 547954
rect -2934 547398 -2698 547634
rect -2614 547398 -2378 547634
rect -2934 511718 -2698 511954
rect -2614 511718 -2378 511954
rect -2934 511398 -2698 511634
rect -2614 511398 -2378 511634
rect -2934 475718 -2698 475954
rect -2614 475718 -2378 475954
rect -2934 475398 -2698 475634
rect -2614 475398 -2378 475634
rect -2934 439718 -2698 439954
rect -2614 439718 -2378 439954
rect -2934 439398 -2698 439634
rect -2614 439398 -2378 439634
rect -2934 403718 -2698 403954
rect -2614 403718 -2378 403954
rect -2934 403398 -2698 403634
rect -2614 403398 -2378 403634
rect -2934 367718 -2698 367954
rect -2614 367718 -2378 367954
rect -2934 367398 -2698 367634
rect -2614 367398 -2378 367634
rect -2934 331718 -2698 331954
rect -2614 331718 -2378 331954
rect -2934 331398 -2698 331634
rect -2614 331398 -2378 331634
rect -2934 295718 -2698 295954
rect -2614 295718 -2378 295954
rect -2934 295398 -2698 295634
rect -2614 295398 -2378 295634
rect -2934 259718 -2698 259954
rect -2614 259718 -2378 259954
rect -2934 259398 -2698 259634
rect -2614 259398 -2378 259634
rect -2934 223718 -2698 223954
rect -2614 223718 -2378 223954
rect -2934 223398 -2698 223634
rect -2614 223398 -2378 223634
rect -2934 187718 -2698 187954
rect -2614 187718 -2378 187954
rect -2934 187398 -2698 187634
rect -2614 187398 -2378 187634
rect -2934 151718 -2698 151954
rect -2614 151718 -2378 151954
rect -2934 151398 -2698 151634
rect -2614 151398 -2378 151634
rect -2934 115718 -2698 115954
rect -2614 115718 -2378 115954
rect -2934 115398 -2698 115634
rect -2614 115398 -2378 115634
rect -2934 79718 -2698 79954
rect -2614 79718 -2378 79954
rect -2934 79398 -2698 79634
rect -2614 79398 -2378 79634
rect -2934 43718 -2698 43954
rect -2614 43718 -2378 43954
rect -2934 43398 -2698 43634
rect -2614 43398 -2378 43634
rect -2934 7718 -2698 7954
rect -2614 7718 -2378 7954
rect -2934 7398 -2698 7634
rect -2614 7398 -2378 7634
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 6326 705562 6562 705798
rect 6646 705562 6882 705798
rect 6326 705242 6562 705478
rect 6646 705242 6882 705478
rect 6326 691718 6562 691954
rect 6646 691718 6882 691954
rect 6326 691398 6562 691634
rect 6646 691398 6882 691634
rect 6326 655718 6562 655954
rect 6646 655718 6882 655954
rect 6326 655398 6562 655634
rect 6646 655398 6882 655634
rect 6326 619718 6562 619954
rect 6646 619718 6882 619954
rect 6326 619398 6562 619634
rect 6646 619398 6882 619634
rect 6326 583718 6562 583954
rect 6646 583718 6882 583954
rect 6326 583398 6562 583634
rect 6646 583398 6882 583634
rect 6326 547718 6562 547954
rect 6646 547718 6882 547954
rect 6326 547398 6562 547634
rect 6646 547398 6882 547634
rect 6326 511718 6562 511954
rect 6646 511718 6882 511954
rect 6326 511398 6562 511634
rect 6646 511398 6882 511634
rect 6326 475718 6562 475954
rect 6646 475718 6882 475954
rect 6326 475398 6562 475634
rect 6646 475398 6882 475634
rect 6326 439718 6562 439954
rect 6646 439718 6882 439954
rect 6326 439398 6562 439634
rect 6646 439398 6882 439634
rect 6326 403718 6562 403954
rect 6646 403718 6882 403954
rect 6326 403398 6562 403634
rect 6646 403398 6882 403634
rect 6326 367718 6562 367954
rect 6646 367718 6882 367954
rect 6326 367398 6562 367634
rect 6646 367398 6882 367634
rect 6326 331718 6562 331954
rect 6646 331718 6882 331954
rect 6326 331398 6562 331634
rect 6646 331398 6882 331634
rect 6326 295718 6562 295954
rect 6646 295718 6882 295954
rect 6326 295398 6562 295634
rect 6646 295398 6882 295634
rect 6326 259718 6562 259954
rect 6646 259718 6882 259954
rect 6326 259398 6562 259634
rect 6646 259398 6882 259634
rect 6326 223718 6562 223954
rect 6646 223718 6882 223954
rect 6326 223398 6562 223634
rect 6646 223398 6882 223634
rect 6326 187718 6562 187954
rect 6646 187718 6882 187954
rect 6326 187398 6562 187634
rect 6646 187398 6882 187634
rect 6326 151718 6562 151954
rect 6646 151718 6882 151954
rect 6326 151398 6562 151634
rect 6646 151398 6882 151634
rect 6326 115718 6562 115954
rect 6646 115718 6882 115954
rect 6326 115398 6562 115634
rect 6646 115398 6882 115634
rect 6326 79718 6562 79954
rect 6646 79718 6882 79954
rect 6326 79398 6562 79634
rect 6646 79398 6882 79634
rect 6326 43718 6562 43954
rect 6646 43718 6882 43954
rect 6326 43398 6562 43634
rect 6646 43398 6882 43634
rect 6326 7718 6562 7954
rect 6646 7718 6882 7954
rect 6326 7398 6562 7634
rect 6646 7398 6882 7634
rect 6326 -1542 6562 -1306
rect 6646 -1542 6882 -1306
rect 6326 -1862 6562 -1626
rect 6646 -1862 6882 -1626
rect 10826 706522 11062 706758
rect 11146 706522 11382 706758
rect 10826 706202 11062 706438
rect 11146 706202 11382 706438
rect 10826 696218 11062 696454
rect 11146 696218 11382 696454
rect 10826 695898 11062 696134
rect 11146 695898 11382 696134
rect 10826 660218 11062 660454
rect 11146 660218 11382 660454
rect 10826 659898 11062 660134
rect 11146 659898 11382 660134
rect 10826 624218 11062 624454
rect 11146 624218 11382 624454
rect 10826 623898 11062 624134
rect 11146 623898 11382 624134
rect 10826 588218 11062 588454
rect 11146 588218 11382 588454
rect 10826 587898 11062 588134
rect 11146 587898 11382 588134
rect 10826 552218 11062 552454
rect 11146 552218 11382 552454
rect 10826 551898 11062 552134
rect 11146 551898 11382 552134
rect 10826 516218 11062 516454
rect 11146 516218 11382 516454
rect 10826 515898 11062 516134
rect 11146 515898 11382 516134
rect 10826 480218 11062 480454
rect 11146 480218 11382 480454
rect 10826 479898 11062 480134
rect 11146 479898 11382 480134
rect 10826 444218 11062 444454
rect 11146 444218 11382 444454
rect 10826 443898 11062 444134
rect 11146 443898 11382 444134
rect 10826 408218 11062 408454
rect 11146 408218 11382 408454
rect 10826 407898 11062 408134
rect 11146 407898 11382 408134
rect 10826 372218 11062 372454
rect 11146 372218 11382 372454
rect 10826 371898 11062 372134
rect 11146 371898 11382 372134
rect 10826 336218 11062 336454
rect 11146 336218 11382 336454
rect 10826 335898 11062 336134
rect 11146 335898 11382 336134
rect 10826 300218 11062 300454
rect 11146 300218 11382 300454
rect 10826 299898 11062 300134
rect 11146 299898 11382 300134
rect 10826 264218 11062 264454
rect 11146 264218 11382 264454
rect 10826 263898 11062 264134
rect 11146 263898 11382 264134
rect 10826 228218 11062 228454
rect 11146 228218 11382 228454
rect 10826 227898 11062 228134
rect 11146 227898 11382 228134
rect 10826 192218 11062 192454
rect 11146 192218 11382 192454
rect 10826 191898 11062 192134
rect 11146 191898 11382 192134
rect 10826 156218 11062 156454
rect 11146 156218 11382 156454
rect 10826 155898 11062 156134
rect 11146 155898 11382 156134
rect 10826 120218 11062 120454
rect 11146 120218 11382 120454
rect 10826 119898 11062 120134
rect 11146 119898 11382 120134
rect 10826 84218 11062 84454
rect 11146 84218 11382 84454
rect 10826 83898 11062 84134
rect 11146 83898 11382 84134
rect 10826 48218 11062 48454
rect 11146 48218 11382 48454
rect 10826 47898 11062 48134
rect 11146 47898 11382 48134
rect 10826 12218 11062 12454
rect 11146 12218 11382 12454
rect 10826 11898 11062 12134
rect 11146 11898 11382 12134
rect 10826 -2502 11062 -2266
rect 11146 -2502 11382 -2266
rect 10826 -2822 11062 -2586
rect 11146 -2822 11382 -2586
rect 15326 707482 15562 707718
rect 15646 707482 15882 707718
rect 15326 707162 15562 707398
rect 15646 707162 15882 707398
rect 15326 700718 15562 700954
rect 15646 700718 15882 700954
rect 15326 700398 15562 700634
rect 15646 700398 15882 700634
rect 15326 664718 15562 664954
rect 15646 664718 15882 664954
rect 15326 664398 15562 664634
rect 15646 664398 15882 664634
rect 15326 628718 15562 628954
rect 15646 628718 15882 628954
rect 15326 628398 15562 628634
rect 15646 628398 15882 628634
rect 15326 592718 15562 592954
rect 15646 592718 15882 592954
rect 15326 592398 15562 592634
rect 15646 592398 15882 592634
rect 15326 556718 15562 556954
rect 15646 556718 15882 556954
rect 15326 556398 15562 556634
rect 15646 556398 15882 556634
rect 15326 520718 15562 520954
rect 15646 520718 15882 520954
rect 15326 520398 15562 520634
rect 15646 520398 15882 520634
rect 15326 484718 15562 484954
rect 15646 484718 15882 484954
rect 15326 484398 15562 484634
rect 15646 484398 15882 484634
rect 15326 448718 15562 448954
rect 15646 448718 15882 448954
rect 15326 448398 15562 448634
rect 15646 448398 15882 448634
rect 15326 412718 15562 412954
rect 15646 412718 15882 412954
rect 15326 412398 15562 412634
rect 15646 412398 15882 412634
rect 15326 376718 15562 376954
rect 15646 376718 15882 376954
rect 15326 376398 15562 376634
rect 15646 376398 15882 376634
rect 15326 340718 15562 340954
rect 15646 340718 15882 340954
rect 15326 340398 15562 340634
rect 15646 340398 15882 340634
rect 15326 304718 15562 304954
rect 15646 304718 15882 304954
rect 15326 304398 15562 304634
rect 15646 304398 15882 304634
rect 15326 268718 15562 268954
rect 15646 268718 15882 268954
rect 15326 268398 15562 268634
rect 15646 268398 15882 268634
rect 15326 232718 15562 232954
rect 15646 232718 15882 232954
rect 15326 232398 15562 232634
rect 15646 232398 15882 232634
rect 15326 196718 15562 196954
rect 15646 196718 15882 196954
rect 15326 196398 15562 196634
rect 15646 196398 15882 196634
rect 15326 160718 15562 160954
rect 15646 160718 15882 160954
rect 15326 160398 15562 160634
rect 15646 160398 15882 160634
rect 15326 124718 15562 124954
rect 15646 124718 15882 124954
rect 15326 124398 15562 124634
rect 15646 124398 15882 124634
rect 15326 88718 15562 88954
rect 15646 88718 15882 88954
rect 15326 88398 15562 88634
rect 15646 88398 15882 88634
rect 15326 52718 15562 52954
rect 15646 52718 15882 52954
rect 15326 52398 15562 52634
rect 15646 52398 15882 52634
rect 15326 16718 15562 16954
rect 15646 16718 15882 16954
rect 15326 16398 15562 16634
rect 15646 16398 15882 16634
rect 15326 -3462 15562 -3226
rect 15646 -3462 15882 -3226
rect 15326 -3782 15562 -3546
rect 15646 -3782 15882 -3546
rect 19826 708442 20062 708678
rect 20146 708442 20382 708678
rect 19826 708122 20062 708358
rect 20146 708122 20382 708358
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -4422 20062 -4186
rect 20146 -4422 20382 -4186
rect 19826 -4742 20062 -4506
rect 20146 -4742 20382 -4506
rect 24326 709402 24562 709638
rect 24646 709402 24882 709638
rect 24326 709082 24562 709318
rect 24646 709082 24882 709318
rect 24326 673718 24562 673954
rect 24646 673718 24882 673954
rect 24326 673398 24562 673634
rect 24646 673398 24882 673634
rect 24326 637718 24562 637954
rect 24646 637718 24882 637954
rect 24326 637398 24562 637634
rect 24646 637398 24882 637634
rect 24326 601718 24562 601954
rect 24646 601718 24882 601954
rect 24326 601398 24562 601634
rect 24646 601398 24882 601634
rect 24326 565718 24562 565954
rect 24646 565718 24882 565954
rect 24326 565398 24562 565634
rect 24646 565398 24882 565634
rect 24326 529718 24562 529954
rect 24646 529718 24882 529954
rect 24326 529398 24562 529634
rect 24646 529398 24882 529634
rect 24326 493718 24562 493954
rect 24646 493718 24882 493954
rect 24326 493398 24562 493634
rect 24646 493398 24882 493634
rect 24326 457718 24562 457954
rect 24646 457718 24882 457954
rect 24326 457398 24562 457634
rect 24646 457398 24882 457634
rect 24326 421718 24562 421954
rect 24646 421718 24882 421954
rect 24326 421398 24562 421634
rect 24646 421398 24882 421634
rect 24326 385718 24562 385954
rect 24646 385718 24882 385954
rect 24326 385398 24562 385634
rect 24646 385398 24882 385634
rect 24326 349718 24562 349954
rect 24646 349718 24882 349954
rect 24326 349398 24562 349634
rect 24646 349398 24882 349634
rect 24326 313718 24562 313954
rect 24646 313718 24882 313954
rect 24326 313398 24562 313634
rect 24646 313398 24882 313634
rect 24326 277718 24562 277954
rect 24646 277718 24882 277954
rect 24326 277398 24562 277634
rect 24646 277398 24882 277634
rect 24326 241718 24562 241954
rect 24646 241718 24882 241954
rect 24326 241398 24562 241634
rect 24646 241398 24882 241634
rect 24326 205718 24562 205954
rect 24646 205718 24882 205954
rect 24326 205398 24562 205634
rect 24646 205398 24882 205634
rect 24326 169718 24562 169954
rect 24646 169718 24882 169954
rect 24326 169398 24562 169634
rect 24646 169398 24882 169634
rect 24326 133718 24562 133954
rect 24646 133718 24882 133954
rect 24326 133398 24562 133634
rect 24646 133398 24882 133634
rect 24326 97718 24562 97954
rect 24646 97718 24882 97954
rect 24326 97398 24562 97634
rect 24646 97398 24882 97634
rect 24326 61718 24562 61954
rect 24646 61718 24882 61954
rect 24326 61398 24562 61634
rect 24646 61398 24882 61634
rect 24326 25718 24562 25954
rect 24646 25718 24882 25954
rect 24326 25398 24562 25634
rect 24646 25398 24882 25634
rect 24326 -5382 24562 -5146
rect 24646 -5382 24882 -5146
rect 24326 -5702 24562 -5466
rect 24646 -5702 24882 -5466
rect 28826 710362 29062 710598
rect 29146 710362 29382 710598
rect 28826 710042 29062 710278
rect 29146 710042 29382 710278
rect 28826 678218 29062 678454
rect 29146 678218 29382 678454
rect 28826 677898 29062 678134
rect 29146 677898 29382 678134
rect 28826 642218 29062 642454
rect 29146 642218 29382 642454
rect 28826 641898 29062 642134
rect 29146 641898 29382 642134
rect 28826 606218 29062 606454
rect 29146 606218 29382 606454
rect 28826 605898 29062 606134
rect 29146 605898 29382 606134
rect 28826 570218 29062 570454
rect 29146 570218 29382 570454
rect 28826 569898 29062 570134
rect 29146 569898 29382 570134
rect 28826 534218 29062 534454
rect 29146 534218 29382 534454
rect 28826 533898 29062 534134
rect 29146 533898 29382 534134
rect 28826 498218 29062 498454
rect 29146 498218 29382 498454
rect 28826 497898 29062 498134
rect 29146 497898 29382 498134
rect 28826 462218 29062 462454
rect 29146 462218 29382 462454
rect 28826 461898 29062 462134
rect 29146 461898 29382 462134
rect 28826 426218 29062 426454
rect 29146 426218 29382 426454
rect 28826 425898 29062 426134
rect 29146 425898 29382 426134
rect 28826 390218 29062 390454
rect 29146 390218 29382 390454
rect 28826 389898 29062 390134
rect 29146 389898 29382 390134
rect 28826 354218 29062 354454
rect 29146 354218 29382 354454
rect 28826 353898 29062 354134
rect 29146 353898 29382 354134
rect 28826 318218 29062 318454
rect 29146 318218 29382 318454
rect 28826 317898 29062 318134
rect 29146 317898 29382 318134
rect 28826 282218 29062 282454
rect 29146 282218 29382 282454
rect 28826 281898 29062 282134
rect 29146 281898 29382 282134
rect 28826 246218 29062 246454
rect 29146 246218 29382 246454
rect 28826 245898 29062 246134
rect 29146 245898 29382 246134
rect 28826 210218 29062 210454
rect 29146 210218 29382 210454
rect 28826 209898 29062 210134
rect 29146 209898 29382 210134
rect 28826 174218 29062 174454
rect 29146 174218 29382 174454
rect 28826 173898 29062 174134
rect 29146 173898 29382 174134
rect 28826 138218 29062 138454
rect 29146 138218 29382 138454
rect 28826 137898 29062 138134
rect 29146 137898 29382 138134
rect 28826 102218 29062 102454
rect 29146 102218 29382 102454
rect 28826 101898 29062 102134
rect 29146 101898 29382 102134
rect 28826 66218 29062 66454
rect 29146 66218 29382 66454
rect 28826 65898 29062 66134
rect 29146 65898 29382 66134
rect 28826 30218 29062 30454
rect 29146 30218 29382 30454
rect 28826 29898 29062 30134
rect 29146 29898 29382 30134
rect 28826 -6342 29062 -6106
rect 29146 -6342 29382 -6106
rect 28826 -6662 29062 -6426
rect 29146 -6662 29382 -6426
rect 33326 711322 33562 711558
rect 33646 711322 33882 711558
rect 33326 711002 33562 711238
rect 33646 711002 33882 711238
rect 33326 682718 33562 682954
rect 33646 682718 33882 682954
rect 33326 682398 33562 682634
rect 33646 682398 33882 682634
rect 33326 646718 33562 646954
rect 33646 646718 33882 646954
rect 33326 646398 33562 646634
rect 33646 646398 33882 646634
rect 33326 610718 33562 610954
rect 33646 610718 33882 610954
rect 33326 610398 33562 610634
rect 33646 610398 33882 610634
rect 33326 574718 33562 574954
rect 33646 574718 33882 574954
rect 33326 574398 33562 574634
rect 33646 574398 33882 574634
rect 33326 538718 33562 538954
rect 33646 538718 33882 538954
rect 33326 538398 33562 538634
rect 33646 538398 33882 538634
rect 33326 502718 33562 502954
rect 33646 502718 33882 502954
rect 33326 502398 33562 502634
rect 33646 502398 33882 502634
rect 33326 466718 33562 466954
rect 33646 466718 33882 466954
rect 33326 466398 33562 466634
rect 33646 466398 33882 466634
rect 33326 430718 33562 430954
rect 33646 430718 33882 430954
rect 33326 430398 33562 430634
rect 33646 430398 33882 430634
rect 33326 394718 33562 394954
rect 33646 394718 33882 394954
rect 33326 394398 33562 394634
rect 33646 394398 33882 394634
rect 33326 358718 33562 358954
rect 33646 358718 33882 358954
rect 33326 358398 33562 358634
rect 33646 358398 33882 358634
rect 33326 322718 33562 322954
rect 33646 322718 33882 322954
rect 33326 322398 33562 322634
rect 33646 322398 33882 322634
rect 33326 286718 33562 286954
rect 33646 286718 33882 286954
rect 33326 286398 33562 286634
rect 33646 286398 33882 286634
rect 33326 250718 33562 250954
rect 33646 250718 33882 250954
rect 33326 250398 33562 250634
rect 33646 250398 33882 250634
rect 33326 214718 33562 214954
rect 33646 214718 33882 214954
rect 33326 214398 33562 214634
rect 33646 214398 33882 214634
rect 33326 178718 33562 178954
rect 33646 178718 33882 178954
rect 33326 178398 33562 178634
rect 33646 178398 33882 178634
rect 33326 142718 33562 142954
rect 33646 142718 33882 142954
rect 33326 142398 33562 142634
rect 33646 142398 33882 142634
rect 33326 106718 33562 106954
rect 33646 106718 33882 106954
rect 33326 106398 33562 106634
rect 33646 106398 33882 106634
rect 33326 70718 33562 70954
rect 33646 70718 33882 70954
rect 33326 70398 33562 70634
rect 33646 70398 33882 70634
rect 33326 34718 33562 34954
rect 33646 34718 33882 34954
rect 33326 34398 33562 34634
rect 33646 34398 33882 34634
rect 33326 -7302 33562 -7066
rect 33646 -7302 33882 -7066
rect 33326 -7622 33562 -7386
rect 33646 -7622 33882 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 42326 705562 42562 705798
rect 42646 705562 42882 705798
rect 42326 705242 42562 705478
rect 42646 705242 42882 705478
rect 42326 691718 42562 691954
rect 42646 691718 42882 691954
rect 42326 691398 42562 691634
rect 42646 691398 42882 691634
rect 42326 655718 42562 655954
rect 42646 655718 42882 655954
rect 42326 655398 42562 655634
rect 42646 655398 42882 655634
rect 42326 619718 42562 619954
rect 42646 619718 42882 619954
rect 42326 619398 42562 619634
rect 42646 619398 42882 619634
rect 42326 583718 42562 583954
rect 42646 583718 42882 583954
rect 42326 583398 42562 583634
rect 42646 583398 42882 583634
rect 42326 547718 42562 547954
rect 42646 547718 42882 547954
rect 42326 547398 42562 547634
rect 42646 547398 42882 547634
rect 42326 511718 42562 511954
rect 42646 511718 42882 511954
rect 42326 511398 42562 511634
rect 42646 511398 42882 511634
rect 42326 475718 42562 475954
rect 42646 475718 42882 475954
rect 42326 475398 42562 475634
rect 42646 475398 42882 475634
rect 42326 439718 42562 439954
rect 42646 439718 42882 439954
rect 42326 439398 42562 439634
rect 42646 439398 42882 439634
rect 42326 403718 42562 403954
rect 42646 403718 42882 403954
rect 42326 403398 42562 403634
rect 42646 403398 42882 403634
rect 42326 367718 42562 367954
rect 42646 367718 42882 367954
rect 42326 367398 42562 367634
rect 42646 367398 42882 367634
rect 42326 331718 42562 331954
rect 42646 331718 42882 331954
rect 42326 331398 42562 331634
rect 42646 331398 42882 331634
rect 42326 295718 42562 295954
rect 42646 295718 42882 295954
rect 42326 295398 42562 295634
rect 42646 295398 42882 295634
rect 42326 259718 42562 259954
rect 42646 259718 42882 259954
rect 42326 259398 42562 259634
rect 42646 259398 42882 259634
rect 42326 223718 42562 223954
rect 42646 223718 42882 223954
rect 42326 223398 42562 223634
rect 42646 223398 42882 223634
rect 42326 187718 42562 187954
rect 42646 187718 42882 187954
rect 42326 187398 42562 187634
rect 42646 187398 42882 187634
rect 42326 151718 42562 151954
rect 42646 151718 42882 151954
rect 42326 151398 42562 151634
rect 42646 151398 42882 151634
rect 42326 115718 42562 115954
rect 42646 115718 42882 115954
rect 42326 115398 42562 115634
rect 42646 115398 42882 115634
rect 42326 79718 42562 79954
rect 42646 79718 42882 79954
rect 42326 79398 42562 79634
rect 42646 79398 42882 79634
rect 42326 43718 42562 43954
rect 42646 43718 42882 43954
rect 42326 43398 42562 43634
rect 42646 43398 42882 43634
rect 42326 7718 42562 7954
rect 42646 7718 42882 7954
rect 42326 7398 42562 7634
rect 42646 7398 42882 7634
rect 42326 -1542 42562 -1306
rect 42646 -1542 42882 -1306
rect 42326 -1862 42562 -1626
rect 42646 -1862 42882 -1626
rect 46826 706522 47062 706758
rect 47146 706522 47382 706758
rect 46826 706202 47062 706438
rect 47146 706202 47382 706438
rect 46826 696218 47062 696454
rect 47146 696218 47382 696454
rect 46826 695898 47062 696134
rect 47146 695898 47382 696134
rect 46826 660218 47062 660454
rect 47146 660218 47382 660454
rect 46826 659898 47062 660134
rect 47146 659898 47382 660134
rect 46826 624218 47062 624454
rect 47146 624218 47382 624454
rect 46826 623898 47062 624134
rect 47146 623898 47382 624134
rect 46826 588218 47062 588454
rect 47146 588218 47382 588454
rect 46826 587898 47062 588134
rect 47146 587898 47382 588134
rect 46826 552218 47062 552454
rect 47146 552218 47382 552454
rect 46826 551898 47062 552134
rect 47146 551898 47382 552134
rect 46826 516218 47062 516454
rect 47146 516218 47382 516454
rect 46826 515898 47062 516134
rect 47146 515898 47382 516134
rect 46826 480218 47062 480454
rect 47146 480218 47382 480454
rect 46826 479898 47062 480134
rect 47146 479898 47382 480134
rect 46826 444218 47062 444454
rect 47146 444218 47382 444454
rect 46826 443898 47062 444134
rect 47146 443898 47382 444134
rect 46826 408218 47062 408454
rect 47146 408218 47382 408454
rect 46826 407898 47062 408134
rect 47146 407898 47382 408134
rect 46826 372218 47062 372454
rect 47146 372218 47382 372454
rect 46826 371898 47062 372134
rect 47146 371898 47382 372134
rect 46826 336218 47062 336454
rect 47146 336218 47382 336454
rect 46826 335898 47062 336134
rect 47146 335898 47382 336134
rect 46826 300218 47062 300454
rect 47146 300218 47382 300454
rect 46826 299898 47062 300134
rect 47146 299898 47382 300134
rect 46826 264218 47062 264454
rect 47146 264218 47382 264454
rect 46826 263898 47062 264134
rect 47146 263898 47382 264134
rect 46826 228218 47062 228454
rect 47146 228218 47382 228454
rect 46826 227898 47062 228134
rect 47146 227898 47382 228134
rect 46826 192218 47062 192454
rect 47146 192218 47382 192454
rect 46826 191898 47062 192134
rect 47146 191898 47382 192134
rect 46826 156218 47062 156454
rect 47146 156218 47382 156454
rect 46826 155898 47062 156134
rect 47146 155898 47382 156134
rect 46826 120218 47062 120454
rect 47146 120218 47382 120454
rect 46826 119898 47062 120134
rect 47146 119898 47382 120134
rect 46826 84218 47062 84454
rect 47146 84218 47382 84454
rect 46826 83898 47062 84134
rect 47146 83898 47382 84134
rect 46826 48218 47062 48454
rect 47146 48218 47382 48454
rect 46826 47898 47062 48134
rect 47146 47898 47382 48134
rect 46826 12218 47062 12454
rect 47146 12218 47382 12454
rect 46826 11898 47062 12134
rect 47146 11898 47382 12134
rect 46826 -2502 47062 -2266
rect 47146 -2502 47382 -2266
rect 46826 -2822 47062 -2586
rect 47146 -2822 47382 -2586
rect 51326 707482 51562 707718
rect 51646 707482 51882 707718
rect 51326 707162 51562 707398
rect 51646 707162 51882 707398
rect 51326 700718 51562 700954
rect 51646 700718 51882 700954
rect 51326 700398 51562 700634
rect 51646 700398 51882 700634
rect 51326 664718 51562 664954
rect 51646 664718 51882 664954
rect 51326 664398 51562 664634
rect 51646 664398 51882 664634
rect 51326 628718 51562 628954
rect 51646 628718 51882 628954
rect 51326 628398 51562 628634
rect 51646 628398 51882 628634
rect 51326 592718 51562 592954
rect 51646 592718 51882 592954
rect 51326 592398 51562 592634
rect 51646 592398 51882 592634
rect 51326 556718 51562 556954
rect 51646 556718 51882 556954
rect 51326 556398 51562 556634
rect 51646 556398 51882 556634
rect 51326 520718 51562 520954
rect 51646 520718 51882 520954
rect 51326 520398 51562 520634
rect 51646 520398 51882 520634
rect 51326 484718 51562 484954
rect 51646 484718 51882 484954
rect 51326 484398 51562 484634
rect 51646 484398 51882 484634
rect 51326 448718 51562 448954
rect 51646 448718 51882 448954
rect 51326 448398 51562 448634
rect 51646 448398 51882 448634
rect 51326 412718 51562 412954
rect 51646 412718 51882 412954
rect 51326 412398 51562 412634
rect 51646 412398 51882 412634
rect 51326 376718 51562 376954
rect 51646 376718 51882 376954
rect 51326 376398 51562 376634
rect 51646 376398 51882 376634
rect 51326 340718 51562 340954
rect 51646 340718 51882 340954
rect 51326 340398 51562 340634
rect 51646 340398 51882 340634
rect 51326 304718 51562 304954
rect 51646 304718 51882 304954
rect 51326 304398 51562 304634
rect 51646 304398 51882 304634
rect 51326 268718 51562 268954
rect 51646 268718 51882 268954
rect 51326 268398 51562 268634
rect 51646 268398 51882 268634
rect 51326 232718 51562 232954
rect 51646 232718 51882 232954
rect 51326 232398 51562 232634
rect 51646 232398 51882 232634
rect 51326 196718 51562 196954
rect 51646 196718 51882 196954
rect 51326 196398 51562 196634
rect 51646 196398 51882 196634
rect 51326 160718 51562 160954
rect 51646 160718 51882 160954
rect 51326 160398 51562 160634
rect 51646 160398 51882 160634
rect 51326 124718 51562 124954
rect 51646 124718 51882 124954
rect 51326 124398 51562 124634
rect 51646 124398 51882 124634
rect 51326 88718 51562 88954
rect 51646 88718 51882 88954
rect 51326 88398 51562 88634
rect 51646 88398 51882 88634
rect 51326 52718 51562 52954
rect 51646 52718 51882 52954
rect 51326 52398 51562 52634
rect 51646 52398 51882 52634
rect 51326 16718 51562 16954
rect 51646 16718 51882 16954
rect 51326 16398 51562 16634
rect 51646 16398 51882 16634
rect 51326 -3462 51562 -3226
rect 51646 -3462 51882 -3226
rect 51326 -3782 51562 -3546
rect 51646 -3782 51882 -3546
rect 55826 708442 56062 708678
rect 56146 708442 56382 708678
rect 55826 708122 56062 708358
rect 56146 708122 56382 708358
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -4422 56062 -4186
rect 56146 -4422 56382 -4186
rect 55826 -4742 56062 -4506
rect 56146 -4742 56382 -4506
rect 60326 709402 60562 709638
rect 60646 709402 60882 709638
rect 60326 709082 60562 709318
rect 60646 709082 60882 709318
rect 60326 673718 60562 673954
rect 60646 673718 60882 673954
rect 60326 673398 60562 673634
rect 60646 673398 60882 673634
rect 60326 637718 60562 637954
rect 60646 637718 60882 637954
rect 60326 637398 60562 637634
rect 60646 637398 60882 637634
rect 60326 601718 60562 601954
rect 60646 601718 60882 601954
rect 60326 601398 60562 601634
rect 60646 601398 60882 601634
rect 60326 565718 60562 565954
rect 60646 565718 60882 565954
rect 60326 565398 60562 565634
rect 60646 565398 60882 565634
rect 60326 529718 60562 529954
rect 60646 529718 60882 529954
rect 60326 529398 60562 529634
rect 60646 529398 60882 529634
rect 60326 493718 60562 493954
rect 60646 493718 60882 493954
rect 60326 493398 60562 493634
rect 60646 493398 60882 493634
rect 60326 457718 60562 457954
rect 60646 457718 60882 457954
rect 60326 457398 60562 457634
rect 60646 457398 60882 457634
rect 60326 421718 60562 421954
rect 60646 421718 60882 421954
rect 60326 421398 60562 421634
rect 60646 421398 60882 421634
rect 60326 385718 60562 385954
rect 60646 385718 60882 385954
rect 60326 385398 60562 385634
rect 60646 385398 60882 385634
rect 60326 349718 60562 349954
rect 60646 349718 60882 349954
rect 60326 349398 60562 349634
rect 60646 349398 60882 349634
rect 60326 313718 60562 313954
rect 60646 313718 60882 313954
rect 60326 313398 60562 313634
rect 60646 313398 60882 313634
rect 60326 277718 60562 277954
rect 60646 277718 60882 277954
rect 60326 277398 60562 277634
rect 60646 277398 60882 277634
rect 60326 241718 60562 241954
rect 60646 241718 60882 241954
rect 60326 241398 60562 241634
rect 60646 241398 60882 241634
rect 60326 205718 60562 205954
rect 60646 205718 60882 205954
rect 60326 205398 60562 205634
rect 60646 205398 60882 205634
rect 60326 169718 60562 169954
rect 60646 169718 60882 169954
rect 60326 169398 60562 169634
rect 60646 169398 60882 169634
rect 60326 133718 60562 133954
rect 60646 133718 60882 133954
rect 60326 133398 60562 133634
rect 60646 133398 60882 133634
rect 60326 97718 60562 97954
rect 60646 97718 60882 97954
rect 60326 97398 60562 97634
rect 60646 97398 60882 97634
rect 60326 61718 60562 61954
rect 60646 61718 60882 61954
rect 60326 61398 60562 61634
rect 60646 61398 60882 61634
rect 60326 25718 60562 25954
rect 60646 25718 60882 25954
rect 60326 25398 60562 25634
rect 60646 25398 60882 25634
rect 60326 -5382 60562 -5146
rect 60646 -5382 60882 -5146
rect 60326 -5702 60562 -5466
rect 60646 -5702 60882 -5466
rect 64826 710362 65062 710598
rect 65146 710362 65382 710598
rect 64826 710042 65062 710278
rect 65146 710042 65382 710278
rect 64826 678218 65062 678454
rect 65146 678218 65382 678454
rect 64826 677898 65062 678134
rect 65146 677898 65382 678134
rect 64826 642218 65062 642454
rect 65146 642218 65382 642454
rect 64826 641898 65062 642134
rect 65146 641898 65382 642134
rect 64826 606218 65062 606454
rect 65146 606218 65382 606454
rect 64826 605898 65062 606134
rect 65146 605898 65382 606134
rect 64826 570218 65062 570454
rect 65146 570218 65382 570454
rect 64826 569898 65062 570134
rect 65146 569898 65382 570134
rect 64826 534218 65062 534454
rect 65146 534218 65382 534454
rect 64826 533898 65062 534134
rect 65146 533898 65382 534134
rect 64826 498218 65062 498454
rect 65146 498218 65382 498454
rect 64826 497898 65062 498134
rect 65146 497898 65382 498134
rect 64826 462218 65062 462454
rect 65146 462218 65382 462454
rect 64826 461898 65062 462134
rect 65146 461898 65382 462134
rect 64826 426218 65062 426454
rect 65146 426218 65382 426454
rect 64826 425898 65062 426134
rect 65146 425898 65382 426134
rect 64826 390218 65062 390454
rect 65146 390218 65382 390454
rect 64826 389898 65062 390134
rect 65146 389898 65382 390134
rect 64826 354218 65062 354454
rect 65146 354218 65382 354454
rect 64826 353898 65062 354134
rect 65146 353898 65382 354134
rect 64826 318218 65062 318454
rect 65146 318218 65382 318454
rect 64826 317898 65062 318134
rect 65146 317898 65382 318134
rect 64826 282218 65062 282454
rect 65146 282218 65382 282454
rect 64826 281898 65062 282134
rect 65146 281898 65382 282134
rect 64826 246218 65062 246454
rect 65146 246218 65382 246454
rect 64826 245898 65062 246134
rect 65146 245898 65382 246134
rect 64826 210218 65062 210454
rect 65146 210218 65382 210454
rect 64826 209898 65062 210134
rect 65146 209898 65382 210134
rect 64826 174218 65062 174454
rect 65146 174218 65382 174454
rect 64826 173898 65062 174134
rect 65146 173898 65382 174134
rect 64826 138218 65062 138454
rect 65146 138218 65382 138454
rect 64826 137898 65062 138134
rect 65146 137898 65382 138134
rect 64826 102218 65062 102454
rect 65146 102218 65382 102454
rect 64826 101898 65062 102134
rect 65146 101898 65382 102134
rect 64826 66218 65062 66454
rect 65146 66218 65382 66454
rect 64826 65898 65062 66134
rect 65146 65898 65382 66134
rect 64826 30218 65062 30454
rect 65146 30218 65382 30454
rect 64826 29898 65062 30134
rect 65146 29898 65382 30134
rect 64826 -6342 65062 -6106
rect 65146 -6342 65382 -6106
rect 64826 -6662 65062 -6426
rect 65146 -6662 65382 -6426
rect 69326 711322 69562 711558
rect 69646 711322 69882 711558
rect 69326 711002 69562 711238
rect 69646 711002 69882 711238
rect 69326 682718 69562 682954
rect 69646 682718 69882 682954
rect 69326 682398 69562 682634
rect 69646 682398 69882 682634
rect 69326 646718 69562 646954
rect 69646 646718 69882 646954
rect 69326 646398 69562 646634
rect 69646 646398 69882 646634
rect 69326 610718 69562 610954
rect 69646 610718 69882 610954
rect 69326 610398 69562 610634
rect 69646 610398 69882 610634
rect 69326 574718 69562 574954
rect 69646 574718 69882 574954
rect 69326 574398 69562 574634
rect 69646 574398 69882 574634
rect 69326 538718 69562 538954
rect 69646 538718 69882 538954
rect 69326 538398 69562 538634
rect 69646 538398 69882 538634
rect 69326 502718 69562 502954
rect 69646 502718 69882 502954
rect 69326 502398 69562 502634
rect 69646 502398 69882 502634
rect 69326 466718 69562 466954
rect 69646 466718 69882 466954
rect 69326 466398 69562 466634
rect 69646 466398 69882 466634
rect 69326 430718 69562 430954
rect 69646 430718 69882 430954
rect 69326 430398 69562 430634
rect 69646 430398 69882 430634
rect 69326 394718 69562 394954
rect 69646 394718 69882 394954
rect 69326 394398 69562 394634
rect 69646 394398 69882 394634
rect 69326 358718 69562 358954
rect 69646 358718 69882 358954
rect 69326 358398 69562 358634
rect 69646 358398 69882 358634
rect 69326 322718 69562 322954
rect 69646 322718 69882 322954
rect 69326 322398 69562 322634
rect 69646 322398 69882 322634
rect 69326 286718 69562 286954
rect 69646 286718 69882 286954
rect 69326 286398 69562 286634
rect 69646 286398 69882 286634
rect 69326 250718 69562 250954
rect 69646 250718 69882 250954
rect 69326 250398 69562 250634
rect 69646 250398 69882 250634
rect 69326 214718 69562 214954
rect 69646 214718 69882 214954
rect 69326 214398 69562 214634
rect 69646 214398 69882 214634
rect 69326 178718 69562 178954
rect 69646 178718 69882 178954
rect 69326 178398 69562 178634
rect 69646 178398 69882 178634
rect 69326 142718 69562 142954
rect 69646 142718 69882 142954
rect 69326 142398 69562 142634
rect 69646 142398 69882 142634
rect 69326 106718 69562 106954
rect 69646 106718 69882 106954
rect 69326 106398 69562 106634
rect 69646 106398 69882 106634
rect 69326 70718 69562 70954
rect 69646 70718 69882 70954
rect 69326 70398 69562 70634
rect 69646 70398 69882 70634
rect 69326 34718 69562 34954
rect 69646 34718 69882 34954
rect 69326 34398 69562 34634
rect 69646 34398 69882 34634
rect 69326 -7302 69562 -7066
rect 69646 -7302 69882 -7066
rect 69326 -7622 69562 -7386
rect 69646 -7622 69882 -7386
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 78326 705562 78562 705798
rect 78646 705562 78882 705798
rect 78326 705242 78562 705478
rect 78646 705242 78882 705478
rect 78326 691718 78562 691954
rect 78646 691718 78882 691954
rect 78326 691398 78562 691634
rect 78646 691398 78882 691634
rect 78326 655718 78562 655954
rect 78646 655718 78882 655954
rect 78326 655398 78562 655634
rect 78646 655398 78882 655634
rect 78326 619718 78562 619954
rect 78646 619718 78882 619954
rect 78326 619398 78562 619634
rect 78646 619398 78882 619634
rect 78326 583718 78562 583954
rect 78646 583718 78882 583954
rect 78326 583398 78562 583634
rect 78646 583398 78882 583634
rect 78326 547718 78562 547954
rect 78646 547718 78882 547954
rect 78326 547398 78562 547634
rect 78646 547398 78882 547634
rect 78326 511718 78562 511954
rect 78646 511718 78882 511954
rect 78326 511398 78562 511634
rect 78646 511398 78882 511634
rect 78326 475718 78562 475954
rect 78646 475718 78882 475954
rect 78326 475398 78562 475634
rect 78646 475398 78882 475634
rect 78326 439718 78562 439954
rect 78646 439718 78882 439954
rect 78326 439398 78562 439634
rect 78646 439398 78882 439634
rect 78326 403718 78562 403954
rect 78646 403718 78882 403954
rect 78326 403398 78562 403634
rect 78646 403398 78882 403634
rect 78326 367718 78562 367954
rect 78646 367718 78882 367954
rect 78326 367398 78562 367634
rect 78646 367398 78882 367634
rect 78326 331718 78562 331954
rect 78646 331718 78882 331954
rect 78326 331398 78562 331634
rect 78646 331398 78882 331634
rect 78326 295718 78562 295954
rect 78646 295718 78882 295954
rect 78326 295398 78562 295634
rect 78646 295398 78882 295634
rect 78326 259718 78562 259954
rect 78646 259718 78882 259954
rect 78326 259398 78562 259634
rect 78646 259398 78882 259634
rect 78326 223718 78562 223954
rect 78646 223718 78882 223954
rect 78326 223398 78562 223634
rect 78646 223398 78882 223634
rect 78326 187718 78562 187954
rect 78646 187718 78882 187954
rect 78326 187398 78562 187634
rect 78646 187398 78882 187634
rect 78326 151718 78562 151954
rect 78646 151718 78882 151954
rect 78326 151398 78562 151634
rect 78646 151398 78882 151634
rect 78326 115718 78562 115954
rect 78646 115718 78882 115954
rect 78326 115398 78562 115634
rect 78646 115398 78882 115634
rect 78326 79718 78562 79954
rect 78646 79718 78882 79954
rect 78326 79398 78562 79634
rect 78646 79398 78882 79634
rect 78326 43718 78562 43954
rect 78646 43718 78882 43954
rect 78326 43398 78562 43634
rect 78646 43398 78882 43634
rect 78326 7718 78562 7954
rect 78646 7718 78882 7954
rect 78326 7398 78562 7634
rect 78646 7398 78882 7634
rect 78326 -1542 78562 -1306
rect 78646 -1542 78882 -1306
rect 78326 -1862 78562 -1626
rect 78646 -1862 78882 -1626
rect 82826 706522 83062 706758
rect 83146 706522 83382 706758
rect 82826 706202 83062 706438
rect 83146 706202 83382 706438
rect 82826 696218 83062 696454
rect 83146 696218 83382 696454
rect 82826 695898 83062 696134
rect 83146 695898 83382 696134
rect 82826 660218 83062 660454
rect 83146 660218 83382 660454
rect 82826 659898 83062 660134
rect 83146 659898 83382 660134
rect 82826 624218 83062 624454
rect 83146 624218 83382 624454
rect 82826 623898 83062 624134
rect 83146 623898 83382 624134
rect 82826 588218 83062 588454
rect 83146 588218 83382 588454
rect 82826 587898 83062 588134
rect 83146 587898 83382 588134
rect 82826 552218 83062 552454
rect 83146 552218 83382 552454
rect 82826 551898 83062 552134
rect 83146 551898 83382 552134
rect 82826 516218 83062 516454
rect 83146 516218 83382 516454
rect 82826 515898 83062 516134
rect 83146 515898 83382 516134
rect 82826 480218 83062 480454
rect 83146 480218 83382 480454
rect 82826 479898 83062 480134
rect 83146 479898 83382 480134
rect 82826 444218 83062 444454
rect 83146 444218 83382 444454
rect 82826 443898 83062 444134
rect 83146 443898 83382 444134
rect 82826 408218 83062 408454
rect 83146 408218 83382 408454
rect 82826 407898 83062 408134
rect 83146 407898 83382 408134
rect 82826 372218 83062 372454
rect 83146 372218 83382 372454
rect 82826 371898 83062 372134
rect 83146 371898 83382 372134
rect 82826 336218 83062 336454
rect 83146 336218 83382 336454
rect 82826 335898 83062 336134
rect 83146 335898 83382 336134
rect 82826 300218 83062 300454
rect 83146 300218 83382 300454
rect 82826 299898 83062 300134
rect 83146 299898 83382 300134
rect 82826 264218 83062 264454
rect 83146 264218 83382 264454
rect 82826 263898 83062 264134
rect 83146 263898 83382 264134
rect 82826 228218 83062 228454
rect 83146 228218 83382 228454
rect 82826 227898 83062 228134
rect 83146 227898 83382 228134
rect 82826 192218 83062 192454
rect 83146 192218 83382 192454
rect 82826 191898 83062 192134
rect 83146 191898 83382 192134
rect 82826 156218 83062 156454
rect 83146 156218 83382 156454
rect 82826 155898 83062 156134
rect 83146 155898 83382 156134
rect 82826 120218 83062 120454
rect 83146 120218 83382 120454
rect 82826 119898 83062 120134
rect 83146 119898 83382 120134
rect 82826 84218 83062 84454
rect 83146 84218 83382 84454
rect 82826 83898 83062 84134
rect 83146 83898 83382 84134
rect 82826 48218 83062 48454
rect 83146 48218 83382 48454
rect 82826 47898 83062 48134
rect 83146 47898 83382 48134
rect 82826 12218 83062 12454
rect 83146 12218 83382 12454
rect 82826 11898 83062 12134
rect 83146 11898 83382 12134
rect 82826 -2502 83062 -2266
rect 83146 -2502 83382 -2266
rect 82826 -2822 83062 -2586
rect 83146 -2822 83382 -2586
rect 87326 707482 87562 707718
rect 87646 707482 87882 707718
rect 87326 707162 87562 707398
rect 87646 707162 87882 707398
rect 87326 700718 87562 700954
rect 87646 700718 87882 700954
rect 87326 700398 87562 700634
rect 87646 700398 87882 700634
rect 87326 664718 87562 664954
rect 87646 664718 87882 664954
rect 87326 664398 87562 664634
rect 87646 664398 87882 664634
rect 87326 628718 87562 628954
rect 87646 628718 87882 628954
rect 87326 628398 87562 628634
rect 87646 628398 87882 628634
rect 87326 592718 87562 592954
rect 87646 592718 87882 592954
rect 87326 592398 87562 592634
rect 87646 592398 87882 592634
rect 87326 556718 87562 556954
rect 87646 556718 87882 556954
rect 87326 556398 87562 556634
rect 87646 556398 87882 556634
rect 87326 520718 87562 520954
rect 87646 520718 87882 520954
rect 87326 520398 87562 520634
rect 87646 520398 87882 520634
rect 87326 484718 87562 484954
rect 87646 484718 87882 484954
rect 87326 484398 87562 484634
rect 87646 484398 87882 484634
rect 87326 448718 87562 448954
rect 87646 448718 87882 448954
rect 87326 448398 87562 448634
rect 87646 448398 87882 448634
rect 87326 412718 87562 412954
rect 87646 412718 87882 412954
rect 87326 412398 87562 412634
rect 87646 412398 87882 412634
rect 87326 376718 87562 376954
rect 87646 376718 87882 376954
rect 87326 376398 87562 376634
rect 87646 376398 87882 376634
rect 87326 340718 87562 340954
rect 87646 340718 87882 340954
rect 87326 340398 87562 340634
rect 87646 340398 87882 340634
rect 87326 304718 87562 304954
rect 87646 304718 87882 304954
rect 87326 304398 87562 304634
rect 87646 304398 87882 304634
rect 87326 268718 87562 268954
rect 87646 268718 87882 268954
rect 87326 268398 87562 268634
rect 87646 268398 87882 268634
rect 87326 232718 87562 232954
rect 87646 232718 87882 232954
rect 87326 232398 87562 232634
rect 87646 232398 87882 232634
rect 87326 196718 87562 196954
rect 87646 196718 87882 196954
rect 87326 196398 87562 196634
rect 87646 196398 87882 196634
rect 87326 160718 87562 160954
rect 87646 160718 87882 160954
rect 87326 160398 87562 160634
rect 87646 160398 87882 160634
rect 87326 124718 87562 124954
rect 87646 124718 87882 124954
rect 87326 124398 87562 124634
rect 87646 124398 87882 124634
rect 87326 88718 87562 88954
rect 87646 88718 87882 88954
rect 87326 88398 87562 88634
rect 87646 88398 87882 88634
rect 87326 52718 87562 52954
rect 87646 52718 87882 52954
rect 87326 52398 87562 52634
rect 87646 52398 87882 52634
rect 87326 16718 87562 16954
rect 87646 16718 87882 16954
rect 87326 16398 87562 16634
rect 87646 16398 87882 16634
rect 87326 -3462 87562 -3226
rect 87646 -3462 87882 -3226
rect 87326 -3782 87562 -3546
rect 87646 -3782 87882 -3546
rect 91826 708442 92062 708678
rect 92146 708442 92382 708678
rect 91826 708122 92062 708358
rect 92146 708122 92382 708358
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 91826 129218 92062 129454
rect 92146 129218 92382 129454
rect 91826 128898 92062 129134
rect 92146 128898 92382 129134
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -4422 92062 -4186
rect 92146 -4422 92382 -4186
rect 91826 -4742 92062 -4506
rect 92146 -4742 92382 -4506
rect 96326 709402 96562 709638
rect 96646 709402 96882 709638
rect 96326 709082 96562 709318
rect 96646 709082 96882 709318
rect 96326 673718 96562 673954
rect 96646 673718 96882 673954
rect 96326 673398 96562 673634
rect 96646 673398 96882 673634
rect 96326 637718 96562 637954
rect 96646 637718 96882 637954
rect 96326 637398 96562 637634
rect 96646 637398 96882 637634
rect 96326 601718 96562 601954
rect 96646 601718 96882 601954
rect 96326 601398 96562 601634
rect 96646 601398 96882 601634
rect 96326 565718 96562 565954
rect 96646 565718 96882 565954
rect 96326 565398 96562 565634
rect 96646 565398 96882 565634
rect 96326 529718 96562 529954
rect 96646 529718 96882 529954
rect 96326 529398 96562 529634
rect 96646 529398 96882 529634
rect 96326 493718 96562 493954
rect 96646 493718 96882 493954
rect 96326 493398 96562 493634
rect 96646 493398 96882 493634
rect 96326 457718 96562 457954
rect 96646 457718 96882 457954
rect 96326 457398 96562 457634
rect 96646 457398 96882 457634
rect 96326 421718 96562 421954
rect 96646 421718 96882 421954
rect 96326 421398 96562 421634
rect 96646 421398 96882 421634
rect 96326 385718 96562 385954
rect 96646 385718 96882 385954
rect 96326 385398 96562 385634
rect 96646 385398 96882 385634
rect 96326 349718 96562 349954
rect 96646 349718 96882 349954
rect 96326 349398 96562 349634
rect 96646 349398 96882 349634
rect 96326 313718 96562 313954
rect 96646 313718 96882 313954
rect 96326 313398 96562 313634
rect 96646 313398 96882 313634
rect 96326 277718 96562 277954
rect 96646 277718 96882 277954
rect 96326 277398 96562 277634
rect 96646 277398 96882 277634
rect 96326 241718 96562 241954
rect 96646 241718 96882 241954
rect 96326 241398 96562 241634
rect 96646 241398 96882 241634
rect 96326 205718 96562 205954
rect 96646 205718 96882 205954
rect 96326 205398 96562 205634
rect 96646 205398 96882 205634
rect 96326 169718 96562 169954
rect 96646 169718 96882 169954
rect 96326 169398 96562 169634
rect 96646 169398 96882 169634
rect 96326 133718 96562 133954
rect 96646 133718 96882 133954
rect 96326 133398 96562 133634
rect 96646 133398 96882 133634
rect 96326 97718 96562 97954
rect 96646 97718 96882 97954
rect 96326 97398 96562 97634
rect 96646 97398 96882 97634
rect 96326 61718 96562 61954
rect 96646 61718 96882 61954
rect 96326 61398 96562 61634
rect 96646 61398 96882 61634
rect 96326 25718 96562 25954
rect 96646 25718 96882 25954
rect 96326 25398 96562 25634
rect 96646 25398 96882 25634
rect 96326 -5382 96562 -5146
rect 96646 -5382 96882 -5146
rect 96326 -5702 96562 -5466
rect 96646 -5702 96882 -5466
rect 100826 710362 101062 710598
rect 101146 710362 101382 710598
rect 100826 710042 101062 710278
rect 101146 710042 101382 710278
rect 100826 678218 101062 678454
rect 101146 678218 101382 678454
rect 100826 677898 101062 678134
rect 101146 677898 101382 678134
rect 100826 642218 101062 642454
rect 101146 642218 101382 642454
rect 100826 641898 101062 642134
rect 101146 641898 101382 642134
rect 100826 606218 101062 606454
rect 101146 606218 101382 606454
rect 100826 605898 101062 606134
rect 101146 605898 101382 606134
rect 100826 570218 101062 570454
rect 101146 570218 101382 570454
rect 100826 569898 101062 570134
rect 101146 569898 101382 570134
rect 100826 534218 101062 534454
rect 101146 534218 101382 534454
rect 100826 533898 101062 534134
rect 101146 533898 101382 534134
rect 100826 498218 101062 498454
rect 101146 498218 101382 498454
rect 100826 497898 101062 498134
rect 101146 497898 101382 498134
rect 100826 462218 101062 462454
rect 101146 462218 101382 462454
rect 100826 461898 101062 462134
rect 101146 461898 101382 462134
rect 100826 426218 101062 426454
rect 101146 426218 101382 426454
rect 100826 425898 101062 426134
rect 101146 425898 101382 426134
rect 100826 390218 101062 390454
rect 101146 390218 101382 390454
rect 100826 389898 101062 390134
rect 101146 389898 101382 390134
rect 100826 354218 101062 354454
rect 101146 354218 101382 354454
rect 100826 353898 101062 354134
rect 101146 353898 101382 354134
rect 100826 318218 101062 318454
rect 101146 318218 101382 318454
rect 100826 317898 101062 318134
rect 101146 317898 101382 318134
rect 100826 282218 101062 282454
rect 101146 282218 101382 282454
rect 100826 281898 101062 282134
rect 101146 281898 101382 282134
rect 100826 246218 101062 246454
rect 101146 246218 101382 246454
rect 100826 245898 101062 246134
rect 101146 245898 101382 246134
rect 100826 210218 101062 210454
rect 101146 210218 101382 210454
rect 100826 209898 101062 210134
rect 101146 209898 101382 210134
rect 100826 174218 101062 174454
rect 101146 174218 101382 174454
rect 100826 173898 101062 174134
rect 101146 173898 101382 174134
rect 100826 138218 101062 138454
rect 101146 138218 101382 138454
rect 100826 137898 101062 138134
rect 101146 137898 101382 138134
rect 100826 102218 101062 102454
rect 101146 102218 101382 102454
rect 100826 101898 101062 102134
rect 101146 101898 101382 102134
rect 100826 66218 101062 66454
rect 101146 66218 101382 66454
rect 100826 65898 101062 66134
rect 101146 65898 101382 66134
rect 100826 30218 101062 30454
rect 101146 30218 101382 30454
rect 100826 29898 101062 30134
rect 101146 29898 101382 30134
rect 100826 -6342 101062 -6106
rect 101146 -6342 101382 -6106
rect 100826 -6662 101062 -6426
rect 101146 -6662 101382 -6426
rect 105326 711322 105562 711558
rect 105646 711322 105882 711558
rect 105326 711002 105562 711238
rect 105646 711002 105882 711238
rect 105326 682718 105562 682954
rect 105646 682718 105882 682954
rect 105326 682398 105562 682634
rect 105646 682398 105882 682634
rect 105326 646718 105562 646954
rect 105646 646718 105882 646954
rect 105326 646398 105562 646634
rect 105646 646398 105882 646634
rect 105326 610718 105562 610954
rect 105646 610718 105882 610954
rect 105326 610398 105562 610634
rect 105646 610398 105882 610634
rect 105326 574718 105562 574954
rect 105646 574718 105882 574954
rect 105326 574398 105562 574634
rect 105646 574398 105882 574634
rect 105326 538718 105562 538954
rect 105646 538718 105882 538954
rect 105326 538398 105562 538634
rect 105646 538398 105882 538634
rect 105326 502718 105562 502954
rect 105646 502718 105882 502954
rect 105326 502398 105562 502634
rect 105646 502398 105882 502634
rect 105326 466718 105562 466954
rect 105646 466718 105882 466954
rect 105326 466398 105562 466634
rect 105646 466398 105882 466634
rect 105326 430718 105562 430954
rect 105646 430718 105882 430954
rect 105326 430398 105562 430634
rect 105646 430398 105882 430634
rect 105326 394718 105562 394954
rect 105646 394718 105882 394954
rect 105326 394398 105562 394634
rect 105646 394398 105882 394634
rect 105326 358718 105562 358954
rect 105646 358718 105882 358954
rect 105326 358398 105562 358634
rect 105646 358398 105882 358634
rect 105326 322718 105562 322954
rect 105646 322718 105882 322954
rect 105326 322398 105562 322634
rect 105646 322398 105882 322634
rect 105326 286718 105562 286954
rect 105646 286718 105882 286954
rect 105326 286398 105562 286634
rect 105646 286398 105882 286634
rect 105326 250718 105562 250954
rect 105646 250718 105882 250954
rect 105326 250398 105562 250634
rect 105646 250398 105882 250634
rect 105326 214718 105562 214954
rect 105646 214718 105882 214954
rect 105326 214398 105562 214634
rect 105646 214398 105882 214634
rect 105326 178718 105562 178954
rect 105646 178718 105882 178954
rect 105326 178398 105562 178634
rect 105646 178398 105882 178634
rect 105326 142718 105562 142954
rect 105646 142718 105882 142954
rect 105326 142398 105562 142634
rect 105646 142398 105882 142634
rect 105326 106718 105562 106954
rect 105646 106718 105882 106954
rect 105326 106398 105562 106634
rect 105646 106398 105882 106634
rect 105326 70718 105562 70954
rect 105646 70718 105882 70954
rect 105326 70398 105562 70634
rect 105646 70398 105882 70634
rect 105326 34718 105562 34954
rect 105646 34718 105882 34954
rect 105326 34398 105562 34634
rect 105646 34398 105882 34634
rect 105326 -7302 105562 -7066
rect 105646 -7302 105882 -7066
rect 105326 -7622 105562 -7386
rect 105646 -7622 105882 -7386
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 114326 705562 114562 705798
rect 114646 705562 114882 705798
rect 114326 705242 114562 705478
rect 114646 705242 114882 705478
rect 114326 691718 114562 691954
rect 114646 691718 114882 691954
rect 114326 691398 114562 691634
rect 114646 691398 114882 691634
rect 114326 655718 114562 655954
rect 114646 655718 114882 655954
rect 114326 655398 114562 655634
rect 114646 655398 114882 655634
rect 114326 619718 114562 619954
rect 114646 619718 114882 619954
rect 114326 619398 114562 619634
rect 114646 619398 114882 619634
rect 114326 583718 114562 583954
rect 114646 583718 114882 583954
rect 114326 583398 114562 583634
rect 114646 583398 114882 583634
rect 114326 547718 114562 547954
rect 114646 547718 114882 547954
rect 114326 547398 114562 547634
rect 114646 547398 114882 547634
rect 114326 511718 114562 511954
rect 114646 511718 114882 511954
rect 114326 511398 114562 511634
rect 114646 511398 114882 511634
rect 114326 475718 114562 475954
rect 114646 475718 114882 475954
rect 114326 475398 114562 475634
rect 114646 475398 114882 475634
rect 114326 439718 114562 439954
rect 114646 439718 114882 439954
rect 114326 439398 114562 439634
rect 114646 439398 114882 439634
rect 114326 403718 114562 403954
rect 114646 403718 114882 403954
rect 114326 403398 114562 403634
rect 114646 403398 114882 403634
rect 114326 367718 114562 367954
rect 114646 367718 114882 367954
rect 114326 367398 114562 367634
rect 114646 367398 114882 367634
rect 114326 331718 114562 331954
rect 114646 331718 114882 331954
rect 114326 331398 114562 331634
rect 114646 331398 114882 331634
rect 114326 295718 114562 295954
rect 114646 295718 114882 295954
rect 114326 295398 114562 295634
rect 114646 295398 114882 295634
rect 114326 259718 114562 259954
rect 114646 259718 114882 259954
rect 114326 259398 114562 259634
rect 114646 259398 114882 259634
rect 114326 223718 114562 223954
rect 114646 223718 114882 223954
rect 114326 223398 114562 223634
rect 114646 223398 114882 223634
rect 114326 187718 114562 187954
rect 114646 187718 114882 187954
rect 114326 187398 114562 187634
rect 114646 187398 114882 187634
rect 114326 151718 114562 151954
rect 114646 151718 114882 151954
rect 114326 151398 114562 151634
rect 114646 151398 114882 151634
rect 118826 706522 119062 706758
rect 119146 706522 119382 706758
rect 118826 706202 119062 706438
rect 119146 706202 119382 706438
rect 118826 696218 119062 696454
rect 119146 696218 119382 696454
rect 118826 695898 119062 696134
rect 119146 695898 119382 696134
rect 118826 660218 119062 660454
rect 119146 660218 119382 660454
rect 118826 659898 119062 660134
rect 119146 659898 119382 660134
rect 118826 624218 119062 624454
rect 119146 624218 119382 624454
rect 118826 623898 119062 624134
rect 119146 623898 119382 624134
rect 118826 588218 119062 588454
rect 119146 588218 119382 588454
rect 118826 587898 119062 588134
rect 119146 587898 119382 588134
rect 118826 552218 119062 552454
rect 119146 552218 119382 552454
rect 118826 551898 119062 552134
rect 119146 551898 119382 552134
rect 118826 516218 119062 516454
rect 119146 516218 119382 516454
rect 118826 515898 119062 516134
rect 119146 515898 119382 516134
rect 118826 480218 119062 480454
rect 119146 480218 119382 480454
rect 118826 479898 119062 480134
rect 119146 479898 119382 480134
rect 118826 444218 119062 444454
rect 119146 444218 119382 444454
rect 118826 443898 119062 444134
rect 119146 443898 119382 444134
rect 118826 408218 119062 408454
rect 119146 408218 119382 408454
rect 118826 407898 119062 408134
rect 119146 407898 119382 408134
rect 118826 372218 119062 372454
rect 119146 372218 119382 372454
rect 118826 371898 119062 372134
rect 119146 371898 119382 372134
rect 118826 336218 119062 336454
rect 119146 336218 119382 336454
rect 118826 335898 119062 336134
rect 119146 335898 119382 336134
rect 118826 300218 119062 300454
rect 119146 300218 119382 300454
rect 118826 299898 119062 300134
rect 119146 299898 119382 300134
rect 118826 264218 119062 264454
rect 119146 264218 119382 264454
rect 118826 263898 119062 264134
rect 119146 263898 119382 264134
rect 118826 228218 119062 228454
rect 119146 228218 119382 228454
rect 118826 227898 119062 228134
rect 119146 227898 119382 228134
rect 118826 192218 119062 192454
rect 119146 192218 119382 192454
rect 118826 191898 119062 192134
rect 119146 191898 119382 192134
rect 118826 156218 119062 156454
rect 119146 156218 119382 156454
rect 118826 155898 119062 156134
rect 119146 155898 119382 156134
rect 123326 707482 123562 707718
rect 123646 707482 123882 707718
rect 123326 707162 123562 707398
rect 123646 707162 123882 707398
rect 123326 700718 123562 700954
rect 123646 700718 123882 700954
rect 123326 700398 123562 700634
rect 123646 700398 123882 700634
rect 123326 664718 123562 664954
rect 123646 664718 123882 664954
rect 123326 664398 123562 664634
rect 123646 664398 123882 664634
rect 123326 628718 123562 628954
rect 123646 628718 123882 628954
rect 123326 628398 123562 628634
rect 123646 628398 123882 628634
rect 123326 592718 123562 592954
rect 123646 592718 123882 592954
rect 123326 592398 123562 592634
rect 123646 592398 123882 592634
rect 123326 556718 123562 556954
rect 123646 556718 123882 556954
rect 123326 556398 123562 556634
rect 123646 556398 123882 556634
rect 123326 520718 123562 520954
rect 123646 520718 123882 520954
rect 123326 520398 123562 520634
rect 123646 520398 123882 520634
rect 123326 484718 123562 484954
rect 123646 484718 123882 484954
rect 123326 484398 123562 484634
rect 123646 484398 123882 484634
rect 123326 448718 123562 448954
rect 123646 448718 123882 448954
rect 123326 448398 123562 448634
rect 123646 448398 123882 448634
rect 123326 412718 123562 412954
rect 123646 412718 123882 412954
rect 123326 412398 123562 412634
rect 123646 412398 123882 412634
rect 123326 376718 123562 376954
rect 123646 376718 123882 376954
rect 123326 376398 123562 376634
rect 123646 376398 123882 376634
rect 123326 340718 123562 340954
rect 123646 340718 123882 340954
rect 123326 340398 123562 340634
rect 123646 340398 123882 340634
rect 123326 304718 123562 304954
rect 123646 304718 123882 304954
rect 123326 304398 123562 304634
rect 123646 304398 123882 304634
rect 123326 268718 123562 268954
rect 123646 268718 123882 268954
rect 123326 268398 123562 268634
rect 123646 268398 123882 268634
rect 123326 232718 123562 232954
rect 123646 232718 123882 232954
rect 123326 232398 123562 232634
rect 123646 232398 123882 232634
rect 123326 196718 123562 196954
rect 123646 196718 123882 196954
rect 123326 196398 123562 196634
rect 123646 196398 123882 196634
rect 123326 160718 123562 160954
rect 123646 160718 123882 160954
rect 123326 160398 123562 160634
rect 123646 160398 123882 160634
rect 127826 708442 128062 708678
rect 128146 708442 128382 708678
rect 127826 708122 128062 708358
rect 128146 708122 128382 708358
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 127826 165218 128062 165454
rect 128146 165218 128382 165454
rect 127826 164898 128062 165134
rect 128146 164898 128382 165134
rect 132326 709402 132562 709638
rect 132646 709402 132882 709638
rect 132326 709082 132562 709318
rect 132646 709082 132882 709318
rect 132326 673718 132562 673954
rect 132646 673718 132882 673954
rect 132326 673398 132562 673634
rect 132646 673398 132882 673634
rect 132326 637718 132562 637954
rect 132646 637718 132882 637954
rect 132326 637398 132562 637634
rect 132646 637398 132882 637634
rect 132326 601718 132562 601954
rect 132646 601718 132882 601954
rect 132326 601398 132562 601634
rect 132646 601398 132882 601634
rect 132326 565718 132562 565954
rect 132646 565718 132882 565954
rect 132326 565398 132562 565634
rect 132646 565398 132882 565634
rect 132326 529718 132562 529954
rect 132646 529718 132882 529954
rect 132326 529398 132562 529634
rect 132646 529398 132882 529634
rect 132326 493718 132562 493954
rect 132646 493718 132882 493954
rect 132326 493398 132562 493634
rect 132646 493398 132882 493634
rect 132326 457718 132562 457954
rect 132646 457718 132882 457954
rect 132326 457398 132562 457634
rect 132646 457398 132882 457634
rect 132326 421718 132562 421954
rect 132646 421718 132882 421954
rect 132326 421398 132562 421634
rect 132646 421398 132882 421634
rect 132326 385718 132562 385954
rect 132646 385718 132882 385954
rect 132326 385398 132562 385634
rect 132646 385398 132882 385634
rect 132326 349718 132562 349954
rect 132646 349718 132882 349954
rect 132326 349398 132562 349634
rect 132646 349398 132882 349634
rect 132326 313718 132562 313954
rect 132646 313718 132882 313954
rect 132326 313398 132562 313634
rect 132646 313398 132882 313634
rect 132326 277718 132562 277954
rect 132646 277718 132882 277954
rect 132326 277398 132562 277634
rect 132646 277398 132882 277634
rect 132326 241718 132562 241954
rect 132646 241718 132882 241954
rect 132326 241398 132562 241634
rect 132646 241398 132882 241634
rect 132326 205718 132562 205954
rect 132646 205718 132882 205954
rect 132326 205398 132562 205634
rect 132646 205398 132882 205634
rect 132326 169718 132562 169954
rect 132646 169718 132882 169954
rect 132326 169398 132562 169634
rect 132646 169398 132882 169634
rect 136826 710362 137062 710598
rect 137146 710362 137382 710598
rect 136826 710042 137062 710278
rect 137146 710042 137382 710278
rect 136826 678218 137062 678454
rect 137146 678218 137382 678454
rect 136826 677898 137062 678134
rect 137146 677898 137382 678134
rect 136826 642218 137062 642454
rect 137146 642218 137382 642454
rect 136826 641898 137062 642134
rect 137146 641898 137382 642134
rect 136826 606218 137062 606454
rect 137146 606218 137382 606454
rect 136826 605898 137062 606134
rect 137146 605898 137382 606134
rect 136826 570218 137062 570454
rect 137146 570218 137382 570454
rect 136826 569898 137062 570134
rect 137146 569898 137382 570134
rect 136826 534218 137062 534454
rect 137146 534218 137382 534454
rect 136826 533898 137062 534134
rect 137146 533898 137382 534134
rect 136826 498218 137062 498454
rect 137146 498218 137382 498454
rect 136826 497898 137062 498134
rect 137146 497898 137382 498134
rect 136826 462218 137062 462454
rect 137146 462218 137382 462454
rect 136826 461898 137062 462134
rect 137146 461898 137382 462134
rect 136826 426218 137062 426454
rect 137146 426218 137382 426454
rect 136826 425898 137062 426134
rect 137146 425898 137382 426134
rect 136826 390218 137062 390454
rect 137146 390218 137382 390454
rect 136826 389898 137062 390134
rect 137146 389898 137382 390134
rect 136826 354218 137062 354454
rect 137146 354218 137382 354454
rect 136826 353898 137062 354134
rect 137146 353898 137382 354134
rect 136826 318218 137062 318454
rect 137146 318218 137382 318454
rect 136826 317898 137062 318134
rect 137146 317898 137382 318134
rect 136826 282218 137062 282454
rect 137146 282218 137382 282454
rect 136826 281898 137062 282134
rect 137146 281898 137382 282134
rect 136826 246218 137062 246454
rect 137146 246218 137382 246454
rect 136826 245898 137062 246134
rect 137146 245898 137382 246134
rect 136826 210218 137062 210454
rect 137146 210218 137382 210454
rect 136826 209898 137062 210134
rect 137146 209898 137382 210134
rect 136826 174218 137062 174454
rect 137146 174218 137382 174454
rect 136826 173898 137062 174134
rect 137146 173898 137382 174134
rect 141326 711322 141562 711558
rect 141646 711322 141882 711558
rect 141326 711002 141562 711238
rect 141646 711002 141882 711238
rect 141326 682718 141562 682954
rect 141646 682718 141882 682954
rect 141326 682398 141562 682634
rect 141646 682398 141882 682634
rect 141326 646718 141562 646954
rect 141646 646718 141882 646954
rect 141326 646398 141562 646634
rect 141646 646398 141882 646634
rect 141326 610718 141562 610954
rect 141646 610718 141882 610954
rect 141326 610398 141562 610634
rect 141646 610398 141882 610634
rect 141326 574718 141562 574954
rect 141646 574718 141882 574954
rect 141326 574398 141562 574634
rect 141646 574398 141882 574634
rect 141326 538718 141562 538954
rect 141646 538718 141882 538954
rect 141326 538398 141562 538634
rect 141646 538398 141882 538634
rect 141326 502718 141562 502954
rect 141646 502718 141882 502954
rect 141326 502398 141562 502634
rect 141646 502398 141882 502634
rect 141326 466718 141562 466954
rect 141646 466718 141882 466954
rect 141326 466398 141562 466634
rect 141646 466398 141882 466634
rect 141326 430718 141562 430954
rect 141646 430718 141882 430954
rect 141326 430398 141562 430634
rect 141646 430398 141882 430634
rect 141326 394718 141562 394954
rect 141646 394718 141882 394954
rect 141326 394398 141562 394634
rect 141646 394398 141882 394634
rect 141326 358718 141562 358954
rect 141646 358718 141882 358954
rect 141326 358398 141562 358634
rect 141646 358398 141882 358634
rect 141326 322718 141562 322954
rect 141646 322718 141882 322954
rect 141326 322398 141562 322634
rect 141646 322398 141882 322634
rect 141326 286718 141562 286954
rect 141646 286718 141882 286954
rect 141326 286398 141562 286634
rect 141646 286398 141882 286634
rect 141326 250718 141562 250954
rect 141646 250718 141882 250954
rect 141326 250398 141562 250634
rect 141646 250398 141882 250634
rect 141326 214718 141562 214954
rect 141646 214718 141882 214954
rect 141326 214398 141562 214634
rect 141646 214398 141882 214634
rect 141326 178718 141562 178954
rect 141646 178718 141882 178954
rect 141326 178398 141562 178634
rect 141646 178398 141882 178634
rect 141326 142718 141562 142954
rect 141646 142718 141882 142954
rect 141326 142398 141562 142634
rect 141646 142398 141882 142634
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 150326 705562 150562 705798
rect 150646 705562 150882 705798
rect 150326 705242 150562 705478
rect 150646 705242 150882 705478
rect 150326 691718 150562 691954
rect 150646 691718 150882 691954
rect 150326 691398 150562 691634
rect 150646 691398 150882 691634
rect 150326 655718 150562 655954
rect 150646 655718 150882 655954
rect 150326 655398 150562 655634
rect 150646 655398 150882 655634
rect 150326 619718 150562 619954
rect 150646 619718 150882 619954
rect 150326 619398 150562 619634
rect 150646 619398 150882 619634
rect 150326 583718 150562 583954
rect 150646 583718 150882 583954
rect 150326 583398 150562 583634
rect 150646 583398 150882 583634
rect 150326 547718 150562 547954
rect 150646 547718 150882 547954
rect 150326 547398 150562 547634
rect 150646 547398 150882 547634
rect 150326 511718 150562 511954
rect 150646 511718 150882 511954
rect 150326 511398 150562 511634
rect 150646 511398 150882 511634
rect 150326 475718 150562 475954
rect 150646 475718 150882 475954
rect 150326 475398 150562 475634
rect 150646 475398 150882 475634
rect 150326 439718 150562 439954
rect 150646 439718 150882 439954
rect 150326 439398 150562 439634
rect 150646 439398 150882 439634
rect 150326 403718 150562 403954
rect 150646 403718 150882 403954
rect 150326 403398 150562 403634
rect 150646 403398 150882 403634
rect 150326 367718 150562 367954
rect 150646 367718 150882 367954
rect 150326 367398 150562 367634
rect 150646 367398 150882 367634
rect 150326 331718 150562 331954
rect 150646 331718 150882 331954
rect 150326 331398 150562 331634
rect 150646 331398 150882 331634
rect 150326 295718 150562 295954
rect 150646 295718 150882 295954
rect 150326 295398 150562 295634
rect 150646 295398 150882 295634
rect 150326 259718 150562 259954
rect 150646 259718 150882 259954
rect 150326 259398 150562 259634
rect 150646 259398 150882 259634
rect 150326 223718 150562 223954
rect 150646 223718 150882 223954
rect 150326 223398 150562 223634
rect 150646 223398 150882 223634
rect 150326 187718 150562 187954
rect 150646 187718 150882 187954
rect 150326 187398 150562 187634
rect 150646 187398 150882 187634
rect 150326 151718 150562 151954
rect 150646 151718 150882 151954
rect 150326 151398 150562 151634
rect 150646 151398 150882 151634
rect 154826 706522 155062 706758
rect 155146 706522 155382 706758
rect 154826 706202 155062 706438
rect 155146 706202 155382 706438
rect 154826 696218 155062 696454
rect 155146 696218 155382 696454
rect 154826 695898 155062 696134
rect 155146 695898 155382 696134
rect 154826 660218 155062 660454
rect 155146 660218 155382 660454
rect 154826 659898 155062 660134
rect 155146 659898 155382 660134
rect 154826 624218 155062 624454
rect 155146 624218 155382 624454
rect 154826 623898 155062 624134
rect 155146 623898 155382 624134
rect 154826 588218 155062 588454
rect 155146 588218 155382 588454
rect 154826 587898 155062 588134
rect 155146 587898 155382 588134
rect 154826 552218 155062 552454
rect 155146 552218 155382 552454
rect 154826 551898 155062 552134
rect 155146 551898 155382 552134
rect 154826 516218 155062 516454
rect 155146 516218 155382 516454
rect 154826 515898 155062 516134
rect 155146 515898 155382 516134
rect 154826 480218 155062 480454
rect 155146 480218 155382 480454
rect 154826 479898 155062 480134
rect 155146 479898 155382 480134
rect 154826 444218 155062 444454
rect 155146 444218 155382 444454
rect 154826 443898 155062 444134
rect 155146 443898 155382 444134
rect 154826 408218 155062 408454
rect 155146 408218 155382 408454
rect 154826 407898 155062 408134
rect 155146 407898 155382 408134
rect 154826 372218 155062 372454
rect 155146 372218 155382 372454
rect 154826 371898 155062 372134
rect 155146 371898 155382 372134
rect 154826 336218 155062 336454
rect 155146 336218 155382 336454
rect 154826 335898 155062 336134
rect 155146 335898 155382 336134
rect 154826 300218 155062 300454
rect 155146 300218 155382 300454
rect 154826 299898 155062 300134
rect 155146 299898 155382 300134
rect 154826 264218 155062 264454
rect 155146 264218 155382 264454
rect 154826 263898 155062 264134
rect 155146 263898 155382 264134
rect 154826 228218 155062 228454
rect 155146 228218 155382 228454
rect 154826 227898 155062 228134
rect 155146 227898 155382 228134
rect 154826 192218 155062 192454
rect 155146 192218 155382 192454
rect 154826 191898 155062 192134
rect 155146 191898 155382 192134
rect 154826 156218 155062 156454
rect 155146 156218 155382 156454
rect 154826 155898 155062 156134
rect 155146 155898 155382 156134
rect 159326 707482 159562 707718
rect 159646 707482 159882 707718
rect 159326 707162 159562 707398
rect 159646 707162 159882 707398
rect 159326 700718 159562 700954
rect 159646 700718 159882 700954
rect 159326 700398 159562 700634
rect 159646 700398 159882 700634
rect 159326 664718 159562 664954
rect 159646 664718 159882 664954
rect 159326 664398 159562 664634
rect 159646 664398 159882 664634
rect 159326 628718 159562 628954
rect 159646 628718 159882 628954
rect 159326 628398 159562 628634
rect 159646 628398 159882 628634
rect 159326 592718 159562 592954
rect 159646 592718 159882 592954
rect 159326 592398 159562 592634
rect 159646 592398 159882 592634
rect 159326 556718 159562 556954
rect 159646 556718 159882 556954
rect 159326 556398 159562 556634
rect 159646 556398 159882 556634
rect 159326 520718 159562 520954
rect 159646 520718 159882 520954
rect 159326 520398 159562 520634
rect 159646 520398 159882 520634
rect 159326 484718 159562 484954
rect 159646 484718 159882 484954
rect 159326 484398 159562 484634
rect 159646 484398 159882 484634
rect 159326 448718 159562 448954
rect 159646 448718 159882 448954
rect 159326 448398 159562 448634
rect 159646 448398 159882 448634
rect 159326 412718 159562 412954
rect 159646 412718 159882 412954
rect 159326 412398 159562 412634
rect 159646 412398 159882 412634
rect 159326 376718 159562 376954
rect 159646 376718 159882 376954
rect 159326 376398 159562 376634
rect 159646 376398 159882 376634
rect 159326 340718 159562 340954
rect 159646 340718 159882 340954
rect 159326 340398 159562 340634
rect 159646 340398 159882 340634
rect 159326 304718 159562 304954
rect 159646 304718 159882 304954
rect 159326 304398 159562 304634
rect 159646 304398 159882 304634
rect 159326 268718 159562 268954
rect 159646 268718 159882 268954
rect 159326 268398 159562 268634
rect 159646 268398 159882 268634
rect 159326 232718 159562 232954
rect 159646 232718 159882 232954
rect 159326 232398 159562 232634
rect 159646 232398 159882 232634
rect 159326 196718 159562 196954
rect 159646 196718 159882 196954
rect 159326 196398 159562 196634
rect 159646 196398 159882 196634
rect 159326 160718 159562 160954
rect 159646 160718 159882 160954
rect 159326 160398 159562 160634
rect 159646 160398 159882 160634
rect 163826 708442 164062 708678
rect 164146 708442 164382 708678
rect 163826 708122 164062 708358
rect 164146 708122 164382 708358
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 163826 165218 164062 165454
rect 164146 165218 164382 165454
rect 163826 164898 164062 165134
rect 164146 164898 164382 165134
rect 168326 709402 168562 709638
rect 168646 709402 168882 709638
rect 168326 709082 168562 709318
rect 168646 709082 168882 709318
rect 168326 673718 168562 673954
rect 168646 673718 168882 673954
rect 168326 673398 168562 673634
rect 168646 673398 168882 673634
rect 168326 637718 168562 637954
rect 168646 637718 168882 637954
rect 168326 637398 168562 637634
rect 168646 637398 168882 637634
rect 168326 601718 168562 601954
rect 168646 601718 168882 601954
rect 168326 601398 168562 601634
rect 168646 601398 168882 601634
rect 168326 565718 168562 565954
rect 168646 565718 168882 565954
rect 168326 565398 168562 565634
rect 168646 565398 168882 565634
rect 168326 529718 168562 529954
rect 168646 529718 168882 529954
rect 168326 529398 168562 529634
rect 168646 529398 168882 529634
rect 168326 493718 168562 493954
rect 168646 493718 168882 493954
rect 168326 493398 168562 493634
rect 168646 493398 168882 493634
rect 168326 457718 168562 457954
rect 168646 457718 168882 457954
rect 168326 457398 168562 457634
rect 168646 457398 168882 457634
rect 168326 421718 168562 421954
rect 168646 421718 168882 421954
rect 168326 421398 168562 421634
rect 168646 421398 168882 421634
rect 168326 385718 168562 385954
rect 168646 385718 168882 385954
rect 168326 385398 168562 385634
rect 168646 385398 168882 385634
rect 168326 349718 168562 349954
rect 168646 349718 168882 349954
rect 168326 349398 168562 349634
rect 168646 349398 168882 349634
rect 168326 313718 168562 313954
rect 168646 313718 168882 313954
rect 168326 313398 168562 313634
rect 168646 313398 168882 313634
rect 168326 277718 168562 277954
rect 168646 277718 168882 277954
rect 168326 277398 168562 277634
rect 168646 277398 168882 277634
rect 168326 241718 168562 241954
rect 168646 241718 168882 241954
rect 168326 241398 168562 241634
rect 168646 241398 168882 241634
rect 168326 205718 168562 205954
rect 168646 205718 168882 205954
rect 168326 205398 168562 205634
rect 168646 205398 168882 205634
rect 168326 169718 168562 169954
rect 168646 169718 168882 169954
rect 168326 169398 168562 169634
rect 168646 169398 168882 169634
rect 172826 710362 173062 710598
rect 173146 710362 173382 710598
rect 172826 710042 173062 710278
rect 173146 710042 173382 710278
rect 172826 678218 173062 678454
rect 173146 678218 173382 678454
rect 172826 677898 173062 678134
rect 173146 677898 173382 678134
rect 172826 642218 173062 642454
rect 173146 642218 173382 642454
rect 172826 641898 173062 642134
rect 173146 641898 173382 642134
rect 172826 606218 173062 606454
rect 173146 606218 173382 606454
rect 172826 605898 173062 606134
rect 173146 605898 173382 606134
rect 172826 570218 173062 570454
rect 173146 570218 173382 570454
rect 172826 569898 173062 570134
rect 173146 569898 173382 570134
rect 172826 534218 173062 534454
rect 173146 534218 173382 534454
rect 172826 533898 173062 534134
rect 173146 533898 173382 534134
rect 172826 498218 173062 498454
rect 173146 498218 173382 498454
rect 172826 497898 173062 498134
rect 173146 497898 173382 498134
rect 172826 462218 173062 462454
rect 173146 462218 173382 462454
rect 172826 461898 173062 462134
rect 173146 461898 173382 462134
rect 172826 426218 173062 426454
rect 173146 426218 173382 426454
rect 172826 425898 173062 426134
rect 173146 425898 173382 426134
rect 172826 390218 173062 390454
rect 173146 390218 173382 390454
rect 172826 389898 173062 390134
rect 173146 389898 173382 390134
rect 172826 354218 173062 354454
rect 173146 354218 173382 354454
rect 172826 353898 173062 354134
rect 173146 353898 173382 354134
rect 172826 318218 173062 318454
rect 173146 318218 173382 318454
rect 172826 317898 173062 318134
rect 173146 317898 173382 318134
rect 172826 282218 173062 282454
rect 173146 282218 173382 282454
rect 172826 281898 173062 282134
rect 173146 281898 173382 282134
rect 172826 246218 173062 246454
rect 173146 246218 173382 246454
rect 172826 245898 173062 246134
rect 173146 245898 173382 246134
rect 172826 210218 173062 210454
rect 173146 210218 173382 210454
rect 172826 209898 173062 210134
rect 173146 209898 173382 210134
rect 172826 174218 173062 174454
rect 173146 174218 173382 174454
rect 172826 173898 173062 174134
rect 173146 173898 173382 174134
rect 177326 711322 177562 711558
rect 177646 711322 177882 711558
rect 177326 711002 177562 711238
rect 177646 711002 177882 711238
rect 177326 682718 177562 682954
rect 177646 682718 177882 682954
rect 177326 682398 177562 682634
rect 177646 682398 177882 682634
rect 177326 646718 177562 646954
rect 177646 646718 177882 646954
rect 177326 646398 177562 646634
rect 177646 646398 177882 646634
rect 177326 610718 177562 610954
rect 177646 610718 177882 610954
rect 177326 610398 177562 610634
rect 177646 610398 177882 610634
rect 177326 574718 177562 574954
rect 177646 574718 177882 574954
rect 177326 574398 177562 574634
rect 177646 574398 177882 574634
rect 177326 538718 177562 538954
rect 177646 538718 177882 538954
rect 177326 538398 177562 538634
rect 177646 538398 177882 538634
rect 177326 502718 177562 502954
rect 177646 502718 177882 502954
rect 177326 502398 177562 502634
rect 177646 502398 177882 502634
rect 177326 466718 177562 466954
rect 177646 466718 177882 466954
rect 177326 466398 177562 466634
rect 177646 466398 177882 466634
rect 177326 430718 177562 430954
rect 177646 430718 177882 430954
rect 177326 430398 177562 430634
rect 177646 430398 177882 430634
rect 177326 394718 177562 394954
rect 177646 394718 177882 394954
rect 177326 394398 177562 394634
rect 177646 394398 177882 394634
rect 177326 358718 177562 358954
rect 177646 358718 177882 358954
rect 177326 358398 177562 358634
rect 177646 358398 177882 358634
rect 177326 322718 177562 322954
rect 177646 322718 177882 322954
rect 177326 322398 177562 322634
rect 177646 322398 177882 322634
rect 177326 286718 177562 286954
rect 177646 286718 177882 286954
rect 177326 286398 177562 286634
rect 177646 286398 177882 286634
rect 177326 250718 177562 250954
rect 177646 250718 177882 250954
rect 177326 250398 177562 250634
rect 177646 250398 177882 250634
rect 177326 214718 177562 214954
rect 177646 214718 177882 214954
rect 177326 214398 177562 214634
rect 177646 214398 177882 214634
rect 177326 178718 177562 178954
rect 177646 178718 177882 178954
rect 177326 178398 177562 178634
rect 177646 178398 177882 178634
rect 177326 142718 177562 142954
rect 177646 142718 177882 142954
rect 177326 142398 177562 142634
rect 177646 142398 177882 142634
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 186326 705562 186562 705798
rect 186646 705562 186882 705798
rect 186326 705242 186562 705478
rect 186646 705242 186882 705478
rect 186326 691718 186562 691954
rect 186646 691718 186882 691954
rect 186326 691398 186562 691634
rect 186646 691398 186882 691634
rect 186326 655718 186562 655954
rect 186646 655718 186882 655954
rect 186326 655398 186562 655634
rect 186646 655398 186882 655634
rect 186326 619718 186562 619954
rect 186646 619718 186882 619954
rect 186326 619398 186562 619634
rect 186646 619398 186882 619634
rect 186326 583718 186562 583954
rect 186646 583718 186882 583954
rect 186326 583398 186562 583634
rect 186646 583398 186882 583634
rect 186326 547718 186562 547954
rect 186646 547718 186882 547954
rect 186326 547398 186562 547634
rect 186646 547398 186882 547634
rect 186326 511718 186562 511954
rect 186646 511718 186882 511954
rect 186326 511398 186562 511634
rect 186646 511398 186882 511634
rect 186326 475718 186562 475954
rect 186646 475718 186882 475954
rect 186326 475398 186562 475634
rect 186646 475398 186882 475634
rect 186326 439718 186562 439954
rect 186646 439718 186882 439954
rect 186326 439398 186562 439634
rect 186646 439398 186882 439634
rect 186326 403718 186562 403954
rect 186646 403718 186882 403954
rect 186326 403398 186562 403634
rect 186646 403398 186882 403634
rect 186326 367718 186562 367954
rect 186646 367718 186882 367954
rect 186326 367398 186562 367634
rect 186646 367398 186882 367634
rect 186326 331718 186562 331954
rect 186646 331718 186882 331954
rect 186326 331398 186562 331634
rect 186646 331398 186882 331634
rect 186326 295718 186562 295954
rect 186646 295718 186882 295954
rect 186326 295398 186562 295634
rect 186646 295398 186882 295634
rect 186326 259718 186562 259954
rect 186646 259718 186882 259954
rect 186326 259398 186562 259634
rect 186646 259398 186882 259634
rect 186326 223718 186562 223954
rect 186646 223718 186882 223954
rect 186326 223398 186562 223634
rect 186646 223398 186882 223634
rect 186326 187718 186562 187954
rect 186646 187718 186882 187954
rect 186326 187398 186562 187634
rect 186646 187398 186882 187634
rect 186326 151718 186562 151954
rect 186646 151718 186882 151954
rect 186326 151398 186562 151634
rect 186646 151398 186882 151634
rect 190826 706522 191062 706758
rect 191146 706522 191382 706758
rect 190826 706202 191062 706438
rect 191146 706202 191382 706438
rect 190826 696218 191062 696454
rect 191146 696218 191382 696454
rect 190826 695898 191062 696134
rect 191146 695898 191382 696134
rect 190826 660218 191062 660454
rect 191146 660218 191382 660454
rect 190826 659898 191062 660134
rect 191146 659898 191382 660134
rect 190826 624218 191062 624454
rect 191146 624218 191382 624454
rect 190826 623898 191062 624134
rect 191146 623898 191382 624134
rect 190826 588218 191062 588454
rect 191146 588218 191382 588454
rect 190826 587898 191062 588134
rect 191146 587898 191382 588134
rect 190826 552218 191062 552454
rect 191146 552218 191382 552454
rect 190826 551898 191062 552134
rect 191146 551898 191382 552134
rect 190826 516218 191062 516454
rect 191146 516218 191382 516454
rect 190826 515898 191062 516134
rect 191146 515898 191382 516134
rect 190826 480218 191062 480454
rect 191146 480218 191382 480454
rect 190826 479898 191062 480134
rect 191146 479898 191382 480134
rect 190826 444218 191062 444454
rect 191146 444218 191382 444454
rect 190826 443898 191062 444134
rect 191146 443898 191382 444134
rect 190826 408218 191062 408454
rect 191146 408218 191382 408454
rect 190826 407898 191062 408134
rect 191146 407898 191382 408134
rect 190826 372218 191062 372454
rect 191146 372218 191382 372454
rect 190826 371898 191062 372134
rect 191146 371898 191382 372134
rect 190826 336218 191062 336454
rect 191146 336218 191382 336454
rect 190826 335898 191062 336134
rect 191146 335898 191382 336134
rect 190826 300218 191062 300454
rect 191146 300218 191382 300454
rect 190826 299898 191062 300134
rect 191146 299898 191382 300134
rect 190826 264218 191062 264454
rect 191146 264218 191382 264454
rect 190826 263898 191062 264134
rect 191146 263898 191382 264134
rect 190826 228218 191062 228454
rect 191146 228218 191382 228454
rect 190826 227898 191062 228134
rect 191146 227898 191382 228134
rect 190826 192218 191062 192454
rect 191146 192218 191382 192454
rect 190826 191898 191062 192134
rect 191146 191898 191382 192134
rect 190826 156218 191062 156454
rect 191146 156218 191382 156454
rect 190826 155898 191062 156134
rect 191146 155898 191382 156134
rect 195326 707482 195562 707718
rect 195646 707482 195882 707718
rect 195326 707162 195562 707398
rect 195646 707162 195882 707398
rect 195326 700718 195562 700954
rect 195646 700718 195882 700954
rect 195326 700398 195562 700634
rect 195646 700398 195882 700634
rect 195326 664718 195562 664954
rect 195646 664718 195882 664954
rect 195326 664398 195562 664634
rect 195646 664398 195882 664634
rect 195326 628718 195562 628954
rect 195646 628718 195882 628954
rect 195326 628398 195562 628634
rect 195646 628398 195882 628634
rect 195326 592718 195562 592954
rect 195646 592718 195882 592954
rect 195326 592398 195562 592634
rect 195646 592398 195882 592634
rect 195326 556718 195562 556954
rect 195646 556718 195882 556954
rect 195326 556398 195562 556634
rect 195646 556398 195882 556634
rect 195326 520718 195562 520954
rect 195646 520718 195882 520954
rect 195326 520398 195562 520634
rect 195646 520398 195882 520634
rect 195326 484718 195562 484954
rect 195646 484718 195882 484954
rect 195326 484398 195562 484634
rect 195646 484398 195882 484634
rect 195326 448718 195562 448954
rect 195646 448718 195882 448954
rect 195326 448398 195562 448634
rect 195646 448398 195882 448634
rect 195326 412718 195562 412954
rect 195646 412718 195882 412954
rect 195326 412398 195562 412634
rect 195646 412398 195882 412634
rect 195326 376718 195562 376954
rect 195646 376718 195882 376954
rect 195326 376398 195562 376634
rect 195646 376398 195882 376634
rect 195326 340718 195562 340954
rect 195646 340718 195882 340954
rect 195326 340398 195562 340634
rect 195646 340398 195882 340634
rect 195326 304718 195562 304954
rect 195646 304718 195882 304954
rect 195326 304398 195562 304634
rect 195646 304398 195882 304634
rect 195326 268718 195562 268954
rect 195646 268718 195882 268954
rect 195326 268398 195562 268634
rect 195646 268398 195882 268634
rect 195326 232718 195562 232954
rect 195646 232718 195882 232954
rect 195326 232398 195562 232634
rect 195646 232398 195882 232634
rect 195326 196718 195562 196954
rect 195646 196718 195882 196954
rect 195326 196398 195562 196634
rect 195646 196398 195882 196634
rect 195326 160718 195562 160954
rect 195646 160718 195882 160954
rect 195326 160398 195562 160634
rect 195646 160398 195882 160634
rect 195326 124718 195562 124954
rect 195646 124718 195882 124954
rect 195326 124398 195562 124634
rect 195646 124398 195882 124634
rect 114326 115718 114562 115954
rect 114646 115718 114882 115954
rect 114326 115398 114562 115634
rect 114646 115398 114882 115634
rect 139610 115718 139846 115954
rect 139610 115398 139846 115634
rect 170330 115718 170566 115954
rect 170330 115398 170566 115634
rect 124250 111218 124486 111454
rect 124250 110898 124486 111134
rect 154970 111218 155206 111454
rect 154970 110898 155206 111134
rect 185690 111218 185926 111454
rect 185690 110898 185926 111134
rect 195326 88718 195562 88954
rect 195646 88718 195882 88954
rect 195326 88398 195562 88634
rect 195646 88398 195882 88634
rect 114326 79718 114562 79954
rect 114646 79718 114882 79954
rect 114326 79398 114562 79634
rect 114646 79398 114882 79634
rect 114326 43718 114562 43954
rect 114646 43718 114882 43954
rect 114326 43398 114562 43634
rect 114646 43398 114882 43634
rect 114326 7718 114562 7954
rect 114646 7718 114882 7954
rect 114326 7398 114562 7634
rect 114646 7398 114882 7634
rect 114326 -1542 114562 -1306
rect 114646 -1542 114882 -1306
rect 114326 -1862 114562 -1626
rect 114646 -1862 114882 -1626
rect 118826 48218 119062 48454
rect 119146 48218 119382 48454
rect 118826 47898 119062 48134
rect 119146 47898 119382 48134
rect 118826 12218 119062 12454
rect 119146 12218 119382 12454
rect 118826 11898 119062 12134
rect 119146 11898 119382 12134
rect 118826 -2502 119062 -2266
rect 119146 -2502 119382 -2266
rect 118826 -2822 119062 -2586
rect 119146 -2822 119382 -2586
rect 123326 52718 123562 52954
rect 123646 52718 123882 52954
rect 123326 52398 123562 52634
rect 123646 52398 123882 52634
rect 123326 16718 123562 16954
rect 123646 16718 123882 16954
rect 123326 16398 123562 16634
rect 123646 16398 123882 16634
rect 123326 -3462 123562 -3226
rect 123646 -3462 123882 -3226
rect 123326 -3782 123562 -3546
rect 123646 -3782 123882 -3546
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 132326 61718 132562 61954
rect 132646 61718 132882 61954
rect 132326 61398 132562 61634
rect 132646 61398 132882 61634
rect 132326 25718 132562 25954
rect 132646 25718 132882 25954
rect 132326 25398 132562 25634
rect 132646 25398 132882 25634
rect 127826 -4422 128062 -4186
rect 128146 -4422 128382 -4186
rect 127826 -4742 128062 -4506
rect 128146 -4742 128382 -4506
rect 136826 66218 137062 66454
rect 137146 66218 137382 66454
rect 136826 65898 137062 66134
rect 137146 65898 137382 66134
rect 136826 30218 137062 30454
rect 137146 30218 137382 30454
rect 136826 29898 137062 30134
rect 137146 29898 137382 30134
rect 132326 -5382 132562 -5146
rect 132646 -5382 132882 -5146
rect 132326 -5702 132562 -5466
rect 132646 -5702 132882 -5466
rect 141326 70718 141562 70954
rect 141646 70718 141882 70954
rect 141326 70398 141562 70634
rect 141646 70398 141882 70634
rect 141326 34718 141562 34954
rect 141646 34718 141882 34954
rect 141326 34398 141562 34634
rect 141646 34398 141882 34634
rect 136826 -6342 137062 -6106
rect 137146 -6342 137382 -6106
rect 136826 -6662 137062 -6426
rect 137146 -6662 137382 -6426
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 150326 43718 150562 43954
rect 150646 43718 150882 43954
rect 150326 43398 150562 43634
rect 150646 43398 150882 43634
rect 150326 7718 150562 7954
rect 150646 7718 150882 7954
rect 150326 7398 150562 7634
rect 150646 7398 150882 7634
rect 141326 -7302 141562 -7066
rect 141646 -7302 141882 -7066
rect 141326 -7622 141562 -7386
rect 141646 -7622 141882 -7386
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 154826 48218 155062 48454
rect 155146 48218 155382 48454
rect 154826 47898 155062 48134
rect 155146 47898 155382 48134
rect 154826 12218 155062 12454
rect 155146 12218 155382 12454
rect 154826 11898 155062 12134
rect 155146 11898 155382 12134
rect 150326 -1542 150562 -1306
rect 150646 -1542 150882 -1306
rect 150326 -1862 150562 -1626
rect 150646 -1862 150882 -1626
rect 159326 52718 159562 52954
rect 159646 52718 159882 52954
rect 159326 52398 159562 52634
rect 159646 52398 159882 52634
rect 159326 16718 159562 16954
rect 159646 16718 159882 16954
rect 159326 16398 159562 16634
rect 159646 16398 159882 16634
rect 154826 -2502 155062 -2266
rect 155146 -2502 155382 -2266
rect 154826 -2822 155062 -2586
rect 155146 -2822 155382 -2586
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 159326 -3462 159562 -3226
rect 159646 -3462 159882 -3226
rect 159326 -3782 159562 -3546
rect 159646 -3782 159882 -3546
rect 168326 61718 168562 61954
rect 168646 61718 168882 61954
rect 168326 61398 168562 61634
rect 168646 61398 168882 61634
rect 168326 25718 168562 25954
rect 168646 25718 168882 25954
rect 168326 25398 168562 25634
rect 168646 25398 168882 25634
rect 163826 -4422 164062 -4186
rect 164146 -4422 164382 -4186
rect 163826 -4742 164062 -4506
rect 164146 -4742 164382 -4506
rect 172826 66218 173062 66454
rect 173146 66218 173382 66454
rect 172826 65898 173062 66134
rect 173146 65898 173382 66134
rect 172826 30218 173062 30454
rect 173146 30218 173382 30454
rect 172826 29898 173062 30134
rect 173146 29898 173382 30134
rect 168326 -5382 168562 -5146
rect 168646 -5382 168882 -5146
rect 168326 -5702 168562 -5466
rect 168646 -5702 168882 -5466
rect 177326 70718 177562 70954
rect 177646 70718 177882 70954
rect 177326 70398 177562 70634
rect 177646 70398 177882 70634
rect 177326 34718 177562 34954
rect 177646 34718 177882 34954
rect 177326 34398 177562 34634
rect 177646 34398 177882 34634
rect 172826 -6342 173062 -6106
rect 173146 -6342 173382 -6106
rect 172826 -6662 173062 -6426
rect 173146 -6662 173382 -6426
rect 177326 -7302 177562 -7066
rect 177646 -7302 177882 -7066
rect 177326 -7622 177562 -7386
rect 177646 -7622 177882 -7386
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 186326 43718 186562 43954
rect 186646 43718 186882 43954
rect 186326 43398 186562 43634
rect 186646 43398 186882 43634
rect 186326 7718 186562 7954
rect 186646 7718 186882 7954
rect 186326 7398 186562 7634
rect 186646 7398 186882 7634
rect 186326 -1542 186562 -1306
rect 186646 -1542 186882 -1306
rect 186326 -1862 186562 -1626
rect 186646 -1862 186882 -1626
rect 190826 48218 191062 48454
rect 191146 48218 191382 48454
rect 190826 47898 191062 48134
rect 191146 47898 191382 48134
rect 190826 12218 191062 12454
rect 191146 12218 191382 12454
rect 190826 11898 191062 12134
rect 191146 11898 191382 12134
rect 190826 -2502 191062 -2266
rect 191146 -2502 191382 -2266
rect 190826 -2822 191062 -2586
rect 191146 -2822 191382 -2586
rect 195326 52718 195562 52954
rect 195646 52718 195882 52954
rect 195326 52398 195562 52634
rect 195646 52398 195882 52634
rect 195326 16718 195562 16954
rect 195646 16718 195882 16954
rect 195326 16398 195562 16634
rect 195646 16398 195882 16634
rect 195326 -3462 195562 -3226
rect 195646 -3462 195882 -3226
rect 195326 -3782 195562 -3546
rect 195646 -3782 195882 -3546
rect 199826 708442 200062 708678
rect 200146 708442 200382 708678
rect 199826 708122 200062 708358
rect 200146 708122 200382 708358
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -4422 200062 -4186
rect 200146 -4422 200382 -4186
rect 199826 -4742 200062 -4506
rect 200146 -4742 200382 -4506
rect 204326 709402 204562 709638
rect 204646 709402 204882 709638
rect 204326 709082 204562 709318
rect 204646 709082 204882 709318
rect 204326 673718 204562 673954
rect 204646 673718 204882 673954
rect 204326 673398 204562 673634
rect 204646 673398 204882 673634
rect 204326 637718 204562 637954
rect 204646 637718 204882 637954
rect 204326 637398 204562 637634
rect 204646 637398 204882 637634
rect 204326 601718 204562 601954
rect 204646 601718 204882 601954
rect 204326 601398 204562 601634
rect 204646 601398 204882 601634
rect 204326 565718 204562 565954
rect 204646 565718 204882 565954
rect 204326 565398 204562 565634
rect 204646 565398 204882 565634
rect 204326 529718 204562 529954
rect 204646 529718 204882 529954
rect 204326 529398 204562 529634
rect 204646 529398 204882 529634
rect 204326 493718 204562 493954
rect 204646 493718 204882 493954
rect 204326 493398 204562 493634
rect 204646 493398 204882 493634
rect 204326 457718 204562 457954
rect 204646 457718 204882 457954
rect 204326 457398 204562 457634
rect 204646 457398 204882 457634
rect 204326 421718 204562 421954
rect 204646 421718 204882 421954
rect 204326 421398 204562 421634
rect 204646 421398 204882 421634
rect 204326 385718 204562 385954
rect 204646 385718 204882 385954
rect 204326 385398 204562 385634
rect 204646 385398 204882 385634
rect 204326 349718 204562 349954
rect 204646 349718 204882 349954
rect 204326 349398 204562 349634
rect 204646 349398 204882 349634
rect 204326 313718 204562 313954
rect 204646 313718 204882 313954
rect 204326 313398 204562 313634
rect 204646 313398 204882 313634
rect 204326 277718 204562 277954
rect 204646 277718 204882 277954
rect 204326 277398 204562 277634
rect 204646 277398 204882 277634
rect 204326 241718 204562 241954
rect 204646 241718 204882 241954
rect 204326 241398 204562 241634
rect 204646 241398 204882 241634
rect 204326 205718 204562 205954
rect 204646 205718 204882 205954
rect 204326 205398 204562 205634
rect 204646 205398 204882 205634
rect 204326 169718 204562 169954
rect 204646 169718 204882 169954
rect 204326 169398 204562 169634
rect 204646 169398 204882 169634
rect 204326 133718 204562 133954
rect 204646 133718 204882 133954
rect 204326 133398 204562 133634
rect 204646 133398 204882 133634
rect 204326 97718 204562 97954
rect 204646 97718 204882 97954
rect 204326 97398 204562 97634
rect 204646 97398 204882 97634
rect 204326 61718 204562 61954
rect 204646 61718 204882 61954
rect 204326 61398 204562 61634
rect 204646 61398 204882 61634
rect 204326 25718 204562 25954
rect 204646 25718 204882 25954
rect 204326 25398 204562 25634
rect 204646 25398 204882 25634
rect 204326 -5382 204562 -5146
rect 204646 -5382 204882 -5146
rect 204326 -5702 204562 -5466
rect 204646 -5702 204882 -5466
rect 208826 710362 209062 710598
rect 209146 710362 209382 710598
rect 208826 710042 209062 710278
rect 209146 710042 209382 710278
rect 208826 678218 209062 678454
rect 209146 678218 209382 678454
rect 208826 677898 209062 678134
rect 209146 677898 209382 678134
rect 208826 642218 209062 642454
rect 209146 642218 209382 642454
rect 208826 641898 209062 642134
rect 209146 641898 209382 642134
rect 208826 606218 209062 606454
rect 209146 606218 209382 606454
rect 208826 605898 209062 606134
rect 209146 605898 209382 606134
rect 208826 570218 209062 570454
rect 209146 570218 209382 570454
rect 208826 569898 209062 570134
rect 209146 569898 209382 570134
rect 208826 534218 209062 534454
rect 209146 534218 209382 534454
rect 208826 533898 209062 534134
rect 209146 533898 209382 534134
rect 208826 498218 209062 498454
rect 209146 498218 209382 498454
rect 208826 497898 209062 498134
rect 209146 497898 209382 498134
rect 208826 462218 209062 462454
rect 209146 462218 209382 462454
rect 208826 461898 209062 462134
rect 209146 461898 209382 462134
rect 208826 426218 209062 426454
rect 209146 426218 209382 426454
rect 208826 425898 209062 426134
rect 209146 425898 209382 426134
rect 208826 390218 209062 390454
rect 209146 390218 209382 390454
rect 208826 389898 209062 390134
rect 209146 389898 209382 390134
rect 208826 354218 209062 354454
rect 209146 354218 209382 354454
rect 208826 353898 209062 354134
rect 209146 353898 209382 354134
rect 208826 318218 209062 318454
rect 209146 318218 209382 318454
rect 208826 317898 209062 318134
rect 209146 317898 209382 318134
rect 208826 282218 209062 282454
rect 209146 282218 209382 282454
rect 208826 281898 209062 282134
rect 209146 281898 209382 282134
rect 208826 246218 209062 246454
rect 209146 246218 209382 246454
rect 208826 245898 209062 246134
rect 209146 245898 209382 246134
rect 208826 210218 209062 210454
rect 209146 210218 209382 210454
rect 208826 209898 209062 210134
rect 209146 209898 209382 210134
rect 208826 174218 209062 174454
rect 209146 174218 209382 174454
rect 208826 173898 209062 174134
rect 209146 173898 209382 174134
rect 208826 138218 209062 138454
rect 209146 138218 209382 138454
rect 208826 137898 209062 138134
rect 209146 137898 209382 138134
rect 208826 102218 209062 102454
rect 209146 102218 209382 102454
rect 208826 101898 209062 102134
rect 209146 101898 209382 102134
rect 208826 66218 209062 66454
rect 209146 66218 209382 66454
rect 208826 65898 209062 66134
rect 209146 65898 209382 66134
rect 208826 30218 209062 30454
rect 209146 30218 209382 30454
rect 208826 29898 209062 30134
rect 209146 29898 209382 30134
rect 208826 -6342 209062 -6106
rect 209146 -6342 209382 -6106
rect 208826 -6662 209062 -6426
rect 209146 -6662 209382 -6426
rect 213326 711322 213562 711558
rect 213646 711322 213882 711558
rect 213326 711002 213562 711238
rect 213646 711002 213882 711238
rect 213326 682718 213562 682954
rect 213646 682718 213882 682954
rect 213326 682398 213562 682634
rect 213646 682398 213882 682634
rect 213326 646718 213562 646954
rect 213646 646718 213882 646954
rect 213326 646398 213562 646634
rect 213646 646398 213882 646634
rect 213326 610718 213562 610954
rect 213646 610718 213882 610954
rect 213326 610398 213562 610634
rect 213646 610398 213882 610634
rect 213326 574718 213562 574954
rect 213646 574718 213882 574954
rect 213326 574398 213562 574634
rect 213646 574398 213882 574634
rect 213326 538718 213562 538954
rect 213646 538718 213882 538954
rect 213326 538398 213562 538634
rect 213646 538398 213882 538634
rect 213326 502718 213562 502954
rect 213646 502718 213882 502954
rect 213326 502398 213562 502634
rect 213646 502398 213882 502634
rect 213326 466718 213562 466954
rect 213646 466718 213882 466954
rect 213326 466398 213562 466634
rect 213646 466398 213882 466634
rect 213326 430718 213562 430954
rect 213646 430718 213882 430954
rect 213326 430398 213562 430634
rect 213646 430398 213882 430634
rect 213326 394718 213562 394954
rect 213646 394718 213882 394954
rect 213326 394398 213562 394634
rect 213646 394398 213882 394634
rect 213326 358718 213562 358954
rect 213646 358718 213882 358954
rect 213326 358398 213562 358634
rect 213646 358398 213882 358634
rect 213326 322718 213562 322954
rect 213646 322718 213882 322954
rect 213326 322398 213562 322634
rect 213646 322398 213882 322634
rect 213326 286718 213562 286954
rect 213646 286718 213882 286954
rect 213326 286398 213562 286634
rect 213646 286398 213882 286634
rect 213326 250718 213562 250954
rect 213646 250718 213882 250954
rect 213326 250398 213562 250634
rect 213646 250398 213882 250634
rect 213326 214718 213562 214954
rect 213646 214718 213882 214954
rect 213326 214398 213562 214634
rect 213646 214398 213882 214634
rect 213326 178718 213562 178954
rect 213646 178718 213882 178954
rect 213326 178398 213562 178634
rect 213646 178398 213882 178634
rect 213326 142718 213562 142954
rect 213646 142718 213882 142954
rect 213326 142398 213562 142634
rect 213646 142398 213882 142634
rect 213326 106718 213562 106954
rect 213646 106718 213882 106954
rect 213326 106398 213562 106634
rect 213646 106398 213882 106634
rect 213326 70718 213562 70954
rect 213646 70718 213882 70954
rect 213326 70398 213562 70634
rect 213646 70398 213882 70634
rect 213326 34718 213562 34954
rect 213646 34718 213882 34954
rect 213326 34398 213562 34634
rect 213646 34398 213882 34634
rect 213326 -7302 213562 -7066
rect 213646 -7302 213882 -7066
rect 213326 -7622 213562 -7386
rect 213646 -7622 213882 -7386
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 222326 705562 222562 705798
rect 222646 705562 222882 705798
rect 222326 705242 222562 705478
rect 222646 705242 222882 705478
rect 222326 691718 222562 691954
rect 222646 691718 222882 691954
rect 222326 691398 222562 691634
rect 222646 691398 222882 691634
rect 222326 655718 222562 655954
rect 222646 655718 222882 655954
rect 222326 655398 222562 655634
rect 222646 655398 222882 655634
rect 222326 619718 222562 619954
rect 222646 619718 222882 619954
rect 222326 619398 222562 619634
rect 222646 619398 222882 619634
rect 222326 583718 222562 583954
rect 222646 583718 222882 583954
rect 222326 583398 222562 583634
rect 222646 583398 222882 583634
rect 222326 547718 222562 547954
rect 222646 547718 222882 547954
rect 222326 547398 222562 547634
rect 222646 547398 222882 547634
rect 222326 511718 222562 511954
rect 222646 511718 222882 511954
rect 222326 511398 222562 511634
rect 222646 511398 222882 511634
rect 222326 475718 222562 475954
rect 222646 475718 222882 475954
rect 222326 475398 222562 475634
rect 222646 475398 222882 475634
rect 222326 439718 222562 439954
rect 222646 439718 222882 439954
rect 222326 439398 222562 439634
rect 222646 439398 222882 439634
rect 222326 403718 222562 403954
rect 222646 403718 222882 403954
rect 222326 403398 222562 403634
rect 222646 403398 222882 403634
rect 222326 367718 222562 367954
rect 222646 367718 222882 367954
rect 222326 367398 222562 367634
rect 222646 367398 222882 367634
rect 222326 331718 222562 331954
rect 222646 331718 222882 331954
rect 222326 331398 222562 331634
rect 222646 331398 222882 331634
rect 222326 295718 222562 295954
rect 222646 295718 222882 295954
rect 222326 295398 222562 295634
rect 222646 295398 222882 295634
rect 222326 259718 222562 259954
rect 222646 259718 222882 259954
rect 222326 259398 222562 259634
rect 222646 259398 222882 259634
rect 222326 223718 222562 223954
rect 222646 223718 222882 223954
rect 222326 223398 222562 223634
rect 222646 223398 222882 223634
rect 222326 187718 222562 187954
rect 222646 187718 222882 187954
rect 222326 187398 222562 187634
rect 222646 187398 222882 187634
rect 222326 151718 222562 151954
rect 222646 151718 222882 151954
rect 222326 151398 222562 151634
rect 222646 151398 222882 151634
rect 222326 115718 222562 115954
rect 222646 115718 222882 115954
rect 222326 115398 222562 115634
rect 222646 115398 222882 115634
rect 222326 79718 222562 79954
rect 222646 79718 222882 79954
rect 222326 79398 222562 79634
rect 222646 79398 222882 79634
rect 222326 43718 222562 43954
rect 222646 43718 222882 43954
rect 222326 43398 222562 43634
rect 222646 43398 222882 43634
rect 222326 7718 222562 7954
rect 222646 7718 222882 7954
rect 222326 7398 222562 7634
rect 222646 7398 222882 7634
rect 222326 -1542 222562 -1306
rect 222646 -1542 222882 -1306
rect 222326 -1862 222562 -1626
rect 222646 -1862 222882 -1626
rect 226826 706522 227062 706758
rect 227146 706522 227382 706758
rect 226826 706202 227062 706438
rect 227146 706202 227382 706438
rect 226826 696218 227062 696454
rect 227146 696218 227382 696454
rect 226826 695898 227062 696134
rect 227146 695898 227382 696134
rect 226826 660218 227062 660454
rect 227146 660218 227382 660454
rect 226826 659898 227062 660134
rect 227146 659898 227382 660134
rect 226826 624218 227062 624454
rect 227146 624218 227382 624454
rect 226826 623898 227062 624134
rect 227146 623898 227382 624134
rect 226826 588218 227062 588454
rect 227146 588218 227382 588454
rect 226826 587898 227062 588134
rect 227146 587898 227382 588134
rect 226826 552218 227062 552454
rect 227146 552218 227382 552454
rect 226826 551898 227062 552134
rect 227146 551898 227382 552134
rect 226826 516218 227062 516454
rect 227146 516218 227382 516454
rect 226826 515898 227062 516134
rect 227146 515898 227382 516134
rect 226826 480218 227062 480454
rect 227146 480218 227382 480454
rect 226826 479898 227062 480134
rect 227146 479898 227382 480134
rect 226826 444218 227062 444454
rect 227146 444218 227382 444454
rect 226826 443898 227062 444134
rect 227146 443898 227382 444134
rect 226826 408218 227062 408454
rect 227146 408218 227382 408454
rect 226826 407898 227062 408134
rect 227146 407898 227382 408134
rect 226826 372218 227062 372454
rect 227146 372218 227382 372454
rect 226826 371898 227062 372134
rect 227146 371898 227382 372134
rect 226826 336218 227062 336454
rect 227146 336218 227382 336454
rect 226826 335898 227062 336134
rect 227146 335898 227382 336134
rect 226826 300218 227062 300454
rect 227146 300218 227382 300454
rect 226826 299898 227062 300134
rect 227146 299898 227382 300134
rect 226826 264218 227062 264454
rect 227146 264218 227382 264454
rect 226826 263898 227062 264134
rect 227146 263898 227382 264134
rect 226826 228218 227062 228454
rect 227146 228218 227382 228454
rect 226826 227898 227062 228134
rect 227146 227898 227382 228134
rect 226826 192218 227062 192454
rect 227146 192218 227382 192454
rect 226826 191898 227062 192134
rect 227146 191898 227382 192134
rect 226826 156218 227062 156454
rect 227146 156218 227382 156454
rect 226826 155898 227062 156134
rect 227146 155898 227382 156134
rect 226826 120218 227062 120454
rect 227146 120218 227382 120454
rect 226826 119898 227062 120134
rect 227146 119898 227382 120134
rect 226826 84218 227062 84454
rect 227146 84218 227382 84454
rect 226826 83898 227062 84134
rect 227146 83898 227382 84134
rect 226826 48218 227062 48454
rect 227146 48218 227382 48454
rect 226826 47898 227062 48134
rect 227146 47898 227382 48134
rect 226826 12218 227062 12454
rect 227146 12218 227382 12454
rect 226826 11898 227062 12134
rect 227146 11898 227382 12134
rect 226826 -2502 227062 -2266
rect 227146 -2502 227382 -2266
rect 226826 -2822 227062 -2586
rect 227146 -2822 227382 -2586
rect 231326 707482 231562 707718
rect 231646 707482 231882 707718
rect 231326 707162 231562 707398
rect 231646 707162 231882 707398
rect 231326 700718 231562 700954
rect 231646 700718 231882 700954
rect 231326 700398 231562 700634
rect 231646 700398 231882 700634
rect 231326 664718 231562 664954
rect 231646 664718 231882 664954
rect 231326 664398 231562 664634
rect 231646 664398 231882 664634
rect 231326 628718 231562 628954
rect 231646 628718 231882 628954
rect 231326 628398 231562 628634
rect 231646 628398 231882 628634
rect 231326 592718 231562 592954
rect 231646 592718 231882 592954
rect 231326 592398 231562 592634
rect 231646 592398 231882 592634
rect 231326 556718 231562 556954
rect 231646 556718 231882 556954
rect 231326 556398 231562 556634
rect 231646 556398 231882 556634
rect 231326 520718 231562 520954
rect 231646 520718 231882 520954
rect 231326 520398 231562 520634
rect 231646 520398 231882 520634
rect 231326 484718 231562 484954
rect 231646 484718 231882 484954
rect 231326 484398 231562 484634
rect 231646 484398 231882 484634
rect 231326 448718 231562 448954
rect 231646 448718 231882 448954
rect 231326 448398 231562 448634
rect 231646 448398 231882 448634
rect 231326 412718 231562 412954
rect 231646 412718 231882 412954
rect 231326 412398 231562 412634
rect 231646 412398 231882 412634
rect 231326 376718 231562 376954
rect 231646 376718 231882 376954
rect 231326 376398 231562 376634
rect 231646 376398 231882 376634
rect 231326 340718 231562 340954
rect 231646 340718 231882 340954
rect 231326 340398 231562 340634
rect 231646 340398 231882 340634
rect 231326 304718 231562 304954
rect 231646 304718 231882 304954
rect 231326 304398 231562 304634
rect 231646 304398 231882 304634
rect 231326 268718 231562 268954
rect 231646 268718 231882 268954
rect 231326 268398 231562 268634
rect 231646 268398 231882 268634
rect 231326 232718 231562 232954
rect 231646 232718 231882 232954
rect 231326 232398 231562 232634
rect 231646 232398 231882 232634
rect 231326 196718 231562 196954
rect 231646 196718 231882 196954
rect 231326 196398 231562 196634
rect 231646 196398 231882 196634
rect 231326 160718 231562 160954
rect 231646 160718 231882 160954
rect 231326 160398 231562 160634
rect 231646 160398 231882 160634
rect 231326 124718 231562 124954
rect 231646 124718 231882 124954
rect 231326 124398 231562 124634
rect 231646 124398 231882 124634
rect 231326 88718 231562 88954
rect 231646 88718 231882 88954
rect 231326 88398 231562 88634
rect 231646 88398 231882 88634
rect 231326 52718 231562 52954
rect 231646 52718 231882 52954
rect 231326 52398 231562 52634
rect 231646 52398 231882 52634
rect 231326 16718 231562 16954
rect 231646 16718 231882 16954
rect 231326 16398 231562 16634
rect 231646 16398 231882 16634
rect 231326 -3462 231562 -3226
rect 231646 -3462 231882 -3226
rect 231326 -3782 231562 -3546
rect 231646 -3782 231882 -3546
rect 235826 708442 236062 708678
rect 236146 708442 236382 708678
rect 235826 708122 236062 708358
rect 236146 708122 236382 708358
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 235826 273218 236062 273454
rect 236146 273218 236382 273454
rect 235826 272898 236062 273134
rect 236146 272898 236382 273134
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -4422 236062 -4186
rect 236146 -4422 236382 -4186
rect 235826 -4742 236062 -4506
rect 236146 -4742 236382 -4506
rect 240326 709402 240562 709638
rect 240646 709402 240882 709638
rect 240326 709082 240562 709318
rect 240646 709082 240882 709318
rect 240326 673718 240562 673954
rect 240646 673718 240882 673954
rect 240326 673398 240562 673634
rect 240646 673398 240882 673634
rect 240326 637718 240562 637954
rect 240646 637718 240882 637954
rect 240326 637398 240562 637634
rect 240646 637398 240882 637634
rect 240326 601718 240562 601954
rect 240646 601718 240882 601954
rect 240326 601398 240562 601634
rect 240646 601398 240882 601634
rect 240326 565718 240562 565954
rect 240646 565718 240882 565954
rect 240326 565398 240562 565634
rect 240646 565398 240882 565634
rect 240326 529718 240562 529954
rect 240646 529718 240882 529954
rect 240326 529398 240562 529634
rect 240646 529398 240882 529634
rect 240326 493718 240562 493954
rect 240646 493718 240882 493954
rect 240326 493398 240562 493634
rect 240646 493398 240882 493634
rect 240326 457718 240562 457954
rect 240646 457718 240882 457954
rect 240326 457398 240562 457634
rect 240646 457398 240882 457634
rect 240326 421718 240562 421954
rect 240646 421718 240882 421954
rect 240326 421398 240562 421634
rect 240646 421398 240882 421634
rect 240326 385718 240562 385954
rect 240646 385718 240882 385954
rect 240326 385398 240562 385634
rect 240646 385398 240882 385634
rect 240326 349718 240562 349954
rect 240646 349718 240882 349954
rect 240326 349398 240562 349634
rect 240646 349398 240882 349634
rect 240326 313718 240562 313954
rect 240646 313718 240882 313954
rect 240326 313398 240562 313634
rect 240646 313398 240882 313634
rect 240326 277718 240562 277954
rect 240646 277718 240882 277954
rect 240326 277398 240562 277634
rect 240646 277398 240882 277634
rect 240326 241718 240562 241954
rect 240646 241718 240882 241954
rect 240326 241398 240562 241634
rect 240646 241398 240882 241634
rect 240326 205718 240562 205954
rect 240646 205718 240882 205954
rect 240326 205398 240562 205634
rect 240646 205398 240882 205634
rect 240326 169718 240562 169954
rect 240646 169718 240882 169954
rect 240326 169398 240562 169634
rect 240646 169398 240882 169634
rect 240326 133718 240562 133954
rect 240646 133718 240882 133954
rect 240326 133398 240562 133634
rect 240646 133398 240882 133634
rect 240326 97718 240562 97954
rect 240646 97718 240882 97954
rect 240326 97398 240562 97634
rect 240646 97398 240882 97634
rect 240326 61718 240562 61954
rect 240646 61718 240882 61954
rect 240326 61398 240562 61634
rect 240646 61398 240882 61634
rect 240326 25718 240562 25954
rect 240646 25718 240882 25954
rect 240326 25398 240562 25634
rect 240646 25398 240882 25634
rect 240326 -5382 240562 -5146
rect 240646 -5382 240882 -5146
rect 240326 -5702 240562 -5466
rect 240646 -5702 240882 -5466
rect 244826 710362 245062 710598
rect 245146 710362 245382 710598
rect 244826 710042 245062 710278
rect 245146 710042 245382 710278
rect 244826 678218 245062 678454
rect 245146 678218 245382 678454
rect 244826 677898 245062 678134
rect 245146 677898 245382 678134
rect 244826 642218 245062 642454
rect 245146 642218 245382 642454
rect 244826 641898 245062 642134
rect 245146 641898 245382 642134
rect 244826 606218 245062 606454
rect 245146 606218 245382 606454
rect 244826 605898 245062 606134
rect 245146 605898 245382 606134
rect 244826 570218 245062 570454
rect 245146 570218 245382 570454
rect 244826 569898 245062 570134
rect 245146 569898 245382 570134
rect 244826 534218 245062 534454
rect 245146 534218 245382 534454
rect 244826 533898 245062 534134
rect 245146 533898 245382 534134
rect 244826 498218 245062 498454
rect 245146 498218 245382 498454
rect 244826 497898 245062 498134
rect 245146 497898 245382 498134
rect 244826 462218 245062 462454
rect 245146 462218 245382 462454
rect 244826 461898 245062 462134
rect 245146 461898 245382 462134
rect 244826 426218 245062 426454
rect 245146 426218 245382 426454
rect 244826 425898 245062 426134
rect 245146 425898 245382 426134
rect 244826 390218 245062 390454
rect 245146 390218 245382 390454
rect 244826 389898 245062 390134
rect 245146 389898 245382 390134
rect 244826 354218 245062 354454
rect 245146 354218 245382 354454
rect 244826 353898 245062 354134
rect 245146 353898 245382 354134
rect 244826 318218 245062 318454
rect 245146 318218 245382 318454
rect 244826 317898 245062 318134
rect 245146 317898 245382 318134
rect 244826 282218 245062 282454
rect 245146 282218 245382 282454
rect 244826 281898 245062 282134
rect 245146 281898 245382 282134
rect 244826 246218 245062 246454
rect 245146 246218 245382 246454
rect 244826 245898 245062 246134
rect 245146 245898 245382 246134
rect 244826 210218 245062 210454
rect 245146 210218 245382 210454
rect 244826 209898 245062 210134
rect 245146 209898 245382 210134
rect 244826 174218 245062 174454
rect 245146 174218 245382 174454
rect 244826 173898 245062 174134
rect 245146 173898 245382 174134
rect 244826 138218 245062 138454
rect 245146 138218 245382 138454
rect 244826 137898 245062 138134
rect 245146 137898 245382 138134
rect 244826 102218 245062 102454
rect 245146 102218 245382 102454
rect 244826 101898 245062 102134
rect 245146 101898 245382 102134
rect 244826 66218 245062 66454
rect 245146 66218 245382 66454
rect 244826 65898 245062 66134
rect 245146 65898 245382 66134
rect 244826 30218 245062 30454
rect 245146 30218 245382 30454
rect 244826 29898 245062 30134
rect 245146 29898 245382 30134
rect 244826 -6342 245062 -6106
rect 245146 -6342 245382 -6106
rect 244826 -6662 245062 -6426
rect 245146 -6662 245382 -6426
rect 249326 711322 249562 711558
rect 249646 711322 249882 711558
rect 249326 711002 249562 711238
rect 249646 711002 249882 711238
rect 249326 682718 249562 682954
rect 249646 682718 249882 682954
rect 249326 682398 249562 682634
rect 249646 682398 249882 682634
rect 249326 646718 249562 646954
rect 249646 646718 249882 646954
rect 249326 646398 249562 646634
rect 249646 646398 249882 646634
rect 249326 610718 249562 610954
rect 249646 610718 249882 610954
rect 249326 610398 249562 610634
rect 249646 610398 249882 610634
rect 249326 574718 249562 574954
rect 249646 574718 249882 574954
rect 249326 574398 249562 574634
rect 249646 574398 249882 574634
rect 249326 538718 249562 538954
rect 249646 538718 249882 538954
rect 249326 538398 249562 538634
rect 249646 538398 249882 538634
rect 249326 502718 249562 502954
rect 249646 502718 249882 502954
rect 249326 502398 249562 502634
rect 249646 502398 249882 502634
rect 249326 466718 249562 466954
rect 249646 466718 249882 466954
rect 249326 466398 249562 466634
rect 249646 466398 249882 466634
rect 249326 430718 249562 430954
rect 249646 430718 249882 430954
rect 249326 430398 249562 430634
rect 249646 430398 249882 430634
rect 249326 394718 249562 394954
rect 249646 394718 249882 394954
rect 249326 394398 249562 394634
rect 249646 394398 249882 394634
rect 249326 358718 249562 358954
rect 249646 358718 249882 358954
rect 249326 358398 249562 358634
rect 249646 358398 249882 358634
rect 249326 322718 249562 322954
rect 249646 322718 249882 322954
rect 249326 322398 249562 322634
rect 249646 322398 249882 322634
rect 249326 286718 249562 286954
rect 249646 286718 249882 286954
rect 249326 286398 249562 286634
rect 249646 286398 249882 286634
rect 249326 250718 249562 250954
rect 249646 250718 249882 250954
rect 249326 250398 249562 250634
rect 249646 250398 249882 250634
rect 249326 214718 249562 214954
rect 249646 214718 249882 214954
rect 249326 214398 249562 214634
rect 249646 214398 249882 214634
rect 249326 178718 249562 178954
rect 249646 178718 249882 178954
rect 249326 178398 249562 178634
rect 249646 178398 249882 178634
rect 249326 142718 249562 142954
rect 249646 142718 249882 142954
rect 249326 142398 249562 142634
rect 249646 142398 249882 142634
rect 249326 106718 249562 106954
rect 249646 106718 249882 106954
rect 249326 106398 249562 106634
rect 249646 106398 249882 106634
rect 249326 70718 249562 70954
rect 249646 70718 249882 70954
rect 249326 70398 249562 70634
rect 249646 70398 249882 70634
rect 249326 34718 249562 34954
rect 249646 34718 249882 34954
rect 249326 34398 249562 34634
rect 249646 34398 249882 34634
rect 249326 -7302 249562 -7066
rect 249646 -7302 249882 -7066
rect 249326 -7622 249562 -7386
rect 249646 -7622 249882 -7386
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 258326 705562 258562 705798
rect 258646 705562 258882 705798
rect 258326 705242 258562 705478
rect 258646 705242 258882 705478
rect 258326 691718 258562 691954
rect 258646 691718 258882 691954
rect 258326 691398 258562 691634
rect 258646 691398 258882 691634
rect 258326 655718 258562 655954
rect 258646 655718 258882 655954
rect 258326 655398 258562 655634
rect 258646 655398 258882 655634
rect 258326 619718 258562 619954
rect 258646 619718 258882 619954
rect 258326 619398 258562 619634
rect 258646 619398 258882 619634
rect 258326 583718 258562 583954
rect 258646 583718 258882 583954
rect 258326 583398 258562 583634
rect 258646 583398 258882 583634
rect 258326 547718 258562 547954
rect 258646 547718 258882 547954
rect 258326 547398 258562 547634
rect 258646 547398 258882 547634
rect 258326 511718 258562 511954
rect 258646 511718 258882 511954
rect 258326 511398 258562 511634
rect 258646 511398 258882 511634
rect 258326 475718 258562 475954
rect 258646 475718 258882 475954
rect 258326 475398 258562 475634
rect 258646 475398 258882 475634
rect 258326 439718 258562 439954
rect 258646 439718 258882 439954
rect 258326 439398 258562 439634
rect 258646 439398 258882 439634
rect 258326 403718 258562 403954
rect 258646 403718 258882 403954
rect 258326 403398 258562 403634
rect 258646 403398 258882 403634
rect 258326 367718 258562 367954
rect 258646 367718 258882 367954
rect 258326 367398 258562 367634
rect 258646 367398 258882 367634
rect 258326 331718 258562 331954
rect 258646 331718 258882 331954
rect 258326 331398 258562 331634
rect 258646 331398 258882 331634
rect 258326 295718 258562 295954
rect 258646 295718 258882 295954
rect 258326 295398 258562 295634
rect 258646 295398 258882 295634
rect 258326 259718 258562 259954
rect 258646 259718 258882 259954
rect 258326 259398 258562 259634
rect 258646 259398 258882 259634
rect 258326 223718 258562 223954
rect 258646 223718 258882 223954
rect 258326 223398 258562 223634
rect 258646 223398 258882 223634
rect 258326 187718 258562 187954
rect 258646 187718 258882 187954
rect 258326 187398 258562 187634
rect 258646 187398 258882 187634
rect 258326 151718 258562 151954
rect 258646 151718 258882 151954
rect 258326 151398 258562 151634
rect 258646 151398 258882 151634
rect 258326 115718 258562 115954
rect 258646 115718 258882 115954
rect 258326 115398 258562 115634
rect 258646 115398 258882 115634
rect 258326 79718 258562 79954
rect 258646 79718 258882 79954
rect 258326 79398 258562 79634
rect 258646 79398 258882 79634
rect 258326 43718 258562 43954
rect 258646 43718 258882 43954
rect 258326 43398 258562 43634
rect 258646 43398 258882 43634
rect 258326 7718 258562 7954
rect 258646 7718 258882 7954
rect 258326 7398 258562 7634
rect 258646 7398 258882 7634
rect 258326 -1542 258562 -1306
rect 258646 -1542 258882 -1306
rect 258326 -1862 258562 -1626
rect 258646 -1862 258882 -1626
rect 262826 706522 263062 706758
rect 263146 706522 263382 706758
rect 262826 706202 263062 706438
rect 263146 706202 263382 706438
rect 262826 696218 263062 696454
rect 263146 696218 263382 696454
rect 262826 695898 263062 696134
rect 263146 695898 263382 696134
rect 262826 660218 263062 660454
rect 263146 660218 263382 660454
rect 262826 659898 263062 660134
rect 263146 659898 263382 660134
rect 262826 624218 263062 624454
rect 263146 624218 263382 624454
rect 262826 623898 263062 624134
rect 263146 623898 263382 624134
rect 262826 588218 263062 588454
rect 263146 588218 263382 588454
rect 262826 587898 263062 588134
rect 263146 587898 263382 588134
rect 262826 552218 263062 552454
rect 263146 552218 263382 552454
rect 262826 551898 263062 552134
rect 263146 551898 263382 552134
rect 262826 516218 263062 516454
rect 263146 516218 263382 516454
rect 262826 515898 263062 516134
rect 263146 515898 263382 516134
rect 262826 480218 263062 480454
rect 263146 480218 263382 480454
rect 262826 479898 263062 480134
rect 263146 479898 263382 480134
rect 262826 444218 263062 444454
rect 263146 444218 263382 444454
rect 262826 443898 263062 444134
rect 263146 443898 263382 444134
rect 262826 408218 263062 408454
rect 263146 408218 263382 408454
rect 262826 407898 263062 408134
rect 263146 407898 263382 408134
rect 262826 372218 263062 372454
rect 263146 372218 263382 372454
rect 262826 371898 263062 372134
rect 263146 371898 263382 372134
rect 262826 336218 263062 336454
rect 263146 336218 263382 336454
rect 262826 335898 263062 336134
rect 263146 335898 263382 336134
rect 262826 300218 263062 300454
rect 263146 300218 263382 300454
rect 262826 299898 263062 300134
rect 263146 299898 263382 300134
rect 262826 264218 263062 264454
rect 263146 264218 263382 264454
rect 262826 263898 263062 264134
rect 263146 263898 263382 264134
rect 262826 228218 263062 228454
rect 263146 228218 263382 228454
rect 262826 227898 263062 228134
rect 263146 227898 263382 228134
rect 262826 192218 263062 192454
rect 263146 192218 263382 192454
rect 262826 191898 263062 192134
rect 263146 191898 263382 192134
rect 262826 156218 263062 156454
rect 263146 156218 263382 156454
rect 262826 155898 263062 156134
rect 263146 155898 263382 156134
rect 262826 120218 263062 120454
rect 263146 120218 263382 120454
rect 262826 119898 263062 120134
rect 263146 119898 263382 120134
rect 262826 84218 263062 84454
rect 263146 84218 263382 84454
rect 262826 83898 263062 84134
rect 263146 83898 263382 84134
rect 262826 48218 263062 48454
rect 263146 48218 263382 48454
rect 262826 47898 263062 48134
rect 263146 47898 263382 48134
rect 262826 12218 263062 12454
rect 263146 12218 263382 12454
rect 262826 11898 263062 12134
rect 263146 11898 263382 12134
rect 262826 -2502 263062 -2266
rect 263146 -2502 263382 -2266
rect 262826 -2822 263062 -2586
rect 263146 -2822 263382 -2586
rect 267326 707482 267562 707718
rect 267646 707482 267882 707718
rect 267326 707162 267562 707398
rect 267646 707162 267882 707398
rect 267326 700718 267562 700954
rect 267646 700718 267882 700954
rect 267326 700398 267562 700634
rect 267646 700398 267882 700634
rect 267326 664718 267562 664954
rect 267646 664718 267882 664954
rect 267326 664398 267562 664634
rect 267646 664398 267882 664634
rect 267326 628718 267562 628954
rect 267646 628718 267882 628954
rect 267326 628398 267562 628634
rect 267646 628398 267882 628634
rect 267326 592718 267562 592954
rect 267646 592718 267882 592954
rect 267326 592398 267562 592634
rect 267646 592398 267882 592634
rect 267326 556718 267562 556954
rect 267646 556718 267882 556954
rect 267326 556398 267562 556634
rect 267646 556398 267882 556634
rect 267326 520718 267562 520954
rect 267646 520718 267882 520954
rect 267326 520398 267562 520634
rect 267646 520398 267882 520634
rect 267326 484718 267562 484954
rect 267646 484718 267882 484954
rect 267326 484398 267562 484634
rect 267646 484398 267882 484634
rect 267326 448718 267562 448954
rect 267646 448718 267882 448954
rect 267326 448398 267562 448634
rect 267646 448398 267882 448634
rect 267326 412718 267562 412954
rect 267646 412718 267882 412954
rect 267326 412398 267562 412634
rect 267646 412398 267882 412634
rect 267326 376718 267562 376954
rect 267646 376718 267882 376954
rect 267326 376398 267562 376634
rect 267646 376398 267882 376634
rect 267326 340718 267562 340954
rect 267646 340718 267882 340954
rect 267326 340398 267562 340634
rect 267646 340398 267882 340634
rect 267326 304718 267562 304954
rect 267646 304718 267882 304954
rect 267326 304398 267562 304634
rect 267646 304398 267882 304634
rect 267326 268718 267562 268954
rect 267646 268718 267882 268954
rect 267326 268398 267562 268634
rect 267646 268398 267882 268634
rect 267326 232718 267562 232954
rect 267646 232718 267882 232954
rect 267326 232398 267562 232634
rect 267646 232398 267882 232634
rect 267326 196718 267562 196954
rect 267646 196718 267882 196954
rect 267326 196398 267562 196634
rect 267646 196398 267882 196634
rect 267326 160718 267562 160954
rect 267646 160718 267882 160954
rect 267326 160398 267562 160634
rect 267646 160398 267882 160634
rect 267326 124718 267562 124954
rect 267646 124718 267882 124954
rect 267326 124398 267562 124634
rect 267646 124398 267882 124634
rect 267326 88718 267562 88954
rect 267646 88718 267882 88954
rect 267326 88398 267562 88634
rect 267646 88398 267882 88634
rect 267326 52718 267562 52954
rect 267646 52718 267882 52954
rect 267326 52398 267562 52634
rect 267646 52398 267882 52634
rect 267326 16718 267562 16954
rect 267646 16718 267882 16954
rect 267326 16398 267562 16634
rect 267646 16398 267882 16634
rect 267326 -3462 267562 -3226
rect 267646 -3462 267882 -3226
rect 267326 -3782 267562 -3546
rect 267646 -3782 267882 -3546
rect 271826 708442 272062 708678
rect 272146 708442 272382 708678
rect 271826 708122 272062 708358
rect 272146 708122 272382 708358
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -4422 272062 -4186
rect 272146 -4422 272382 -4186
rect 271826 -4742 272062 -4506
rect 272146 -4742 272382 -4506
rect 276326 709402 276562 709638
rect 276646 709402 276882 709638
rect 276326 709082 276562 709318
rect 276646 709082 276882 709318
rect 276326 673718 276562 673954
rect 276646 673718 276882 673954
rect 276326 673398 276562 673634
rect 276646 673398 276882 673634
rect 276326 637718 276562 637954
rect 276646 637718 276882 637954
rect 276326 637398 276562 637634
rect 276646 637398 276882 637634
rect 276326 601718 276562 601954
rect 276646 601718 276882 601954
rect 276326 601398 276562 601634
rect 276646 601398 276882 601634
rect 276326 565718 276562 565954
rect 276646 565718 276882 565954
rect 276326 565398 276562 565634
rect 276646 565398 276882 565634
rect 276326 529718 276562 529954
rect 276646 529718 276882 529954
rect 276326 529398 276562 529634
rect 276646 529398 276882 529634
rect 276326 493718 276562 493954
rect 276646 493718 276882 493954
rect 276326 493398 276562 493634
rect 276646 493398 276882 493634
rect 276326 457718 276562 457954
rect 276646 457718 276882 457954
rect 276326 457398 276562 457634
rect 276646 457398 276882 457634
rect 276326 421718 276562 421954
rect 276646 421718 276882 421954
rect 276326 421398 276562 421634
rect 276646 421398 276882 421634
rect 276326 385718 276562 385954
rect 276646 385718 276882 385954
rect 276326 385398 276562 385634
rect 276646 385398 276882 385634
rect 276326 349718 276562 349954
rect 276646 349718 276882 349954
rect 276326 349398 276562 349634
rect 276646 349398 276882 349634
rect 276326 313718 276562 313954
rect 276646 313718 276882 313954
rect 276326 313398 276562 313634
rect 276646 313398 276882 313634
rect 276326 277718 276562 277954
rect 276646 277718 276882 277954
rect 276326 277398 276562 277634
rect 276646 277398 276882 277634
rect 276326 241718 276562 241954
rect 276646 241718 276882 241954
rect 276326 241398 276562 241634
rect 276646 241398 276882 241634
rect 276326 205718 276562 205954
rect 276646 205718 276882 205954
rect 276326 205398 276562 205634
rect 276646 205398 276882 205634
rect 276326 169718 276562 169954
rect 276646 169718 276882 169954
rect 276326 169398 276562 169634
rect 276646 169398 276882 169634
rect 276326 133718 276562 133954
rect 276646 133718 276882 133954
rect 276326 133398 276562 133634
rect 276646 133398 276882 133634
rect 276326 97718 276562 97954
rect 276646 97718 276882 97954
rect 276326 97398 276562 97634
rect 276646 97398 276882 97634
rect 276326 61718 276562 61954
rect 276646 61718 276882 61954
rect 276326 61398 276562 61634
rect 276646 61398 276882 61634
rect 276326 25718 276562 25954
rect 276646 25718 276882 25954
rect 276326 25398 276562 25634
rect 276646 25398 276882 25634
rect 276326 -5382 276562 -5146
rect 276646 -5382 276882 -5146
rect 276326 -5702 276562 -5466
rect 276646 -5702 276882 -5466
rect 280826 710362 281062 710598
rect 281146 710362 281382 710598
rect 280826 710042 281062 710278
rect 281146 710042 281382 710278
rect 280826 678218 281062 678454
rect 281146 678218 281382 678454
rect 280826 677898 281062 678134
rect 281146 677898 281382 678134
rect 280826 642218 281062 642454
rect 281146 642218 281382 642454
rect 280826 641898 281062 642134
rect 281146 641898 281382 642134
rect 280826 606218 281062 606454
rect 281146 606218 281382 606454
rect 280826 605898 281062 606134
rect 281146 605898 281382 606134
rect 280826 570218 281062 570454
rect 281146 570218 281382 570454
rect 280826 569898 281062 570134
rect 281146 569898 281382 570134
rect 280826 534218 281062 534454
rect 281146 534218 281382 534454
rect 280826 533898 281062 534134
rect 281146 533898 281382 534134
rect 280826 498218 281062 498454
rect 281146 498218 281382 498454
rect 280826 497898 281062 498134
rect 281146 497898 281382 498134
rect 280826 462218 281062 462454
rect 281146 462218 281382 462454
rect 280826 461898 281062 462134
rect 281146 461898 281382 462134
rect 280826 426218 281062 426454
rect 281146 426218 281382 426454
rect 280826 425898 281062 426134
rect 281146 425898 281382 426134
rect 280826 390218 281062 390454
rect 281146 390218 281382 390454
rect 280826 389898 281062 390134
rect 281146 389898 281382 390134
rect 280826 354218 281062 354454
rect 281146 354218 281382 354454
rect 280826 353898 281062 354134
rect 281146 353898 281382 354134
rect 280826 318218 281062 318454
rect 281146 318218 281382 318454
rect 280826 317898 281062 318134
rect 281146 317898 281382 318134
rect 280826 282218 281062 282454
rect 281146 282218 281382 282454
rect 280826 281898 281062 282134
rect 281146 281898 281382 282134
rect 280826 246218 281062 246454
rect 281146 246218 281382 246454
rect 280826 245898 281062 246134
rect 281146 245898 281382 246134
rect 280826 210218 281062 210454
rect 281146 210218 281382 210454
rect 280826 209898 281062 210134
rect 281146 209898 281382 210134
rect 280826 174218 281062 174454
rect 281146 174218 281382 174454
rect 280826 173898 281062 174134
rect 281146 173898 281382 174134
rect 280826 138218 281062 138454
rect 281146 138218 281382 138454
rect 280826 137898 281062 138134
rect 281146 137898 281382 138134
rect 280826 102218 281062 102454
rect 281146 102218 281382 102454
rect 280826 101898 281062 102134
rect 281146 101898 281382 102134
rect 280826 66218 281062 66454
rect 281146 66218 281382 66454
rect 280826 65898 281062 66134
rect 281146 65898 281382 66134
rect 280826 30218 281062 30454
rect 281146 30218 281382 30454
rect 280826 29898 281062 30134
rect 281146 29898 281382 30134
rect 280826 -6342 281062 -6106
rect 281146 -6342 281382 -6106
rect 280826 -6662 281062 -6426
rect 281146 -6662 281382 -6426
rect 285326 711322 285562 711558
rect 285646 711322 285882 711558
rect 285326 711002 285562 711238
rect 285646 711002 285882 711238
rect 285326 682718 285562 682954
rect 285646 682718 285882 682954
rect 285326 682398 285562 682634
rect 285646 682398 285882 682634
rect 285326 646718 285562 646954
rect 285646 646718 285882 646954
rect 285326 646398 285562 646634
rect 285646 646398 285882 646634
rect 285326 610718 285562 610954
rect 285646 610718 285882 610954
rect 285326 610398 285562 610634
rect 285646 610398 285882 610634
rect 285326 574718 285562 574954
rect 285646 574718 285882 574954
rect 285326 574398 285562 574634
rect 285646 574398 285882 574634
rect 285326 538718 285562 538954
rect 285646 538718 285882 538954
rect 285326 538398 285562 538634
rect 285646 538398 285882 538634
rect 285326 502718 285562 502954
rect 285646 502718 285882 502954
rect 285326 502398 285562 502634
rect 285646 502398 285882 502634
rect 285326 466718 285562 466954
rect 285646 466718 285882 466954
rect 285326 466398 285562 466634
rect 285646 466398 285882 466634
rect 285326 430718 285562 430954
rect 285646 430718 285882 430954
rect 285326 430398 285562 430634
rect 285646 430398 285882 430634
rect 285326 394718 285562 394954
rect 285646 394718 285882 394954
rect 285326 394398 285562 394634
rect 285646 394398 285882 394634
rect 285326 358718 285562 358954
rect 285646 358718 285882 358954
rect 285326 358398 285562 358634
rect 285646 358398 285882 358634
rect 285326 322718 285562 322954
rect 285646 322718 285882 322954
rect 285326 322398 285562 322634
rect 285646 322398 285882 322634
rect 285326 286718 285562 286954
rect 285646 286718 285882 286954
rect 285326 286398 285562 286634
rect 285646 286398 285882 286634
rect 285326 250718 285562 250954
rect 285646 250718 285882 250954
rect 285326 250398 285562 250634
rect 285646 250398 285882 250634
rect 285326 214718 285562 214954
rect 285646 214718 285882 214954
rect 285326 214398 285562 214634
rect 285646 214398 285882 214634
rect 285326 178718 285562 178954
rect 285646 178718 285882 178954
rect 285326 178398 285562 178634
rect 285646 178398 285882 178634
rect 285326 142718 285562 142954
rect 285646 142718 285882 142954
rect 285326 142398 285562 142634
rect 285646 142398 285882 142634
rect 285326 106718 285562 106954
rect 285646 106718 285882 106954
rect 285326 106398 285562 106634
rect 285646 106398 285882 106634
rect 285326 70718 285562 70954
rect 285646 70718 285882 70954
rect 285326 70398 285562 70634
rect 285646 70398 285882 70634
rect 285326 34718 285562 34954
rect 285646 34718 285882 34954
rect 285326 34398 285562 34634
rect 285646 34398 285882 34634
rect 285326 -7302 285562 -7066
rect 285646 -7302 285882 -7066
rect 285326 -7622 285562 -7386
rect 285646 -7622 285882 -7386
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 294326 705562 294562 705798
rect 294646 705562 294882 705798
rect 294326 705242 294562 705478
rect 294646 705242 294882 705478
rect 294326 691718 294562 691954
rect 294646 691718 294882 691954
rect 294326 691398 294562 691634
rect 294646 691398 294882 691634
rect 294326 655718 294562 655954
rect 294646 655718 294882 655954
rect 294326 655398 294562 655634
rect 294646 655398 294882 655634
rect 294326 619718 294562 619954
rect 294646 619718 294882 619954
rect 294326 619398 294562 619634
rect 294646 619398 294882 619634
rect 294326 583718 294562 583954
rect 294646 583718 294882 583954
rect 294326 583398 294562 583634
rect 294646 583398 294882 583634
rect 294326 547718 294562 547954
rect 294646 547718 294882 547954
rect 294326 547398 294562 547634
rect 294646 547398 294882 547634
rect 294326 511718 294562 511954
rect 294646 511718 294882 511954
rect 294326 511398 294562 511634
rect 294646 511398 294882 511634
rect 294326 475718 294562 475954
rect 294646 475718 294882 475954
rect 294326 475398 294562 475634
rect 294646 475398 294882 475634
rect 294326 439718 294562 439954
rect 294646 439718 294882 439954
rect 294326 439398 294562 439634
rect 294646 439398 294882 439634
rect 294326 403718 294562 403954
rect 294646 403718 294882 403954
rect 294326 403398 294562 403634
rect 294646 403398 294882 403634
rect 294326 367718 294562 367954
rect 294646 367718 294882 367954
rect 294326 367398 294562 367634
rect 294646 367398 294882 367634
rect 294326 331718 294562 331954
rect 294646 331718 294882 331954
rect 294326 331398 294562 331634
rect 294646 331398 294882 331634
rect 294326 295718 294562 295954
rect 294646 295718 294882 295954
rect 294326 295398 294562 295634
rect 294646 295398 294882 295634
rect 294326 259718 294562 259954
rect 294646 259718 294882 259954
rect 294326 259398 294562 259634
rect 294646 259398 294882 259634
rect 294326 223718 294562 223954
rect 294646 223718 294882 223954
rect 294326 223398 294562 223634
rect 294646 223398 294882 223634
rect 294326 187718 294562 187954
rect 294646 187718 294882 187954
rect 294326 187398 294562 187634
rect 294646 187398 294882 187634
rect 294326 151718 294562 151954
rect 294646 151718 294882 151954
rect 294326 151398 294562 151634
rect 294646 151398 294882 151634
rect 294326 115718 294562 115954
rect 294646 115718 294882 115954
rect 294326 115398 294562 115634
rect 294646 115398 294882 115634
rect 294326 79718 294562 79954
rect 294646 79718 294882 79954
rect 294326 79398 294562 79634
rect 294646 79398 294882 79634
rect 294326 43718 294562 43954
rect 294646 43718 294882 43954
rect 294326 43398 294562 43634
rect 294646 43398 294882 43634
rect 294326 7718 294562 7954
rect 294646 7718 294882 7954
rect 294326 7398 294562 7634
rect 294646 7398 294882 7634
rect 294326 -1542 294562 -1306
rect 294646 -1542 294882 -1306
rect 294326 -1862 294562 -1626
rect 294646 -1862 294882 -1626
rect 298826 706522 299062 706758
rect 299146 706522 299382 706758
rect 298826 706202 299062 706438
rect 299146 706202 299382 706438
rect 298826 696218 299062 696454
rect 299146 696218 299382 696454
rect 298826 695898 299062 696134
rect 299146 695898 299382 696134
rect 298826 660218 299062 660454
rect 299146 660218 299382 660454
rect 298826 659898 299062 660134
rect 299146 659898 299382 660134
rect 298826 624218 299062 624454
rect 299146 624218 299382 624454
rect 298826 623898 299062 624134
rect 299146 623898 299382 624134
rect 298826 588218 299062 588454
rect 299146 588218 299382 588454
rect 298826 587898 299062 588134
rect 299146 587898 299382 588134
rect 298826 552218 299062 552454
rect 299146 552218 299382 552454
rect 298826 551898 299062 552134
rect 299146 551898 299382 552134
rect 298826 516218 299062 516454
rect 299146 516218 299382 516454
rect 298826 515898 299062 516134
rect 299146 515898 299382 516134
rect 298826 480218 299062 480454
rect 299146 480218 299382 480454
rect 298826 479898 299062 480134
rect 299146 479898 299382 480134
rect 298826 444218 299062 444454
rect 299146 444218 299382 444454
rect 298826 443898 299062 444134
rect 299146 443898 299382 444134
rect 298826 408218 299062 408454
rect 299146 408218 299382 408454
rect 298826 407898 299062 408134
rect 299146 407898 299382 408134
rect 298826 372218 299062 372454
rect 299146 372218 299382 372454
rect 298826 371898 299062 372134
rect 299146 371898 299382 372134
rect 298826 336218 299062 336454
rect 299146 336218 299382 336454
rect 298826 335898 299062 336134
rect 299146 335898 299382 336134
rect 298826 300218 299062 300454
rect 299146 300218 299382 300454
rect 298826 299898 299062 300134
rect 299146 299898 299382 300134
rect 298826 264218 299062 264454
rect 299146 264218 299382 264454
rect 298826 263898 299062 264134
rect 299146 263898 299382 264134
rect 298826 228218 299062 228454
rect 299146 228218 299382 228454
rect 298826 227898 299062 228134
rect 299146 227898 299382 228134
rect 298826 192218 299062 192454
rect 299146 192218 299382 192454
rect 298826 191898 299062 192134
rect 299146 191898 299382 192134
rect 298826 156218 299062 156454
rect 299146 156218 299382 156454
rect 298826 155898 299062 156134
rect 299146 155898 299382 156134
rect 298826 120218 299062 120454
rect 299146 120218 299382 120454
rect 298826 119898 299062 120134
rect 299146 119898 299382 120134
rect 298826 84218 299062 84454
rect 299146 84218 299382 84454
rect 298826 83898 299062 84134
rect 299146 83898 299382 84134
rect 298826 48218 299062 48454
rect 299146 48218 299382 48454
rect 298826 47898 299062 48134
rect 299146 47898 299382 48134
rect 298826 12218 299062 12454
rect 299146 12218 299382 12454
rect 298826 11898 299062 12134
rect 299146 11898 299382 12134
rect 298826 -2502 299062 -2266
rect 299146 -2502 299382 -2266
rect 298826 -2822 299062 -2586
rect 299146 -2822 299382 -2586
rect 303326 707482 303562 707718
rect 303646 707482 303882 707718
rect 303326 707162 303562 707398
rect 303646 707162 303882 707398
rect 303326 700718 303562 700954
rect 303646 700718 303882 700954
rect 303326 700398 303562 700634
rect 303646 700398 303882 700634
rect 303326 664718 303562 664954
rect 303646 664718 303882 664954
rect 303326 664398 303562 664634
rect 303646 664398 303882 664634
rect 303326 628718 303562 628954
rect 303646 628718 303882 628954
rect 303326 628398 303562 628634
rect 303646 628398 303882 628634
rect 303326 592718 303562 592954
rect 303646 592718 303882 592954
rect 303326 592398 303562 592634
rect 303646 592398 303882 592634
rect 303326 556718 303562 556954
rect 303646 556718 303882 556954
rect 303326 556398 303562 556634
rect 303646 556398 303882 556634
rect 303326 520718 303562 520954
rect 303646 520718 303882 520954
rect 303326 520398 303562 520634
rect 303646 520398 303882 520634
rect 303326 484718 303562 484954
rect 303646 484718 303882 484954
rect 303326 484398 303562 484634
rect 303646 484398 303882 484634
rect 303326 448718 303562 448954
rect 303646 448718 303882 448954
rect 303326 448398 303562 448634
rect 303646 448398 303882 448634
rect 303326 412718 303562 412954
rect 303646 412718 303882 412954
rect 303326 412398 303562 412634
rect 303646 412398 303882 412634
rect 303326 376718 303562 376954
rect 303646 376718 303882 376954
rect 303326 376398 303562 376634
rect 303646 376398 303882 376634
rect 303326 340718 303562 340954
rect 303646 340718 303882 340954
rect 303326 340398 303562 340634
rect 303646 340398 303882 340634
rect 303326 304718 303562 304954
rect 303646 304718 303882 304954
rect 303326 304398 303562 304634
rect 303646 304398 303882 304634
rect 303326 268718 303562 268954
rect 303646 268718 303882 268954
rect 303326 268398 303562 268634
rect 303646 268398 303882 268634
rect 303326 232718 303562 232954
rect 303646 232718 303882 232954
rect 303326 232398 303562 232634
rect 303646 232398 303882 232634
rect 303326 196718 303562 196954
rect 303646 196718 303882 196954
rect 303326 196398 303562 196634
rect 303646 196398 303882 196634
rect 303326 160718 303562 160954
rect 303646 160718 303882 160954
rect 303326 160398 303562 160634
rect 303646 160398 303882 160634
rect 303326 124718 303562 124954
rect 303646 124718 303882 124954
rect 303326 124398 303562 124634
rect 303646 124398 303882 124634
rect 303326 88718 303562 88954
rect 303646 88718 303882 88954
rect 303326 88398 303562 88634
rect 303646 88398 303882 88634
rect 303326 52718 303562 52954
rect 303646 52718 303882 52954
rect 303326 52398 303562 52634
rect 303646 52398 303882 52634
rect 303326 16718 303562 16954
rect 303646 16718 303882 16954
rect 303326 16398 303562 16634
rect 303646 16398 303882 16634
rect 303326 -3462 303562 -3226
rect 303646 -3462 303882 -3226
rect 303326 -3782 303562 -3546
rect 303646 -3782 303882 -3546
rect 307826 708442 308062 708678
rect 308146 708442 308382 708678
rect 307826 708122 308062 708358
rect 308146 708122 308382 708358
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -4422 308062 -4186
rect 308146 -4422 308382 -4186
rect 307826 -4742 308062 -4506
rect 308146 -4742 308382 -4506
rect 312326 709402 312562 709638
rect 312646 709402 312882 709638
rect 312326 709082 312562 709318
rect 312646 709082 312882 709318
rect 312326 673718 312562 673954
rect 312646 673718 312882 673954
rect 312326 673398 312562 673634
rect 312646 673398 312882 673634
rect 312326 637718 312562 637954
rect 312646 637718 312882 637954
rect 312326 637398 312562 637634
rect 312646 637398 312882 637634
rect 312326 601718 312562 601954
rect 312646 601718 312882 601954
rect 312326 601398 312562 601634
rect 312646 601398 312882 601634
rect 312326 565718 312562 565954
rect 312646 565718 312882 565954
rect 312326 565398 312562 565634
rect 312646 565398 312882 565634
rect 312326 529718 312562 529954
rect 312646 529718 312882 529954
rect 312326 529398 312562 529634
rect 312646 529398 312882 529634
rect 312326 493718 312562 493954
rect 312646 493718 312882 493954
rect 312326 493398 312562 493634
rect 312646 493398 312882 493634
rect 312326 457718 312562 457954
rect 312646 457718 312882 457954
rect 312326 457398 312562 457634
rect 312646 457398 312882 457634
rect 312326 421718 312562 421954
rect 312646 421718 312882 421954
rect 312326 421398 312562 421634
rect 312646 421398 312882 421634
rect 312326 385718 312562 385954
rect 312646 385718 312882 385954
rect 312326 385398 312562 385634
rect 312646 385398 312882 385634
rect 312326 349718 312562 349954
rect 312646 349718 312882 349954
rect 312326 349398 312562 349634
rect 312646 349398 312882 349634
rect 312326 313718 312562 313954
rect 312646 313718 312882 313954
rect 312326 313398 312562 313634
rect 312646 313398 312882 313634
rect 312326 277718 312562 277954
rect 312646 277718 312882 277954
rect 312326 277398 312562 277634
rect 312646 277398 312882 277634
rect 312326 241718 312562 241954
rect 312646 241718 312882 241954
rect 312326 241398 312562 241634
rect 312646 241398 312882 241634
rect 312326 205718 312562 205954
rect 312646 205718 312882 205954
rect 312326 205398 312562 205634
rect 312646 205398 312882 205634
rect 312326 169718 312562 169954
rect 312646 169718 312882 169954
rect 312326 169398 312562 169634
rect 312646 169398 312882 169634
rect 312326 133718 312562 133954
rect 312646 133718 312882 133954
rect 312326 133398 312562 133634
rect 312646 133398 312882 133634
rect 312326 97718 312562 97954
rect 312646 97718 312882 97954
rect 312326 97398 312562 97634
rect 312646 97398 312882 97634
rect 312326 61718 312562 61954
rect 312646 61718 312882 61954
rect 312326 61398 312562 61634
rect 312646 61398 312882 61634
rect 312326 25718 312562 25954
rect 312646 25718 312882 25954
rect 312326 25398 312562 25634
rect 312646 25398 312882 25634
rect 312326 -5382 312562 -5146
rect 312646 -5382 312882 -5146
rect 312326 -5702 312562 -5466
rect 312646 -5702 312882 -5466
rect 316826 710362 317062 710598
rect 317146 710362 317382 710598
rect 316826 710042 317062 710278
rect 317146 710042 317382 710278
rect 316826 678218 317062 678454
rect 317146 678218 317382 678454
rect 316826 677898 317062 678134
rect 317146 677898 317382 678134
rect 316826 642218 317062 642454
rect 317146 642218 317382 642454
rect 316826 641898 317062 642134
rect 317146 641898 317382 642134
rect 316826 606218 317062 606454
rect 317146 606218 317382 606454
rect 316826 605898 317062 606134
rect 317146 605898 317382 606134
rect 316826 570218 317062 570454
rect 317146 570218 317382 570454
rect 316826 569898 317062 570134
rect 317146 569898 317382 570134
rect 316826 534218 317062 534454
rect 317146 534218 317382 534454
rect 316826 533898 317062 534134
rect 317146 533898 317382 534134
rect 316826 498218 317062 498454
rect 317146 498218 317382 498454
rect 316826 497898 317062 498134
rect 317146 497898 317382 498134
rect 316826 462218 317062 462454
rect 317146 462218 317382 462454
rect 316826 461898 317062 462134
rect 317146 461898 317382 462134
rect 316826 426218 317062 426454
rect 317146 426218 317382 426454
rect 316826 425898 317062 426134
rect 317146 425898 317382 426134
rect 316826 390218 317062 390454
rect 317146 390218 317382 390454
rect 316826 389898 317062 390134
rect 317146 389898 317382 390134
rect 316826 354218 317062 354454
rect 317146 354218 317382 354454
rect 316826 353898 317062 354134
rect 317146 353898 317382 354134
rect 316826 318218 317062 318454
rect 317146 318218 317382 318454
rect 316826 317898 317062 318134
rect 317146 317898 317382 318134
rect 316826 282218 317062 282454
rect 317146 282218 317382 282454
rect 316826 281898 317062 282134
rect 317146 281898 317382 282134
rect 316826 246218 317062 246454
rect 317146 246218 317382 246454
rect 316826 245898 317062 246134
rect 317146 245898 317382 246134
rect 316826 210218 317062 210454
rect 317146 210218 317382 210454
rect 316826 209898 317062 210134
rect 317146 209898 317382 210134
rect 316826 174218 317062 174454
rect 317146 174218 317382 174454
rect 316826 173898 317062 174134
rect 317146 173898 317382 174134
rect 316826 138218 317062 138454
rect 317146 138218 317382 138454
rect 316826 137898 317062 138134
rect 317146 137898 317382 138134
rect 316826 102218 317062 102454
rect 317146 102218 317382 102454
rect 316826 101898 317062 102134
rect 317146 101898 317382 102134
rect 316826 66218 317062 66454
rect 317146 66218 317382 66454
rect 316826 65898 317062 66134
rect 317146 65898 317382 66134
rect 316826 30218 317062 30454
rect 317146 30218 317382 30454
rect 316826 29898 317062 30134
rect 317146 29898 317382 30134
rect 316826 -6342 317062 -6106
rect 317146 -6342 317382 -6106
rect 316826 -6662 317062 -6426
rect 317146 -6662 317382 -6426
rect 321326 711322 321562 711558
rect 321646 711322 321882 711558
rect 321326 711002 321562 711238
rect 321646 711002 321882 711238
rect 321326 682718 321562 682954
rect 321646 682718 321882 682954
rect 321326 682398 321562 682634
rect 321646 682398 321882 682634
rect 321326 646718 321562 646954
rect 321646 646718 321882 646954
rect 321326 646398 321562 646634
rect 321646 646398 321882 646634
rect 321326 610718 321562 610954
rect 321646 610718 321882 610954
rect 321326 610398 321562 610634
rect 321646 610398 321882 610634
rect 321326 574718 321562 574954
rect 321646 574718 321882 574954
rect 321326 574398 321562 574634
rect 321646 574398 321882 574634
rect 321326 538718 321562 538954
rect 321646 538718 321882 538954
rect 321326 538398 321562 538634
rect 321646 538398 321882 538634
rect 321326 502718 321562 502954
rect 321646 502718 321882 502954
rect 321326 502398 321562 502634
rect 321646 502398 321882 502634
rect 321326 466718 321562 466954
rect 321646 466718 321882 466954
rect 321326 466398 321562 466634
rect 321646 466398 321882 466634
rect 321326 430718 321562 430954
rect 321646 430718 321882 430954
rect 321326 430398 321562 430634
rect 321646 430398 321882 430634
rect 321326 394718 321562 394954
rect 321646 394718 321882 394954
rect 321326 394398 321562 394634
rect 321646 394398 321882 394634
rect 321326 358718 321562 358954
rect 321646 358718 321882 358954
rect 321326 358398 321562 358634
rect 321646 358398 321882 358634
rect 321326 322718 321562 322954
rect 321646 322718 321882 322954
rect 321326 322398 321562 322634
rect 321646 322398 321882 322634
rect 321326 286718 321562 286954
rect 321646 286718 321882 286954
rect 321326 286398 321562 286634
rect 321646 286398 321882 286634
rect 321326 250718 321562 250954
rect 321646 250718 321882 250954
rect 321326 250398 321562 250634
rect 321646 250398 321882 250634
rect 321326 214718 321562 214954
rect 321646 214718 321882 214954
rect 321326 214398 321562 214634
rect 321646 214398 321882 214634
rect 321326 178718 321562 178954
rect 321646 178718 321882 178954
rect 321326 178398 321562 178634
rect 321646 178398 321882 178634
rect 321326 142718 321562 142954
rect 321646 142718 321882 142954
rect 321326 142398 321562 142634
rect 321646 142398 321882 142634
rect 321326 106718 321562 106954
rect 321646 106718 321882 106954
rect 321326 106398 321562 106634
rect 321646 106398 321882 106634
rect 321326 70718 321562 70954
rect 321646 70718 321882 70954
rect 321326 70398 321562 70634
rect 321646 70398 321882 70634
rect 321326 34718 321562 34954
rect 321646 34718 321882 34954
rect 321326 34398 321562 34634
rect 321646 34398 321882 34634
rect 321326 -7302 321562 -7066
rect 321646 -7302 321882 -7066
rect 321326 -7622 321562 -7386
rect 321646 -7622 321882 -7386
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 330326 705562 330562 705798
rect 330646 705562 330882 705798
rect 330326 705242 330562 705478
rect 330646 705242 330882 705478
rect 330326 691718 330562 691954
rect 330646 691718 330882 691954
rect 330326 691398 330562 691634
rect 330646 691398 330882 691634
rect 330326 655718 330562 655954
rect 330646 655718 330882 655954
rect 330326 655398 330562 655634
rect 330646 655398 330882 655634
rect 330326 619718 330562 619954
rect 330646 619718 330882 619954
rect 330326 619398 330562 619634
rect 330646 619398 330882 619634
rect 330326 583718 330562 583954
rect 330646 583718 330882 583954
rect 330326 583398 330562 583634
rect 330646 583398 330882 583634
rect 330326 547718 330562 547954
rect 330646 547718 330882 547954
rect 330326 547398 330562 547634
rect 330646 547398 330882 547634
rect 330326 511718 330562 511954
rect 330646 511718 330882 511954
rect 330326 511398 330562 511634
rect 330646 511398 330882 511634
rect 330326 475718 330562 475954
rect 330646 475718 330882 475954
rect 330326 475398 330562 475634
rect 330646 475398 330882 475634
rect 330326 439718 330562 439954
rect 330646 439718 330882 439954
rect 330326 439398 330562 439634
rect 330646 439398 330882 439634
rect 330326 403718 330562 403954
rect 330646 403718 330882 403954
rect 330326 403398 330562 403634
rect 330646 403398 330882 403634
rect 330326 367718 330562 367954
rect 330646 367718 330882 367954
rect 330326 367398 330562 367634
rect 330646 367398 330882 367634
rect 330326 331718 330562 331954
rect 330646 331718 330882 331954
rect 330326 331398 330562 331634
rect 330646 331398 330882 331634
rect 330326 295718 330562 295954
rect 330646 295718 330882 295954
rect 330326 295398 330562 295634
rect 330646 295398 330882 295634
rect 330326 259718 330562 259954
rect 330646 259718 330882 259954
rect 330326 259398 330562 259634
rect 330646 259398 330882 259634
rect 330326 223718 330562 223954
rect 330646 223718 330882 223954
rect 330326 223398 330562 223634
rect 330646 223398 330882 223634
rect 330326 187718 330562 187954
rect 330646 187718 330882 187954
rect 330326 187398 330562 187634
rect 330646 187398 330882 187634
rect 330326 151718 330562 151954
rect 330646 151718 330882 151954
rect 330326 151398 330562 151634
rect 330646 151398 330882 151634
rect 330326 115718 330562 115954
rect 330646 115718 330882 115954
rect 330326 115398 330562 115634
rect 330646 115398 330882 115634
rect 330326 79718 330562 79954
rect 330646 79718 330882 79954
rect 330326 79398 330562 79634
rect 330646 79398 330882 79634
rect 330326 43718 330562 43954
rect 330646 43718 330882 43954
rect 330326 43398 330562 43634
rect 330646 43398 330882 43634
rect 330326 7718 330562 7954
rect 330646 7718 330882 7954
rect 330326 7398 330562 7634
rect 330646 7398 330882 7634
rect 330326 -1542 330562 -1306
rect 330646 -1542 330882 -1306
rect 330326 -1862 330562 -1626
rect 330646 -1862 330882 -1626
rect 334826 706522 335062 706758
rect 335146 706522 335382 706758
rect 334826 706202 335062 706438
rect 335146 706202 335382 706438
rect 334826 696218 335062 696454
rect 335146 696218 335382 696454
rect 334826 695898 335062 696134
rect 335146 695898 335382 696134
rect 334826 660218 335062 660454
rect 335146 660218 335382 660454
rect 334826 659898 335062 660134
rect 335146 659898 335382 660134
rect 334826 624218 335062 624454
rect 335146 624218 335382 624454
rect 334826 623898 335062 624134
rect 335146 623898 335382 624134
rect 334826 588218 335062 588454
rect 335146 588218 335382 588454
rect 334826 587898 335062 588134
rect 335146 587898 335382 588134
rect 334826 552218 335062 552454
rect 335146 552218 335382 552454
rect 334826 551898 335062 552134
rect 335146 551898 335382 552134
rect 334826 516218 335062 516454
rect 335146 516218 335382 516454
rect 334826 515898 335062 516134
rect 335146 515898 335382 516134
rect 334826 480218 335062 480454
rect 335146 480218 335382 480454
rect 334826 479898 335062 480134
rect 335146 479898 335382 480134
rect 334826 444218 335062 444454
rect 335146 444218 335382 444454
rect 334826 443898 335062 444134
rect 335146 443898 335382 444134
rect 334826 408218 335062 408454
rect 335146 408218 335382 408454
rect 334826 407898 335062 408134
rect 335146 407898 335382 408134
rect 334826 372218 335062 372454
rect 335146 372218 335382 372454
rect 334826 371898 335062 372134
rect 335146 371898 335382 372134
rect 334826 336218 335062 336454
rect 335146 336218 335382 336454
rect 334826 335898 335062 336134
rect 335146 335898 335382 336134
rect 334826 300218 335062 300454
rect 335146 300218 335382 300454
rect 334826 299898 335062 300134
rect 335146 299898 335382 300134
rect 334826 264218 335062 264454
rect 335146 264218 335382 264454
rect 334826 263898 335062 264134
rect 335146 263898 335382 264134
rect 334826 228218 335062 228454
rect 335146 228218 335382 228454
rect 334826 227898 335062 228134
rect 335146 227898 335382 228134
rect 334826 192218 335062 192454
rect 335146 192218 335382 192454
rect 334826 191898 335062 192134
rect 335146 191898 335382 192134
rect 334826 156218 335062 156454
rect 335146 156218 335382 156454
rect 334826 155898 335062 156134
rect 335146 155898 335382 156134
rect 334826 120218 335062 120454
rect 335146 120218 335382 120454
rect 334826 119898 335062 120134
rect 335146 119898 335382 120134
rect 334826 84218 335062 84454
rect 335146 84218 335382 84454
rect 334826 83898 335062 84134
rect 335146 83898 335382 84134
rect 334826 48218 335062 48454
rect 335146 48218 335382 48454
rect 334826 47898 335062 48134
rect 335146 47898 335382 48134
rect 334826 12218 335062 12454
rect 335146 12218 335382 12454
rect 334826 11898 335062 12134
rect 335146 11898 335382 12134
rect 334826 -2502 335062 -2266
rect 335146 -2502 335382 -2266
rect 334826 -2822 335062 -2586
rect 335146 -2822 335382 -2586
rect 339326 707482 339562 707718
rect 339646 707482 339882 707718
rect 339326 707162 339562 707398
rect 339646 707162 339882 707398
rect 339326 700718 339562 700954
rect 339646 700718 339882 700954
rect 339326 700398 339562 700634
rect 339646 700398 339882 700634
rect 339326 664718 339562 664954
rect 339646 664718 339882 664954
rect 339326 664398 339562 664634
rect 339646 664398 339882 664634
rect 339326 628718 339562 628954
rect 339646 628718 339882 628954
rect 339326 628398 339562 628634
rect 339646 628398 339882 628634
rect 339326 592718 339562 592954
rect 339646 592718 339882 592954
rect 339326 592398 339562 592634
rect 339646 592398 339882 592634
rect 339326 556718 339562 556954
rect 339646 556718 339882 556954
rect 339326 556398 339562 556634
rect 339646 556398 339882 556634
rect 339326 520718 339562 520954
rect 339646 520718 339882 520954
rect 339326 520398 339562 520634
rect 339646 520398 339882 520634
rect 339326 484718 339562 484954
rect 339646 484718 339882 484954
rect 339326 484398 339562 484634
rect 339646 484398 339882 484634
rect 339326 448718 339562 448954
rect 339646 448718 339882 448954
rect 339326 448398 339562 448634
rect 339646 448398 339882 448634
rect 339326 412718 339562 412954
rect 339646 412718 339882 412954
rect 339326 412398 339562 412634
rect 339646 412398 339882 412634
rect 339326 376718 339562 376954
rect 339646 376718 339882 376954
rect 339326 376398 339562 376634
rect 339646 376398 339882 376634
rect 339326 340718 339562 340954
rect 339646 340718 339882 340954
rect 339326 340398 339562 340634
rect 339646 340398 339882 340634
rect 339326 304718 339562 304954
rect 339646 304718 339882 304954
rect 339326 304398 339562 304634
rect 339646 304398 339882 304634
rect 339326 268718 339562 268954
rect 339646 268718 339882 268954
rect 339326 268398 339562 268634
rect 339646 268398 339882 268634
rect 339326 232718 339562 232954
rect 339646 232718 339882 232954
rect 339326 232398 339562 232634
rect 339646 232398 339882 232634
rect 339326 196718 339562 196954
rect 339646 196718 339882 196954
rect 339326 196398 339562 196634
rect 339646 196398 339882 196634
rect 339326 160718 339562 160954
rect 339646 160718 339882 160954
rect 339326 160398 339562 160634
rect 339646 160398 339882 160634
rect 339326 124718 339562 124954
rect 339646 124718 339882 124954
rect 339326 124398 339562 124634
rect 339646 124398 339882 124634
rect 339326 88718 339562 88954
rect 339646 88718 339882 88954
rect 339326 88398 339562 88634
rect 339646 88398 339882 88634
rect 339326 52718 339562 52954
rect 339646 52718 339882 52954
rect 339326 52398 339562 52634
rect 339646 52398 339882 52634
rect 339326 16718 339562 16954
rect 339646 16718 339882 16954
rect 339326 16398 339562 16634
rect 339646 16398 339882 16634
rect 339326 -3462 339562 -3226
rect 339646 -3462 339882 -3226
rect 339326 -3782 339562 -3546
rect 339646 -3782 339882 -3546
rect 343826 708442 344062 708678
rect 344146 708442 344382 708678
rect 343826 708122 344062 708358
rect 344146 708122 344382 708358
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -4422 344062 -4186
rect 344146 -4422 344382 -4186
rect 343826 -4742 344062 -4506
rect 344146 -4742 344382 -4506
rect 348326 709402 348562 709638
rect 348646 709402 348882 709638
rect 348326 709082 348562 709318
rect 348646 709082 348882 709318
rect 348326 673718 348562 673954
rect 348646 673718 348882 673954
rect 348326 673398 348562 673634
rect 348646 673398 348882 673634
rect 348326 637718 348562 637954
rect 348646 637718 348882 637954
rect 348326 637398 348562 637634
rect 348646 637398 348882 637634
rect 348326 601718 348562 601954
rect 348646 601718 348882 601954
rect 348326 601398 348562 601634
rect 348646 601398 348882 601634
rect 348326 565718 348562 565954
rect 348646 565718 348882 565954
rect 348326 565398 348562 565634
rect 348646 565398 348882 565634
rect 348326 529718 348562 529954
rect 348646 529718 348882 529954
rect 348326 529398 348562 529634
rect 348646 529398 348882 529634
rect 348326 493718 348562 493954
rect 348646 493718 348882 493954
rect 348326 493398 348562 493634
rect 348646 493398 348882 493634
rect 348326 457718 348562 457954
rect 348646 457718 348882 457954
rect 348326 457398 348562 457634
rect 348646 457398 348882 457634
rect 348326 421718 348562 421954
rect 348646 421718 348882 421954
rect 348326 421398 348562 421634
rect 348646 421398 348882 421634
rect 348326 385718 348562 385954
rect 348646 385718 348882 385954
rect 348326 385398 348562 385634
rect 348646 385398 348882 385634
rect 348326 349718 348562 349954
rect 348646 349718 348882 349954
rect 348326 349398 348562 349634
rect 348646 349398 348882 349634
rect 348326 313718 348562 313954
rect 348646 313718 348882 313954
rect 348326 313398 348562 313634
rect 348646 313398 348882 313634
rect 348326 277718 348562 277954
rect 348646 277718 348882 277954
rect 348326 277398 348562 277634
rect 348646 277398 348882 277634
rect 348326 241718 348562 241954
rect 348646 241718 348882 241954
rect 348326 241398 348562 241634
rect 348646 241398 348882 241634
rect 348326 205718 348562 205954
rect 348646 205718 348882 205954
rect 348326 205398 348562 205634
rect 348646 205398 348882 205634
rect 348326 169718 348562 169954
rect 348646 169718 348882 169954
rect 348326 169398 348562 169634
rect 348646 169398 348882 169634
rect 348326 133718 348562 133954
rect 348646 133718 348882 133954
rect 348326 133398 348562 133634
rect 348646 133398 348882 133634
rect 348326 97718 348562 97954
rect 348646 97718 348882 97954
rect 348326 97398 348562 97634
rect 348646 97398 348882 97634
rect 348326 61718 348562 61954
rect 348646 61718 348882 61954
rect 348326 61398 348562 61634
rect 348646 61398 348882 61634
rect 348326 25718 348562 25954
rect 348646 25718 348882 25954
rect 348326 25398 348562 25634
rect 348646 25398 348882 25634
rect 348326 -5382 348562 -5146
rect 348646 -5382 348882 -5146
rect 348326 -5702 348562 -5466
rect 348646 -5702 348882 -5466
rect 352826 710362 353062 710598
rect 353146 710362 353382 710598
rect 352826 710042 353062 710278
rect 353146 710042 353382 710278
rect 352826 678218 353062 678454
rect 353146 678218 353382 678454
rect 352826 677898 353062 678134
rect 353146 677898 353382 678134
rect 352826 642218 353062 642454
rect 353146 642218 353382 642454
rect 352826 641898 353062 642134
rect 353146 641898 353382 642134
rect 352826 606218 353062 606454
rect 353146 606218 353382 606454
rect 352826 605898 353062 606134
rect 353146 605898 353382 606134
rect 352826 570218 353062 570454
rect 353146 570218 353382 570454
rect 352826 569898 353062 570134
rect 353146 569898 353382 570134
rect 352826 534218 353062 534454
rect 353146 534218 353382 534454
rect 352826 533898 353062 534134
rect 353146 533898 353382 534134
rect 352826 498218 353062 498454
rect 353146 498218 353382 498454
rect 352826 497898 353062 498134
rect 353146 497898 353382 498134
rect 352826 462218 353062 462454
rect 353146 462218 353382 462454
rect 352826 461898 353062 462134
rect 353146 461898 353382 462134
rect 352826 426218 353062 426454
rect 353146 426218 353382 426454
rect 352826 425898 353062 426134
rect 353146 425898 353382 426134
rect 352826 390218 353062 390454
rect 353146 390218 353382 390454
rect 352826 389898 353062 390134
rect 353146 389898 353382 390134
rect 352826 354218 353062 354454
rect 353146 354218 353382 354454
rect 352826 353898 353062 354134
rect 353146 353898 353382 354134
rect 352826 318218 353062 318454
rect 353146 318218 353382 318454
rect 352826 317898 353062 318134
rect 353146 317898 353382 318134
rect 352826 282218 353062 282454
rect 353146 282218 353382 282454
rect 352826 281898 353062 282134
rect 353146 281898 353382 282134
rect 352826 246218 353062 246454
rect 353146 246218 353382 246454
rect 352826 245898 353062 246134
rect 353146 245898 353382 246134
rect 352826 210218 353062 210454
rect 353146 210218 353382 210454
rect 352826 209898 353062 210134
rect 353146 209898 353382 210134
rect 352826 174218 353062 174454
rect 353146 174218 353382 174454
rect 352826 173898 353062 174134
rect 353146 173898 353382 174134
rect 352826 138218 353062 138454
rect 353146 138218 353382 138454
rect 352826 137898 353062 138134
rect 353146 137898 353382 138134
rect 352826 102218 353062 102454
rect 353146 102218 353382 102454
rect 352826 101898 353062 102134
rect 353146 101898 353382 102134
rect 352826 66218 353062 66454
rect 353146 66218 353382 66454
rect 352826 65898 353062 66134
rect 353146 65898 353382 66134
rect 352826 30218 353062 30454
rect 353146 30218 353382 30454
rect 352826 29898 353062 30134
rect 353146 29898 353382 30134
rect 352826 -6342 353062 -6106
rect 353146 -6342 353382 -6106
rect 352826 -6662 353062 -6426
rect 353146 -6662 353382 -6426
rect 357326 711322 357562 711558
rect 357646 711322 357882 711558
rect 357326 711002 357562 711238
rect 357646 711002 357882 711238
rect 357326 682718 357562 682954
rect 357646 682718 357882 682954
rect 357326 682398 357562 682634
rect 357646 682398 357882 682634
rect 357326 646718 357562 646954
rect 357646 646718 357882 646954
rect 357326 646398 357562 646634
rect 357646 646398 357882 646634
rect 357326 610718 357562 610954
rect 357646 610718 357882 610954
rect 357326 610398 357562 610634
rect 357646 610398 357882 610634
rect 357326 574718 357562 574954
rect 357646 574718 357882 574954
rect 357326 574398 357562 574634
rect 357646 574398 357882 574634
rect 357326 538718 357562 538954
rect 357646 538718 357882 538954
rect 357326 538398 357562 538634
rect 357646 538398 357882 538634
rect 357326 502718 357562 502954
rect 357646 502718 357882 502954
rect 357326 502398 357562 502634
rect 357646 502398 357882 502634
rect 357326 466718 357562 466954
rect 357646 466718 357882 466954
rect 357326 466398 357562 466634
rect 357646 466398 357882 466634
rect 357326 430718 357562 430954
rect 357646 430718 357882 430954
rect 357326 430398 357562 430634
rect 357646 430398 357882 430634
rect 357326 394718 357562 394954
rect 357646 394718 357882 394954
rect 357326 394398 357562 394634
rect 357646 394398 357882 394634
rect 357326 358718 357562 358954
rect 357646 358718 357882 358954
rect 357326 358398 357562 358634
rect 357646 358398 357882 358634
rect 357326 322718 357562 322954
rect 357646 322718 357882 322954
rect 357326 322398 357562 322634
rect 357646 322398 357882 322634
rect 357326 286718 357562 286954
rect 357646 286718 357882 286954
rect 357326 286398 357562 286634
rect 357646 286398 357882 286634
rect 357326 250718 357562 250954
rect 357646 250718 357882 250954
rect 357326 250398 357562 250634
rect 357646 250398 357882 250634
rect 357326 214718 357562 214954
rect 357646 214718 357882 214954
rect 357326 214398 357562 214634
rect 357646 214398 357882 214634
rect 357326 178718 357562 178954
rect 357646 178718 357882 178954
rect 357326 178398 357562 178634
rect 357646 178398 357882 178634
rect 357326 142718 357562 142954
rect 357646 142718 357882 142954
rect 357326 142398 357562 142634
rect 357646 142398 357882 142634
rect 357326 106718 357562 106954
rect 357646 106718 357882 106954
rect 357326 106398 357562 106634
rect 357646 106398 357882 106634
rect 357326 70718 357562 70954
rect 357646 70718 357882 70954
rect 357326 70398 357562 70634
rect 357646 70398 357882 70634
rect 357326 34718 357562 34954
rect 357646 34718 357882 34954
rect 357326 34398 357562 34634
rect 357646 34398 357882 34634
rect 357326 -7302 357562 -7066
rect 357646 -7302 357882 -7066
rect 357326 -7622 357562 -7386
rect 357646 -7622 357882 -7386
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 366326 705562 366562 705798
rect 366646 705562 366882 705798
rect 366326 705242 366562 705478
rect 366646 705242 366882 705478
rect 366326 691718 366562 691954
rect 366646 691718 366882 691954
rect 366326 691398 366562 691634
rect 366646 691398 366882 691634
rect 366326 655718 366562 655954
rect 366646 655718 366882 655954
rect 366326 655398 366562 655634
rect 366646 655398 366882 655634
rect 366326 619718 366562 619954
rect 366646 619718 366882 619954
rect 366326 619398 366562 619634
rect 366646 619398 366882 619634
rect 366326 583718 366562 583954
rect 366646 583718 366882 583954
rect 366326 583398 366562 583634
rect 366646 583398 366882 583634
rect 366326 547718 366562 547954
rect 366646 547718 366882 547954
rect 366326 547398 366562 547634
rect 366646 547398 366882 547634
rect 366326 511718 366562 511954
rect 366646 511718 366882 511954
rect 366326 511398 366562 511634
rect 366646 511398 366882 511634
rect 366326 475718 366562 475954
rect 366646 475718 366882 475954
rect 366326 475398 366562 475634
rect 366646 475398 366882 475634
rect 366326 439718 366562 439954
rect 366646 439718 366882 439954
rect 366326 439398 366562 439634
rect 366646 439398 366882 439634
rect 366326 403718 366562 403954
rect 366646 403718 366882 403954
rect 366326 403398 366562 403634
rect 366646 403398 366882 403634
rect 366326 367718 366562 367954
rect 366646 367718 366882 367954
rect 366326 367398 366562 367634
rect 366646 367398 366882 367634
rect 366326 331718 366562 331954
rect 366646 331718 366882 331954
rect 366326 331398 366562 331634
rect 366646 331398 366882 331634
rect 366326 295718 366562 295954
rect 366646 295718 366882 295954
rect 366326 295398 366562 295634
rect 366646 295398 366882 295634
rect 366326 259718 366562 259954
rect 366646 259718 366882 259954
rect 366326 259398 366562 259634
rect 366646 259398 366882 259634
rect 366326 223718 366562 223954
rect 366646 223718 366882 223954
rect 366326 223398 366562 223634
rect 366646 223398 366882 223634
rect 366326 187718 366562 187954
rect 366646 187718 366882 187954
rect 366326 187398 366562 187634
rect 366646 187398 366882 187634
rect 366326 151718 366562 151954
rect 366646 151718 366882 151954
rect 366326 151398 366562 151634
rect 366646 151398 366882 151634
rect 366326 115718 366562 115954
rect 366646 115718 366882 115954
rect 366326 115398 366562 115634
rect 366646 115398 366882 115634
rect 366326 79718 366562 79954
rect 366646 79718 366882 79954
rect 366326 79398 366562 79634
rect 366646 79398 366882 79634
rect 366326 43718 366562 43954
rect 366646 43718 366882 43954
rect 366326 43398 366562 43634
rect 366646 43398 366882 43634
rect 366326 7718 366562 7954
rect 366646 7718 366882 7954
rect 366326 7398 366562 7634
rect 366646 7398 366882 7634
rect 366326 -1542 366562 -1306
rect 366646 -1542 366882 -1306
rect 366326 -1862 366562 -1626
rect 366646 -1862 366882 -1626
rect 370826 706522 371062 706758
rect 371146 706522 371382 706758
rect 370826 706202 371062 706438
rect 371146 706202 371382 706438
rect 370826 696218 371062 696454
rect 371146 696218 371382 696454
rect 370826 695898 371062 696134
rect 371146 695898 371382 696134
rect 370826 660218 371062 660454
rect 371146 660218 371382 660454
rect 370826 659898 371062 660134
rect 371146 659898 371382 660134
rect 370826 624218 371062 624454
rect 371146 624218 371382 624454
rect 370826 623898 371062 624134
rect 371146 623898 371382 624134
rect 370826 588218 371062 588454
rect 371146 588218 371382 588454
rect 370826 587898 371062 588134
rect 371146 587898 371382 588134
rect 370826 552218 371062 552454
rect 371146 552218 371382 552454
rect 370826 551898 371062 552134
rect 371146 551898 371382 552134
rect 370826 516218 371062 516454
rect 371146 516218 371382 516454
rect 370826 515898 371062 516134
rect 371146 515898 371382 516134
rect 370826 480218 371062 480454
rect 371146 480218 371382 480454
rect 370826 479898 371062 480134
rect 371146 479898 371382 480134
rect 370826 444218 371062 444454
rect 371146 444218 371382 444454
rect 370826 443898 371062 444134
rect 371146 443898 371382 444134
rect 370826 408218 371062 408454
rect 371146 408218 371382 408454
rect 370826 407898 371062 408134
rect 371146 407898 371382 408134
rect 370826 372218 371062 372454
rect 371146 372218 371382 372454
rect 370826 371898 371062 372134
rect 371146 371898 371382 372134
rect 370826 336218 371062 336454
rect 371146 336218 371382 336454
rect 370826 335898 371062 336134
rect 371146 335898 371382 336134
rect 370826 300218 371062 300454
rect 371146 300218 371382 300454
rect 370826 299898 371062 300134
rect 371146 299898 371382 300134
rect 370826 264218 371062 264454
rect 371146 264218 371382 264454
rect 370826 263898 371062 264134
rect 371146 263898 371382 264134
rect 370826 228218 371062 228454
rect 371146 228218 371382 228454
rect 370826 227898 371062 228134
rect 371146 227898 371382 228134
rect 370826 192218 371062 192454
rect 371146 192218 371382 192454
rect 370826 191898 371062 192134
rect 371146 191898 371382 192134
rect 370826 156218 371062 156454
rect 371146 156218 371382 156454
rect 370826 155898 371062 156134
rect 371146 155898 371382 156134
rect 370826 120218 371062 120454
rect 371146 120218 371382 120454
rect 370826 119898 371062 120134
rect 371146 119898 371382 120134
rect 370826 84218 371062 84454
rect 371146 84218 371382 84454
rect 370826 83898 371062 84134
rect 371146 83898 371382 84134
rect 370826 48218 371062 48454
rect 371146 48218 371382 48454
rect 370826 47898 371062 48134
rect 371146 47898 371382 48134
rect 370826 12218 371062 12454
rect 371146 12218 371382 12454
rect 370826 11898 371062 12134
rect 371146 11898 371382 12134
rect 370826 -2502 371062 -2266
rect 371146 -2502 371382 -2266
rect 370826 -2822 371062 -2586
rect 371146 -2822 371382 -2586
rect 375326 707482 375562 707718
rect 375646 707482 375882 707718
rect 375326 707162 375562 707398
rect 375646 707162 375882 707398
rect 375326 700718 375562 700954
rect 375646 700718 375882 700954
rect 375326 700398 375562 700634
rect 375646 700398 375882 700634
rect 375326 664718 375562 664954
rect 375646 664718 375882 664954
rect 375326 664398 375562 664634
rect 375646 664398 375882 664634
rect 375326 628718 375562 628954
rect 375646 628718 375882 628954
rect 375326 628398 375562 628634
rect 375646 628398 375882 628634
rect 375326 592718 375562 592954
rect 375646 592718 375882 592954
rect 375326 592398 375562 592634
rect 375646 592398 375882 592634
rect 375326 556718 375562 556954
rect 375646 556718 375882 556954
rect 375326 556398 375562 556634
rect 375646 556398 375882 556634
rect 375326 520718 375562 520954
rect 375646 520718 375882 520954
rect 375326 520398 375562 520634
rect 375646 520398 375882 520634
rect 375326 484718 375562 484954
rect 375646 484718 375882 484954
rect 375326 484398 375562 484634
rect 375646 484398 375882 484634
rect 375326 448718 375562 448954
rect 375646 448718 375882 448954
rect 375326 448398 375562 448634
rect 375646 448398 375882 448634
rect 375326 412718 375562 412954
rect 375646 412718 375882 412954
rect 375326 412398 375562 412634
rect 375646 412398 375882 412634
rect 375326 376718 375562 376954
rect 375646 376718 375882 376954
rect 375326 376398 375562 376634
rect 375646 376398 375882 376634
rect 375326 340718 375562 340954
rect 375646 340718 375882 340954
rect 375326 340398 375562 340634
rect 375646 340398 375882 340634
rect 375326 304718 375562 304954
rect 375646 304718 375882 304954
rect 375326 304398 375562 304634
rect 375646 304398 375882 304634
rect 375326 268718 375562 268954
rect 375646 268718 375882 268954
rect 375326 268398 375562 268634
rect 375646 268398 375882 268634
rect 375326 232718 375562 232954
rect 375646 232718 375882 232954
rect 375326 232398 375562 232634
rect 375646 232398 375882 232634
rect 375326 196718 375562 196954
rect 375646 196718 375882 196954
rect 375326 196398 375562 196634
rect 375646 196398 375882 196634
rect 375326 160718 375562 160954
rect 375646 160718 375882 160954
rect 375326 160398 375562 160634
rect 375646 160398 375882 160634
rect 375326 124718 375562 124954
rect 375646 124718 375882 124954
rect 375326 124398 375562 124634
rect 375646 124398 375882 124634
rect 375326 88718 375562 88954
rect 375646 88718 375882 88954
rect 375326 88398 375562 88634
rect 375646 88398 375882 88634
rect 375326 52718 375562 52954
rect 375646 52718 375882 52954
rect 375326 52398 375562 52634
rect 375646 52398 375882 52634
rect 375326 16718 375562 16954
rect 375646 16718 375882 16954
rect 375326 16398 375562 16634
rect 375646 16398 375882 16634
rect 375326 -3462 375562 -3226
rect 375646 -3462 375882 -3226
rect 375326 -3782 375562 -3546
rect 375646 -3782 375882 -3546
rect 379826 708442 380062 708678
rect 380146 708442 380382 708678
rect 379826 708122 380062 708358
rect 380146 708122 380382 708358
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -4422 380062 -4186
rect 380146 -4422 380382 -4186
rect 379826 -4742 380062 -4506
rect 380146 -4742 380382 -4506
rect 384326 709402 384562 709638
rect 384646 709402 384882 709638
rect 384326 709082 384562 709318
rect 384646 709082 384882 709318
rect 384326 673718 384562 673954
rect 384646 673718 384882 673954
rect 384326 673398 384562 673634
rect 384646 673398 384882 673634
rect 384326 637718 384562 637954
rect 384646 637718 384882 637954
rect 384326 637398 384562 637634
rect 384646 637398 384882 637634
rect 384326 601718 384562 601954
rect 384646 601718 384882 601954
rect 384326 601398 384562 601634
rect 384646 601398 384882 601634
rect 384326 565718 384562 565954
rect 384646 565718 384882 565954
rect 384326 565398 384562 565634
rect 384646 565398 384882 565634
rect 384326 529718 384562 529954
rect 384646 529718 384882 529954
rect 384326 529398 384562 529634
rect 384646 529398 384882 529634
rect 384326 493718 384562 493954
rect 384646 493718 384882 493954
rect 384326 493398 384562 493634
rect 384646 493398 384882 493634
rect 384326 457718 384562 457954
rect 384646 457718 384882 457954
rect 384326 457398 384562 457634
rect 384646 457398 384882 457634
rect 384326 421718 384562 421954
rect 384646 421718 384882 421954
rect 384326 421398 384562 421634
rect 384646 421398 384882 421634
rect 384326 385718 384562 385954
rect 384646 385718 384882 385954
rect 384326 385398 384562 385634
rect 384646 385398 384882 385634
rect 384326 349718 384562 349954
rect 384646 349718 384882 349954
rect 384326 349398 384562 349634
rect 384646 349398 384882 349634
rect 384326 313718 384562 313954
rect 384646 313718 384882 313954
rect 384326 313398 384562 313634
rect 384646 313398 384882 313634
rect 384326 277718 384562 277954
rect 384646 277718 384882 277954
rect 384326 277398 384562 277634
rect 384646 277398 384882 277634
rect 384326 241718 384562 241954
rect 384646 241718 384882 241954
rect 384326 241398 384562 241634
rect 384646 241398 384882 241634
rect 384326 205718 384562 205954
rect 384646 205718 384882 205954
rect 384326 205398 384562 205634
rect 384646 205398 384882 205634
rect 384326 169718 384562 169954
rect 384646 169718 384882 169954
rect 384326 169398 384562 169634
rect 384646 169398 384882 169634
rect 384326 133718 384562 133954
rect 384646 133718 384882 133954
rect 384326 133398 384562 133634
rect 384646 133398 384882 133634
rect 384326 97718 384562 97954
rect 384646 97718 384882 97954
rect 384326 97398 384562 97634
rect 384646 97398 384882 97634
rect 384326 61718 384562 61954
rect 384646 61718 384882 61954
rect 384326 61398 384562 61634
rect 384646 61398 384882 61634
rect 384326 25718 384562 25954
rect 384646 25718 384882 25954
rect 384326 25398 384562 25634
rect 384646 25398 384882 25634
rect 384326 -5382 384562 -5146
rect 384646 -5382 384882 -5146
rect 384326 -5702 384562 -5466
rect 384646 -5702 384882 -5466
rect 388826 710362 389062 710598
rect 389146 710362 389382 710598
rect 388826 710042 389062 710278
rect 389146 710042 389382 710278
rect 388826 678218 389062 678454
rect 389146 678218 389382 678454
rect 388826 677898 389062 678134
rect 389146 677898 389382 678134
rect 388826 642218 389062 642454
rect 389146 642218 389382 642454
rect 388826 641898 389062 642134
rect 389146 641898 389382 642134
rect 388826 606218 389062 606454
rect 389146 606218 389382 606454
rect 388826 605898 389062 606134
rect 389146 605898 389382 606134
rect 388826 570218 389062 570454
rect 389146 570218 389382 570454
rect 388826 569898 389062 570134
rect 389146 569898 389382 570134
rect 388826 534218 389062 534454
rect 389146 534218 389382 534454
rect 388826 533898 389062 534134
rect 389146 533898 389382 534134
rect 388826 498218 389062 498454
rect 389146 498218 389382 498454
rect 388826 497898 389062 498134
rect 389146 497898 389382 498134
rect 388826 462218 389062 462454
rect 389146 462218 389382 462454
rect 388826 461898 389062 462134
rect 389146 461898 389382 462134
rect 388826 426218 389062 426454
rect 389146 426218 389382 426454
rect 388826 425898 389062 426134
rect 389146 425898 389382 426134
rect 388826 390218 389062 390454
rect 389146 390218 389382 390454
rect 388826 389898 389062 390134
rect 389146 389898 389382 390134
rect 388826 354218 389062 354454
rect 389146 354218 389382 354454
rect 388826 353898 389062 354134
rect 389146 353898 389382 354134
rect 388826 318218 389062 318454
rect 389146 318218 389382 318454
rect 388826 317898 389062 318134
rect 389146 317898 389382 318134
rect 388826 282218 389062 282454
rect 389146 282218 389382 282454
rect 388826 281898 389062 282134
rect 389146 281898 389382 282134
rect 388826 246218 389062 246454
rect 389146 246218 389382 246454
rect 388826 245898 389062 246134
rect 389146 245898 389382 246134
rect 388826 210218 389062 210454
rect 389146 210218 389382 210454
rect 388826 209898 389062 210134
rect 389146 209898 389382 210134
rect 388826 174218 389062 174454
rect 389146 174218 389382 174454
rect 388826 173898 389062 174134
rect 389146 173898 389382 174134
rect 388826 138218 389062 138454
rect 389146 138218 389382 138454
rect 388826 137898 389062 138134
rect 389146 137898 389382 138134
rect 388826 102218 389062 102454
rect 389146 102218 389382 102454
rect 388826 101898 389062 102134
rect 389146 101898 389382 102134
rect 388826 66218 389062 66454
rect 389146 66218 389382 66454
rect 388826 65898 389062 66134
rect 389146 65898 389382 66134
rect 388826 30218 389062 30454
rect 389146 30218 389382 30454
rect 388826 29898 389062 30134
rect 389146 29898 389382 30134
rect 388826 -6342 389062 -6106
rect 389146 -6342 389382 -6106
rect 388826 -6662 389062 -6426
rect 389146 -6662 389382 -6426
rect 393326 711322 393562 711558
rect 393646 711322 393882 711558
rect 393326 711002 393562 711238
rect 393646 711002 393882 711238
rect 393326 682718 393562 682954
rect 393646 682718 393882 682954
rect 393326 682398 393562 682634
rect 393646 682398 393882 682634
rect 393326 646718 393562 646954
rect 393646 646718 393882 646954
rect 393326 646398 393562 646634
rect 393646 646398 393882 646634
rect 393326 610718 393562 610954
rect 393646 610718 393882 610954
rect 393326 610398 393562 610634
rect 393646 610398 393882 610634
rect 393326 574718 393562 574954
rect 393646 574718 393882 574954
rect 393326 574398 393562 574634
rect 393646 574398 393882 574634
rect 393326 538718 393562 538954
rect 393646 538718 393882 538954
rect 393326 538398 393562 538634
rect 393646 538398 393882 538634
rect 393326 502718 393562 502954
rect 393646 502718 393882 502954
rect 393326 502398 393562 502634
rect 393646 502398 393882 502634
rect 393326 466718 393562 466954
rect 393646 466718 393882 466954
rect 393326 466398 393562 466634
rect 393646 466398 393882 466634
rect 393326 430718 393562 430954
rect 393646 430718 393882 430954
rect 393326 430398 393562 430634
rect 393646 430398 393882 430634
rect 393326 394718 393562 394954
rect 393646 394718 393882 394954
rect 393326 394398 393562 394634
rect 393646 394398 393882 394634
rect 393326 358718 393562 358954
rect 393646 358718 393882 358954
rect 393326 358398 393562 358634
rect 393646 358398 393882 358634
rect 393326 322718 393562 322954
rect 393646 322718 393882 322954
rect 393326 322398 393562 322634
rect 393646 322398 393882 322634
rect 393326 286718 393562 286954
rect 393646 286718 393882 286954
rect 393326 286398 393562 286634
rect 393646 286398 393882 286634
rect 393326 250718 393562 250954
rect 393646 250718 393882 250954
rect 393326 250398 393562 250634
rect 393646 250398 393882 250634
rect 393326 214718 393562 214954
rect 393646 214718 393882 214954
rect 393326 214398 393562 214634
rect 393646 214398 393882 214634
rect 393326 178718 393562 178954
rect 393646 178718 393882 178954
rect 393326 178398 393562 178634
rect 393646 178398 393882 178634
rect 393326 142718 393562 142954
rect 393646 142718 393882 142954
rect 393326 142398 393562 142634
rect 393646 142398 393882 142634
rect 393326 106718 393562 106954
rect 393646 106718 393882 106954
rect 393326 106398 393562 106634
rect 393646 106398 393882 106634
rect 393326 70718 393562 70954
rect 393646 70718 393882 70954
rect 393326 70398 393562 70634
rect 393646 70398 393882 70634
rect 393326 34718 393562 34954
rect 393646 34718 393882 34954
rect 393326 34398 393562 34634
rect 393646 34398 393882 34634
rect 393326 -7302 393562 -7066
rect 393646 -7302 393882 -7066
rect 393326 -7622 393562 -7386
rect 393646 -7622 393882 -7386
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 402326 705562 402562 705798
rect 402646 705562 402882 705798
rect 402326 705242 402562 705478
rect 402646 705242 402882 705478
rect 402326 691718 402562 691954
rect 402646 691718 402882 691954
rect 402326 691398 402562 691634
rect 402646 691398 402882 691634
rect 402326 655718 402562 655954
rect 402646 655718 402882 655954
rect 402326 655398 402562 655634
rect 402646 655398 402882 655634
rect 402326 619718 402562 619954
rect 402646 619718 402882 619954
rect 402326 619398 402562 619634
rect 402646 619398 402882 619634
rect 402326 583718 402562 583954
rect 402646 583718 402882 583954
rect 402326 583398 402562 583634
rect 402646 583398 402882 583634
rect 402326 547718 402562 547954
rect 402646 547718 402882 547954
rect 402326 547398 402562 547634
rect 402646 547398 402882 547634
rect 402326 511718 402562 511954
rect 402646 511718 402882 511954
rect 402326 511398 402562 511634
rect 402646 511398 402882 511634
rect 402326 475718 402562 475954
rect 402646 475718 402882 475954
rect 402326 475398 402562 475634
rect 402646 475398 402882 475634
rect 402326 439718 402562 439954
rect 402646 439718 402882 439954
rect 402326 439398 402562 439634
rect 402646 439398 402882 439634
rect 402326 403718 402562 403954
rect 402646 403718 402882 403954
rect 402326 403398 402562 403634
rect 402646 403398 402882 403634
rect 402326 367718 402562 367954
rect 402646 367718 402882 367954
rect 402326 367398 402562 367634
rect 402646 367398 402882 367634
rect 402326 331718 402562 331954
rect 402646 331718 402882 331954
rect 402326 331398 402562 331634
rect 402646 331398 402882 331634
rect 402326 295718 402562 295954
rect 402646 295718 402882 295954
rect 402326 295398 402562 295634
rect 402646 295398 402882 295634
rect 402326 259718 402562 259954
rect 402646 259718 402882 259954
rect 402326 259398 402562 259634
rect 402646 259398 402882 259634
rect 402326 223718 402562 223954
rect 402646 223718 402882 223954
rect 402326 223398 402562 223634
rect 402646 223398 402882 223634
rect 402326 187718 402562 187954
rect 402646 187718 402882 187954
rect 402326 187398 402562 187634
rect 402646 187398 402882 187634
rect 402326 151718 402562 151954
rect 402646 151718 402882 151954
rect 402326 151398 402562 151634
rect 402646 151398 402882 151634
rect 402326 115718 402562 115954
rect 402646 115718 402882 115954
rect 402326 115398 402562 115634
rect 402646 115398 402882 115634
rect 402326 79718 402562 79954
rect 402646 79718 402882 79954
rect 402326 79398 402562 79634
rect 402646 79398 402882 79634
rect 402326 43718 402562 43954
rect 402646 43718 402882 43954
rect 402326 43398 402562 43634
rect 402646 43398 402882 43634
rect 402326 7718 402562 7954
rect 402646 7718 402882 7954
rect 402326 7398 402562 7634
rect 402646 7398 402882 7634
rect 402326 -1542 402562 -1306
rect 402646 -1542 402882 -1306
rect 402326 -1862 402562 -1626
rect 402646 -1862 402882 -1626
rect 406826 706522 407062 706758
rect 407146 706522 407382 706758
rect 406826 706202 407062 706438
rect 407146 706202 407382 706438
rect 406826 696218 407062 696454
rect 407146 696218 407382 696454
rect 406826 695898 407062 696134
rect 407146 695898 407382 696134
rect 406826 660218 407062 660454
rect 407146 660218 407382 660454
rect 406826 659898 407062 660134
rect 407146 659898 407382 660134
rect 406826 624218 407062 624454
rect 407146 624218 407382 624454
rect 406826 623898 407062 624134
rect 407146 623898 407382 624134
rect 406826 588218 407062 588454
rect 407146 588218 407382 588454
rect 406826 587898 407062 588134
rect 407146 587898 407382 588134
rect 406826 552218 407062 552454
rect 407146 552218 407382 552454
rect 406826 551898 407062 552134
rect 407146 551898 407382 552134
rect 406826 516218 407062 516454
rect 407146 516218 407382 516454
rect 406826 515898 407062 516134
rect 407146 515898 407382 516134
rect 406826 480218 407062 480454
rect 407146 480218 407382 480454
rect 406826 479898 407062 480134
rect 407146 479898 407382 480134
rect 406826 444218 407062 444454
rect 407146 444218 407382 444454
rect 406826 443898 407062 444134
rect 407146 443898 407382 444134
rect 406826 408218 407062 408454
rect 407146 408218 407382 408454
rect 406826 407898 407062 408134
rect 407146 407898 407382 408134
rect 406826 372218 407062 372454
rect 407146 372218 407382 372454
rect 406826 371898 407062 372134
rect 407146 371898 407382 372134
rect 406826 336218 407062 336454
rect 407146 336218 407382 336454
rect 406826 335898 407062 336134
rect 407146 335898 407382 336134
rect 406826 300218 407062 300454
rect 407146 300218 407382 300454
rect 406826 299898 407062 300134
rect 407146 299898 407382 300134
rect 406826 264218 407062 264454
rect 407146 264218 407382 264454
rect 406826 263898 407062 264134
rect 407146 263898 407382 264134
rect 406826 228218 407062 228454
rect 407146 228218 407382 228454
rect 406826 227898 407062 228134
rect 407146 227898 407382 228134
rect 406826 192218 407062 192454
rect 407146 192218 407382 192454
rect 406826 191898 407062 192134
rect 407146 191898 407382 192134
rect 406826 156218 407062 156454
rect 407146 156218 407382 156454
rect 406826 155898 407062 156134
rect 407146 155898 407382 156134
rect 406826 120218 407062 120454
rect 407146 120218 407382 120454
rect 406826 119898 407062 120134
rect 407146 119898 407382 120134
rect 406826 84218 407062 84454
rect 407146 84218 407382 84454
rect 406826 83898 407062 84134
rect 407146 83898 407382 84134
rect 406826 48218 407062 48454
rect 407146 48218 407382 48454
rect 406826 47898 407062 48134
rect 407146 47898 407382 48134
rect 406826 12218 407062 12454
rect 407146 12218 407382 12454
rect 406826 11898 407062 12134
rect 407146 11898 407382 12134
rect 406826 -2502 407062 -2266
rect 407146 -2502 407382 -2266
rect 406826 -2822 407062 -2586
rect 407146 -2822 407382 -2586
rect 411326 707482 411562 707718
rect 411646 707482 411882 707718
rect 411326 707162 411562 707398
rect 411646 707162 411882 707398
rect 411326 700718 411562 700954
rect 411646 700718 411882 700954
rect 411326 700398 411562 700634
rect 411646 700398 411882 700634
rect 411326 664718 411562 664954
rect 411646 664718 411882 664954
rect 411326 664398 411562 664634
rect 411646 664398 411882 664634
rect 411326 628718 411562 628954
rect 411646 628718 411882 628954
rect 411326 628398 411562 628634
rect 411646 628398 411882 628634
rect 411326 592718 411562 592954
rect 411646 592718 411882 592954
rect 411326 592398 411562 592634
rect 411646 592398 411882 592634
rect 411326 556718 411562 556954
rect 411646 556718 411882 556954
rect 411326 556398 411562 556634
rect 411646 556398 411882 556634
rect 411326 520718 411562 520954
rect 411646 520718 411882 520954
rect 411326 520398 411562 520634
rect 411646 520398 411882 520634
rect 411326 484718 411562 484954
rect 411646 484718 411882 484954
rect 411326 484398 411562 484634
rect 411646 484398 411882 484634
rect 411326 448718 411562 448954
rect 411646 448718 411882 448954
rect 411326 448398 411562 448634
rect 411646 448398 411882 448634
rect 411326 412718 411562 412954
rect 411646 412718 411882 412954
rect 411326 412398 411562 412634
rect 411646 412398 411882 412634
rect 411326 376718 411562 376954
rect 411646 376718 411882 376954
rect 411326 376398 411562 376634
rect 411646 376398 411882 376634
rect 411326 340718 411562 340954
rect 411646 340718 411882 340954
rect 411326 340398 411562 340634
rect 411646 340398 411882 340634
rect 411326 304718 411562 304954
rect 411646 304718 411882 304954
rect 411326 304398 411562 304634
rect 411646 304398 411882 304634
rect 411326 268718 411562 268954
rect 411646 268718 411882 268954
rect 411326 268398 411562 268634
rect 411646 268398 411882 268634
rect 411326 232718 411562 232954
rect 411646 232718 411882 232954
rect 411326 232398 411562 232634
rect 411646 232398 411882 232634
rect 411326 196718 411562 196954
rect 411646 196718 411882 196954
rect 411326 196398 411562 196634
rect 411646 196398 411882 196634
rect 411326 160718 411562 160954
rect 411646 160718 411882 160954
rect 411326 160398 411562 160634
rect 411646 160398 411882 160634
rect 411326 124718 411562 124954
rect 411646 124718 411882 124954
rect 411326 124398 411562 124634
rect 411646 124398 411882 124634
rect 411326 88718 411562 88954
rect 411646 88718 411882 88954
rect 411326 88398 411562 88634
rect 411646 88398 411882 88634
rect 411326 52718 411562 52954
rect 411646 52718 411882 52954
rect 411326 52398 411562 52634
rect 411646 52398 411882 52634
rect 411326 16718 411562 16954
rect 411646 16718 411882 16954
rect 411326 16398 411562 16634
rect 411646 16398 411882 16634
rect 411326 -3462 411562 -3226
rect 411646 -3462 411882 -3226
rect 411326 -3782 411562 -3546
rect 411646 -3782 411882 -3546
rect 415826 708442 416062 708678
rect 416146 708442 416382 708678
rect 415826 708122 416062 708358
rect 416146 708122 416382 708358
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -4422 416062 -4186
rect 416146 -4422 416382 -4186
rect 415826 -4742 416062 -4506
rect 416146 -4742 416382 -4506
rect 420326 709402 420562 709638
rect 420646 709402 420882 709638
rect 420326 709082 420562 709318
rect 420646 709082 420882 709318
rect 420326 673718 420562 673954
rect 420646 673718 420882 673954
rect 420326 673398 420562 673634
rect 420646 673398 420882 673634
rect 420326 637718 420562 637954
rect 420646 637718 420882 637954
rect 420326 637398 420562 637634
rect 420646 637398 420882 637634
rect 420326 601718 420562 601954
rect 420646 601718 420882 601954
rect 420326 601398 420562 601634
rect 420646 601398 420882 601634
rect 420326 565718 420562 565954
rect 420646 565718 420882 565954
rect 420326 565398 420562 565634
rect 420646 565398 420882 565634
rect 420326 529718 420562 529954
rect 420646 529718 420882 529954
rect 420326 529398 420562 529634
rect 420646 529398 420882 529634
rect 420326 493718 420562 493954
rect 420646 493718 420882 493954
rect 420326 493398 420562 493634
rect 420646 493398 420882 493634
rect 420326 457718 420562 457954
rect 420646 457718 420882 457954
rect 420326 457398 420562 457634
rect 420646 457398 420882 457634
rect 420326 421718 420562 421954
rect 420646 421718 420882 421954
rect 420326 421398 420562 421634
rect 420646 421398 420882 421634
rect 420326 385718 420562 385954
rect 420646 385718 420882 385954
rect 420326 385398 420562 385634
rect 420646 385398 420882 385634
rect 420326 349718 420562 349954
rect 420646 349718 420882 349954
rect 420326 349398 420562 349634
rect 420646 349398 420882 349634
rect 420326 313718 420562 313954
rect 420646 313718 420882 313954
rect 420326 313398 420562 313634
rect 420646 313398 420882 313634
rect 420326 277718 420562 277954
rect 420646 277718 420882 277954
rect 420326 277398 420562 277634
rect 420646 277398 420882 277634
rect 420326 241718 420562 241954
rect 420646 241718 420882 241954
rect 420326 241398 420562 241634
rect 420646 241398 420882 241634
rect 420326 205718 420562 205954
rect 420646 205718 420882 205954
rect 420326 205398 420562 205634
rect 420646 205398 420882 205634
rect 420326 169718 420562 169954
rect 420646 169718 420882 169954
rect 420326 169398 420562 169634
rect 420646 169398 420882 169634
rect 420326 133718 420562 133954
rect 420646 133718 420882 133954
rect 420326 133398 420562 133634
rect 420646 133398 420882 133634
rect 420326 97718 420562 97954
rect 420646 97718 420882 97954
rect 420326 97398 420562 97634
rect 420646 97398 420882 97634
rect 420326 61718 420562 61954
rect 420646 61718 420882 61954
rect 420326 61398 420562 61634
rect 420646 61398 420882 61634
rect 420326 25718 420562 25954
rect 420646 25718 420882 25954
rect 420326 25398 420562 25634
rect 420646 25398 420882 25634
rect 420326 -5382 420562 -5146
rect 420646 -5382 420882 -5146
rect 420326 -5702 420562 -5466
rect 420646 -5702 420882 -5466
rect 424826 710362 425062 710598
rect 425146 710362 425382 710598
rect 424826 710042 425062 710278
rect 425146 710042 425382 710278
rect 424826 678218 425062 678454
rect 425146 678218 425382 678454
rect 424826 677898 425062 678134
rect 425146 677898 425382 678134
rect 424826 642218 425062 642454
rect 425146 642218 425382 642454
rect 424826 641898 425062 642134
rect 425146 641898 425382 642134
rect 424826 606218 425062 606454
rect 425146 606218 425382 606454
rect 424826 605898 425062 606134
rect 425146 605898 425382 606134
rect 424826 570218 425062 570454
rect 425146 570218 425382 570454
rect 424826 569898 425062 570134
rect 425146 569898 425382 570134
rect 424826 534218 425062 534454
rect 425146 534218 425382 534454
rect 424826 533898 425062 534134
rect 425146 533898 425382 534134
rect 424826 498218 425062 498454
rect 425146 498218 425382 498454
rect 424826 497898 425062 498134
rect 425146 497898 425382 498134
rect 424826 462218 425062 462454
rect 425146 462218 425382 462454
rect 424826 461898 425062 462134
rect 425146 461898 425382 462134
rect 424826 426218 425062 426454
rect 425146 426218 425382 426454
rect 424826 425898 425062 426134
rect 425146 425898 425382 426134
rect 424826 390218 425062 390454
rect 425146 390218 425382 390454
rect 424826 389898 425062 390134
rect 425146 389898 425382 390134
rect 424826 354218 425062 354454
rect 425146 354218 425382 354454
rect 424826 353898 425062 354134
rect 425146 353898 425382 354134
rect 424826 318218 425062 318454
rect 425146 318218 425382 318454
rect 424826 317898 425062 318134
rect 425146 317898 425382 318134
rect 424826 282218 425062 282454
rect 425146 282218 425382 282454
rect 424826 281898 425062 282134
rect 425146 281898 425382 282134
rect 424826 246218 425062 246454
rect 425146 246218 425382 246454
rect 424826 245898 425062 246134
rect 425146 245898 425382 246134
rect 424826 210218 425062 210454
rect 425146 210218 425382 210454
rect 424826 209898 425062 210134
rect 425146 209898 425382 210134
rect 424826 174218 425062 174454
rect 425146 174218 425382 174454
rect 424826 173898 425062 174134
rect 425146 173898 425382 174134
rect 424826 138218 425062 138454
rect 425146 138218 425382 138454
rect 424826 137898 425062 138134
rect 425146 137898 425382 138134
rect 424826 102218 425062 102454
rect 425146 102218 425382 102454
rect 424826 101898 425062 102134
rect 425146 101898 425382 102134
rect 424826 66218 425062 66454
rect 425146 66218 425382 66454
rect 424826 65898 425062 66134
rect 425146 65898 425382 66134
rect 424826 30218 425062 30454
rect 425146 30218 425382 30454
rect 424826 29898 425062 30134
rect 425146 29898 425382 30134
rect 424826 -6342 425062 -6106
rect 425146 -6342 425382 -6106
rect 424826 -6662 425062 -6426
rect 425146 -6662 425382 -6426
rect 429326 711322 429562 711558
rect 429646 711322 429882 711558
rect 429326 711002 429562 711238
rect 429646 711002 429882 711238
rect 429326 682718 429562 682954
rect 429646 682718 429882 682954
rect 429326 682398 429562 682634
rect 429646 682398 429882 682634
rect 429326 646718 429562 646954
rect 429646 646718 429882 646954
rect 429326 646398 429562 646634
rect 429646 646398 429882 646634
rect 429326 610718 429562 610954
rect 429646 610718 429882 610954
rect 429326 610398 429562 610634
rect 429646 610398 429882 610634
rect 429326 574718 429562 574954
rect 429646 574718 429882 574954
rect 429326 574398 429562 574634
rect 429646 574398 429882 574634
rect 429326 538718 429562 538954
rect 429646 538718 429882 538954
rect 429326 538398 429562 538634
rect 429646 538398 429882 538634
rect 429326 502718 429562 502954
rect 429646 502718 429882 502954
rect 429326 502398 429562 502634
rect 429646 502398 429882 502634
rect 429326 466718 429562 466954
rect 429646 466718 429882 466954
rect 429326 466398 429562 466634
rect 429646 466398 429882 466634
rect 429326 430718 429562 430954
rect 429646 430718 429882 430954
rect 429326 430398 429562 430634
rect 429646 430398 429882 430634
rect 429326 394718 429562 394954
rect 429646 394718 429882 394954
rect 429326 394398 429562 394634
rect 429646 394398 429882 394634
rect 429326 358718 429562 358954
rect 429646 358718 429882 358954
rect 429326 358398 429562 358634
rect 429646 358398 429882 358634
rect 429326 322718 429562 322954
rect 429646 322718 429882 322954
rect 429326 322398 429562 322634
rect 429646 322398 429882 322634
rect 429326 286718 429562 286954
rect 429646 286718 429882 286954
rect 429326 286398 429562 286634
rect 429646 286398 429882 286634
rect 429326 250718 429562 250954
rect 429646 250718 429882 250954
rect 429326 250398 429562 250634
rect 429646 250398 429882 250634
rect 429326 214718 429562 214954
rect 429646 214718 429882 214954
rect 429326 214398 429562 214634
rect 429646 214398 429882 214634
rect 429326 178718 429562 178954
rect 429646 178718 429882 178954
rect 429326 178398 429562 178634
rect 429646 178398 429882 178634
rect 429326 142718 429562 142954
rect 429646 142718 429882 142954
rect 429326 142398 429562 142634
rect 429646 142398 429882 142634
rect 429326 106718 429562 106954
rect 429646 106718 429882 106954
rect 429326 106398 429562 106634
rect 429646 106398 429882 106634
rect 429326 70718 429562 70954
rect 429646 70718 429882 70954
rect 429326 70398 429562 70634
rect 429646 70398 429882 70634
rect 429326 34718 429562 34954
rect 429646 34718 429882 34954
rect 429326 34398 429562 34634
rect 429646 34398 429882 34634
rect 429326 -7302 429562 -7066
rect 429646 -7302 429882 -7066
rect 429326 -7622 429562 -7386
rect 429646 -7622 429882 -7386
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 438326 705562 438562 705798
rect 438646 705562 438882 705798
rect 438326 705242 438562 705478
rect 438646 705242 438882 705478
rect 438326 691718 438562 691954
rect 438646 691718 438882 691954
rect 438326 691398 438562 691634
rect 438646 691398 438882 691634
rect 438326 655718 438562 655954
rect 438646 655718 438882 655954
rect 438326 655398 438562 655634
rect 438646 655398 438882 655634
rect 438326 619718 438562 619954
rect 438646 619718 438882 619954
rect 438326 619398 438562 619634
rect 438646 619398 438882 619634
rect 438326 583718 438562 583954
rect 438646 583718 438882 583954
rect 438326 583398 438562 583634
rect 438646 583398 438882 583634
rect 438326 547718 438562 547954
rect 438646 547718 438882 547954
rect 438326 547398 438562 547634
rect 438646 547398 438882 547634
rect 438326 511718 438562 511954
rect 438646 511718 438882 511954
rect 438326 511398 438562 511634
rect 438646 511398 438882 511634
rect 438326 475718 438562 475954
rect 438646 475718 438882 475954
rect 438326 475398 438562 475634
rect 438646 475398 438882 475634
rect 438326 439718 438562 439954
rect 438646 439718 438882 439954
rect 438326 439398 438562 439634
rect 438646 439398 438882 439634
rect 438326 403718 438562 403954
rect 438646 403718 438882 403954
rect 438326 403398 438562 403634
rect 438646 403398 438882 403634
rect 438326 367718 438562 367954
rect 438646 367718 438882 367954
rect 438326 367398 438562 367634
rect 438646 367398 438882 367634
rect 438326 331718 438562 331954
rect 438646 331718 438882 331954
rect 438326 331398 438562 331634
rect 438646 331398 438882 331634
rect 438326 295718 438562 295954
rect 438646 295718 438882 295954
rect 438326 295398 438562 295634
rect 438646 295398 438882 295634
rect 438326 259718 438562 259954
rect 438646 259718 438882 259954
rect 438326 259398 438562 259634
rect 438646 259398 438882 259634
rect 438326 223718 438562 223954
rect 438646 223718 438882 223954
rect 438326 223398 438562 223634
rect 438646 223398 438882 223634
rect 438326 187718 438562 187954
rect 438646 187718 438882 187954
rect 438326 187398 438562 187634
rect 438646 187398 438882 187634
rect 438326 151718 438562 151954
rect 438646 151718 438882 151954
rect 438326 151398 438562 151634
rect 438646 151398 438882 151634
rect 438326 115718 438562 115954
rect 438646 115718 438882 115954
rect 438326 115398 438562 115634
rect 438646 115398 438882 115634
rect 438326 79718 438562 79954
rect 438646 79718 438882 79954
rect 438326 79398 438562 79634
rect 438646 79398 438882 79634
rect 438326 43718 438562 43954
rect 438646 43718 438882 43954
rect 438326 43398 438562 43634
rect 438646 43398 438882 43634
rect 438326 7718 438562 7954
rect 438646 7718 438882 7954
rect 438326 7398 438562 7634
rect 438646 7398 438882 7634
rect 438326 -1542 438562 -1306
rect 438646 -1542 438882 -1306
rect 438326 -1862 438562 -1626
rect 438646 -1862 438882 -1626
rect 442826 706522 443062 706758
rect 443146 706522 443382 706758
rect 442826 706202 443062 706438
rect 443146 706202 443382 706438
rect 442826 696218 443062 696454
rect 443146 696218 443382 696454
rect 442826 695898 443062 696134
rect 443146 695898 443382 696134
rect 442826 660218 443062 660454
rect 443146 660218 443382 660454
rect 442826 659898 443062 660134
rect 443146 659898 443382 660134
rect 442826 624218 443062 624454
rect 443146 624218 443382 624454
rect 442826 623898 443062 624134
rect 443146 623898 443382 624134
rect 442826 588218 443062 588454
rect 443146 588218 443382 588454
rect 442826 587898 443062 588134
rect 443146 587898 443382 588134
rect 442826 552218 443062 552454
rect 443146 552218 443382 552454
rect 442826 551898 443062 552134
rect 443146 551898 443382 552134
rect 442826 516218 443062 516454
rect 443146 516218 443382 516454
rect 442826 515898 443062 516134
rect 443146 515898 443382 516134
rect 442826 480218 443062 480454
rect 443146 480218 443382 480454
rect 442826 479898 443062 480134
rect 443146 479898 443382 480134
rect 442826 444218 443062 444454
rect 443146 444218 443382 444454
rect 442826 443898 443062 444134
rect 443146 443898 443382 444134
rect 442826 408218 443062 408454
rect 443146 408218 443382 408454
rect 442826 407898 443062 408134
rect 443146 407898 443382 408134
rect 442826 372218 443062 372454
rect 443146 372218 443382 372454
rect 442826 371898 443062 372134
rect 443146 371898 443382 372134
rect 442826 336218 443062 336454
rect 443146 336218 443382 336454
rect 442826 335898 443062 336134
rect 443146 335898 443382 336134
rect 442826 300218 443062 300454
rect 443146 300218 443382 300454
rect 442826 299898 443062 300134
rect 443146 299898 443382 300134
rect 442826 264218 443062 264454
rect 443146 264218 443382 264454
rect 442826 263898 443062 264134
rect 443146 263898 443382 264134
rect 442826 228218 443062 228454
rect 443146 228218 443382 228454
rect 442826 227898 443062 228134
rect 443146 227898 443382 228134
rect 442826 192218 443062 192454
rect 443146 192218 443382 192454
rect 442826 191898 443062 192134
rect 443146 191898 443382 192134
rect 442826 156218 443062 156454
rect 443146 156218 443382 156454
rect 442826 155898 443062 156134
rect 443146 155898 443382 156134
rect 442826 120218 443062 120454
rect 443146 120218 443382 120454
rect 442826 119898 443062 120134
rect 443146 119898 443382 120134
rect 442826 84218 443062 84454
rect 443146 84218 443382 84454
rect 442826 83898 443062 84134
rect 443146 83898 443382 84134
rect 442826 48218 443062 48454
rect 443146 48218 443382 48454
rect 442826 47898 443062 48134
rect 443146 47898 443382 48134
rect 442826 12218 443062 12454
rect 443146 12218 443382 12454
rect 442826 11898 443062 12134
rect 443146 11898 443382 12134
rect 442826 -2502 443062 -2266
rect 443146 -2502 443382 -2266
rect 442826 -2822 443062 -2586
rect 443146 -2822 443382 -2586
rect 447326 707482 447562 707718
rect 447646 707482 447882 707718
rect 447326 707162 447562 707398
rect 447646 707162 447882 707398
rect 447326 700718 447562 700954
rect 447646 700718 447882 700954
rect 447326 700398 447562 700634
rect 447646 700398 447882 700634
rect 447326 664718 447562 664954
rect 447646 664718 447882 664954
rect 447326 664398 447562 664634
rect 447646 664398 447882 664634
rect 447326 628718 447562 628954
rect 447646 628718 447882 628954
rect 447326 628398 447562 628634
rect 447646 628398 447882 628634
rect 447326 592718 447562 592954
rect 447646 592718 447882 592954
rect 447326 592398 447562 592634
rect 447646 592398 447882 592634
rect 447326 556718 447562 556954
rect 447646 556718 447882 556954
rect 447326 556398 447562 556634
rect 447646 556398 447882 556634
rect 447326 520718 447562 520954
rect 447646 520718 447882 520954
rect 447326 520398 447562 520634
rect 447646 520398 447882 520634
rect 447326 484718 447562 484954
rect 447646 484718 447882 484954
rect 447326 484398 447562 484634
rect 447646 484398 447882 484634
rect 447326 448718 447562 448954
rect 447646 448718 447882 448954
rect 447326 448398 447562 448634
rect 447646 448398 447882 448634
rect 447326 412718 447562 412954
rect 447646 412718 447882 412954
rect 447326 412398 447562 412634
rect 447646 412398 447882 412634
rect 447326 376718 447562 376954
rect 447646 376718 447882 376954
rect 447326 376398 447562 376634
rect 447646 376398 447882 376634
rect 447326 340718 447562 340954
rect 447646 340718 447882 340954
rect 447326 340398 447562 340634
rect 447646 340398 447882 340634
rect 447326 304718 447562 304954
rect 447646 304718 447882 304954
rect 447326 304398 447562 304634
rect 447646 304398 447882 304634
rect 447326 268718 447562 268954
rect 447646 268718 447882 268954
rect 447326 268398 447562 268634
rect 447646 268398 447882 268634
rect 447326 232718 447562 232954
rect 447646 232718 447882 232954
rect 447326 232398 447562 232634
rect 447646 232398 447882 232634
rect 447326 196718 447562 196954
rect 447646 196718 447882 196954
rect 447326 196398 447562 196634
rect 447646 196398 447882 196634
rect 447326 160718 447562 160954
rect 447646 160718 447882 160954
rect 447326 160398 447562 160634
rect 447646 160398 447882 160634
rect 447326 124718 447562 124954
rect 447646 124718 447882 124954
rect 447326 124398 447562 124634
rect 447646 124398 447882 124634
rect 447326 88718 447562 88954
rect 447646 88718 447882 88954
rect 447326 88398 447562 88634
rect 447646 88398 447882 88634
rect 447326 52718 447562 52954
rect 447646 52718 447882 52954
rect 447326 52398 447562 52634
rect 447646 52398 447882 52634
rect 447326 16718 447562 16954
rect 447646 16718 447882 16954
rect 447326 16398 447562 16634
rect 447646 16398 447882 16634
rect 447326 -3462 447562 -3226
rect 447646 -3462 447882 -3226
rect 447326 -3782 447562 -3546
rect 447646 -3782 447882 -3546
rect 451826 708442 452062 708678
rect 452146 708442 452382 708678
rect 451826 708122 452062 708358
rect 452146 708122 452382 708358
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -4422 452062 -4186
rect 452146 -4422 452382 -4186
rect 451826 -4742 452062 -4506
rect 452146 -4742 452382 -4506
rect 456326 709402 456562 709638
rect 456646 709402 456882 709638
rect 456326 709082 456562 709318
rect 456646 709082 456882 709318
rect 456326 673718 456562 673954
rect 456646 673718 456882 673954
rect 456326 673398 456562 673634
rect 456646 673398 456882 673634
rect 456326 637718 456562 637954
rect 456646 637718 456882 637954
rect 456326 637398 456562 637634
rect 456646 637398 456882 637634
rect 456326 601718 456562 601954
rect 456646 601718 456882 601954
rect 456326 601398 456562 601634
rect 456646 601398 456882 601634
rect 456326 565718 456562 565954
rect 456646 565718 456882 565954
rect 456326 565398 456562 565634
rect 456646 565398 456882 565634
rect 456326 529718 456562 529954
rect 456646 529718 456882 529954
rect 456326 529398 456562 529634
rect 456646 529398 456882 529634
rect 456326 493718 456562 493954
rect 456646 493718 456882 493954
rect 456326 493398 456562 493634
rect 456646 493398 456882 493634
rect 456326 457718 456562 457954
rect 456646 457718 456882 457954
rect 456326 457398 456562 457634
rect 456646 457398 456882 457634
rect 456326 421718 456562 421954
rect 456646 421718 456882 421954
rect 456326 421398 456562 421634
rect 456646 421398 456882 421634
rect 456326 385718 456562 385954
rect 456646 385718 456882 385954
rect 456326 385398 456562 385634
rect 456646 385398 456882 385634
rect 456326 349718 456562 349954
rect 456646 349718 456882 349954
rect 456326 349398 456562 349634
rect 456646 349398 456882 349634
rect 456326 313718 456562 313954
rect 456646 313718 456882 313954
rect 456326 313398 456562 313634
rect 456646 313398 456882 313634
rect 456326 277718 456562 277954
rect 456646 277718 456882 277954
rect 456326 277398 456562 277634
rect 456646 277398 456882 277634
rect 456326 241718 456562 241954
rect 456646 241718 456882 241954
rect 456326 241398 456562 241634
rect 456646 241398 456882 241634
rect 456326 205718 456562 205954
rect 456646 205718 456882 205954
rect 456326 205398 456562 205634
rect 456646 205398 456882 205634
rect 456326 169718 456562 169954
rect 456646 169718 456882 169954
rect 456326 169398 456562 169634
rect 456646 169398 456882 169634
rect 456326 133718 456562 133954
rect 456646 133718 456882 133954
rect 456326 133398 456562 133634
rect 456646 133398 456882 133634
rect 456326 97718 456562 97954
rect 456646 97718 456882 97954
rect 456326 97398 456562 97634
rect 456646 97398 456882 97634
rect 456326 61718 456562 61954
rect 456646 61718 456882 61954
rect 456326 61398 456562 61634
rect 456646 61398 456882 61634
rect 456326 25718 456562 25954
rect 456646 25718 456882 25954
rect 456326 25398 456562 25634
rect 456646 25398 456882 25634
rect 456326 -5382 456562 -5146
rect 456646 -5382 456882 -5146
rect 456326 -5702 456562 -5466
rect 456646 -5702 456882 -5466
rect 460826 710362 461062 710598
rect 461146 710362 461382 710598
rect 460826 710042 461062 710278
rect 461146 710042 461382 710278
rect 460826 678218 461062 678454
rect 461146 678218 461382 678454
rect 460826 677898 461062 678134
rect 461146 677898 461382 678134
rect 460826 642218 461062 642454
rect 461146 642218 461382 642454
rect 460826 641898 461062 642134
rect 461146 641898 461382 642134
rect 460826 606218 461062 606454
rect 461146 606218 461382 606454
rect 460826 605898 461062 606134
rect 461146 605898 461382 606134
rect 460826 570218 461062 570454
rect 461146 570218 461382 570454
rect 460826 569898 461062 570134
rect 461146 569898 461382 570134
rect 460826 534218 461062 534454
rect 461146 534218 461382 534454
rect 460826 533898 461062 534134
rect 461146 533898 461382 534134
rect 460826 498218 461062 498454
rect 461146 498218 461382 498454
rect 460826 497898 461062 498134
rect 461146 497898 461382 498134
rect 460826 462218 461062 462454
rect 461146 462218 461382 462454
rect 460826 461898 461062 462134
rect 461146 461898 461382 462134
rect 460826 426218 461062 426454
rect 461146 426218 461382 426454
rect 460826 425898 461062 426134
rect 461146 425898 461382 426134
rect 460826 390218 461062 390454
rect 461146 390218 461382 390454
rect 460826 389898 461062 390134
rect 461146 389898 461382 390134
rect 460826 354218 461062 354454
rect 461146 354218 461382 354454
rect 460826 353898 461062 354134
rect 461146 353898 461382 354134
rect 460826 318218 461062 318454
rect 461146 318218 461382 318454
rect 460826 317898 461062 318134
rect 461146 317898 461382 318134
rect 460826 282218 461062 282454
rect 461146 282218 461382 282454
rect 460826 281898 461062 282134
rect 461146 281898 461382 282134
rect 460826 246218 461062 246454
rect 461146 246218 461382 246454
rect 460826 245898 461062 246134
rect 461146 245898 461382 246134
rect 460826 210218 461062 210454
rect 461146 210218 461382 210454
rect 460826 209898 461062 210134
rect 461146 209898 461382 210134
rect 460826 174218 461062 174454
rect 461146 174218 461382 174454
rect 460826 173898 461062 174134
rect 461146 173898 461382 174134
rect 460826 138218 461062 138454
rect 461146 138218 461382 138454
rect 460826 137898 461062 138134
rect 461146 137898 461382 138134
rect 460826 102218 461062 102454
rect 461146 102218 461382 102454
rect 460826 101898 461062 102134
rect 461146 101898 461382 102134
rect 460826 66218 461062 66454
rect 461146 66218 461382 66454
rect 460826 65898 461062 66134
rect 461146 65898 461382 66134
rect 460826 30218 461062 30454
rect 461146 30218 461382 30454
rect 460826 29898 461062 30134
rect 461146 29898 461382 30134
rect 460826 -6342 461062 -6106
rect 461146 -6342 461382 -6106
rect 460826 -6662 461062 -6426
rect 461146 -6662 461382 -6426
rect 465326 711322 465562 711558
rect 465646 711322 465882 711558
rect 465326 711002 465562 711238
rect 465646 711002 465882 711238
rect 465326 682718 465562 682954
rect 465646 682718 465882 682954
rect 465326 682398 465562 682634
rect 465646 682398 465882 682634
rect 465326 646718 465562 646954
rect 465646 646718 465882 646954
rect 465326 646398 465562 646634
rect 465646 646398 465882 646634
rect 465326 610718 465562 610954
rect 465646 610718 465882 610954
rect 465326 610398 465562 610634
rect 465646 610398 465882 610634
rect 465326 574718 465562 574954
rect 465646 574718 465882 574954
rect 465326 574398 465562 574634
rect 465646 574398 465882 574634
rect 465326 538718 465562 538954
rect 465646 538718 465882 538954
rect 465326 538398 465562 538634
rect 465646 538398 465882 538634
rect 465326 502718 465562 502954
rect 465646 502718 465882 502954
rect 465326 502398 465562 502634
rect 465646 502398 465882 502634
rect 465326 466718 465562 466954
rect 465646 466718 465882 466954
rect 465326 466398 465562 466634
rect 465646 466398 465882 466634
rect 465326 430718 465562 430954
rect 465646 430718 465882 430954
rect 465326 430398 465562 430634
rect 465646 430398 465882 430634
rect 465326 394718 465562 394954
rect 465646 394718 465882 394954
rect 465326 394398 465562 394634
rect 465646 394398 465882 394634
rect 465326 358718 465562 358954
rect 465646 358718 465882 358954
rect 465326 358398 465562 358634
rect 465646 358398 465882 358634
rect 465326 322718 465562 322954
rect 465646 322718 465882 322954
rect 465326 322398 465562 322634
rect 465646 322398 465882 322634
rect 465326 286718 465562 286954
rect 465646 286718 465882 286954
rect 465326 286398 465562 286634
rect 465646 286398 465882 286634
rect 465326 250718 465562 250954
rect 465646 250718 465882 250954
rect 465326 250398 465562 250634
rect 465646 250398 465882 250634
rect 465326 214718 465562 214954
rect 465646 214718 465882 214954
rect 465326 214398 465562 214634
rect 465646 214398 465882 214634
rect 465326 178718 465562 178954
rect 465646 178718 465882 178954
rect 465326 178398 465562 178634
rect 465646 178398 465882 178634
rect 465326 142718 465562 142954
rect 465646 142718 465882 142954
rect 465326 142398 465562 142634
rect 465646 142398 465882 142634
rect 465326 106718 465562 106954
rect 465646 106718 465882 106954
rect 465326 106398 465562 106634
rect 465646 106398 465882 106634
rect 465326 70718 465562 70954
rect 465646 70718 465882 70954
rect 465326 70398 465562 70634
rect 465646 70398 465882 70634
rect 465326 34718 465562 34954
rect 465646 34718 465882 34954
rect 465326 34398 465562 34634
rect 465646 34398 465882 34634
rect 465326 -7302 465562 -7066
rect 465646 -7302 465882 -7066
rect 465326 -7622 465562 -7386
rect 465646 -7622 465882 -7386
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 474326 705562 474562 705798
rect 474646 705562 474882 705798
rect 474326 705242 474562 705478
rect 474646 705242 474882 705478
rect 474326 691718 474562 691954
rect 474646 691718 474882 691954
rect 474326 691398 474562 691634
rect 474646 691398 474882 691634
rect 474326 655718 474562 655954
rect 474646 655718 474882 655954
rect 474326 655398 474562 655634
rect 474646 655398 474882 655634
rect 474326 619718 474562 619954
rect 474646 619718 474882 619954
rect 474326 619398 474562 619634
rect 474646 619398 474882 619634
rect 474326 583718 474562 583954
rect 474646 583718 474882 583954
rect 474326 583398 474562 583634
rect 474646 583398 474882 583634
rect 474326 547718 474562 547954
rect 474646 547718 474882 547954
rect 474326 547398 474562 547634
rect 474646 547398 474882 547634
rect 474326 511718 474562 511954
rect 474646 511718 474882 511954
rect 474326 511398 474562 511634
rect 474646 511398 474882 511634
rect 474326 475718 474562 475954
rect 474646 475718 474882 475954
rect 474326 475398 474562 475634
rect 474646 475398 474882 475634
rect 474326 439718 474562 439954
rect 474646 439718 474882 439954
rect 474326 439398 474562 439634
rect 474646 439398 474882 439634
rect 474326 403718 474562 403954
rect 474646 403718 474882 403954
rect 474326 403398 474562 403634
rect 474646 403398 474882 403634
rect 474326 367718 474562 367954
rect 474646 367718 474882 367954
rect 474326 367398 474562 367634
rect 474646 367398 474882 367634
rect 474326 331718 474562 331954
rect 474646 331718 474882 331954
rect 474326 331398 474562 331634
rect 474646 331398 474882 331634
rect 474326 295718 474562 295954
rect 474646 295718 474882 295954
rect 474326 295398 474562 295634
rect 474646 295398 474882 295634
rect 474326 259718 474562 259954
rect 474646 259718 474882 259954
rect 474326 259398 474562 259634
rect 474646 259398 474882 259634
rect 474326 223718 474562 223954
rect 474646 223718 474882 223954
rect 474326 223398 474562 223634
rect 474646 223398 474882 223634
rect 474326 187718 474562 187954
rect 474646 187718 474882 187954
rect 474326 187398 474562 187634
rect 474646 187398 474882 187634
rect 474326 151718 474562 151954
rect 474646 151718 474882 151954
rect 474326 151398 474562 151634
rect 474646 151398 474882 151634
rect 474326 115718 474562 115954
rect 474646 115718 474882 115954
rect 474326 115398 474562 115634
rect 474646 115398 474882 115634
rect 474326 79718 474562 79954
rect 474646 79718 474882 79954
rect 474326 79398 474562 79634
rect 474646 79398 474882 79634
rect 474326 43718 474562 43954
rect 474646 43718 474882 43954
rect 474326 43398 474562 43634
rect 474646 43398 474882 43634
rect 474326 7718 474562 7954
rect 474646 7718 474882 7954
rect 474326 7398 474562 7634
rect 474646 7398 474882 7634
rect 474326 -1542 474562 -1306
rect 474646 -1542 474882 -1306
rect 474326 -1862 474562 -1626
rect 474646 -1862 474882 -1626
rect 478826 706522 479062 706758
rect 479146 706522 479382 706758
rect 478826 706202 479062 706438
rect 479146 706202 479382 706438
rect 478826 696218 479062 696454
rect 479146 696218 479382 696454
rect 478826 695898 479062 696134
rect 479146 695898 479382 696134
rect 478826 660218 479062 660454
rect 479146 660218 479382 660454
rect 478826 659898 479062 660134
rect 479146 659898 479382 660134
rect 478826 624218 479062 624454
rect 479146 624218 479382 624454
rect 478826 623898 479062 624134
rect 479146 623898 479382 624134
rect 478826 588218 479062 588454
rect 479146 588218 479382 588454
rect 478826 587898 479062 588134
rect 479146 587898 479382 588134
rect 478826 552218 479062 552454
rect 479146 552218 479382 552454
rect 478826 551898 479062 552134
rect 479146 551898 479382 552134
rect 478826 516218 479062 516454
rect 479146 516218 479382 516454
rect 478826 515898 479062 516134
rect 479146 515898 479382 516134
rect 478826 480218 479062 480454
rect 479146 480218 479382 480454
rect 478826 479898 479062 480134
rect 479146 479898 479382 480134
rect 478826 444218 479062 444454
rect 479146 444218 479382 444454
rect 478826 443898 479062 444134
rect 479146 443898 479382 444134
rect 478826 408218 479062 408454
rect 479146 408218 479382 408454
rect 478826 407898 479062 408134
rect 479146 407898 479382 408134
rect 478826 372218 479062 372454
rect 479146 372218 479382 372454
rect 478826 371898 479062 372134
rect 479146 371898 479382 372134
rect 478826 336218 479062 336454
rect 479146 336218 479382 336454
rect 478826 335898 479062 336134
rect 479146 335898 479382 336134
rect 478826 300218 479062 300454
rect 479146 300218 479382 300454
rect 478826 299898 479062 300134
rect 479146 299898 479382 300134
rect 478826 264218 479062 264454
rect 479146 264218 479382 264454
rect 478826 263898 479062 264134
rect 479146 263898 479382 264134
rect 478826 228218 479062 228454
rect 479146 228218 479382 228454
rect 478826 227898 479062 228134
rect 479146 227898 479382 228134
rect 478826 192218 479062 192454
rect 479146 192218 479382 192454
rect 478826 191898 479062 192134
rect 479146 191898 479382 192134
rect 478826 156218 479062 156454
rect 479146 156218 479382 156454
rect 478826 155898 479062 156134
rect 479146 155898 479382 156134
rect 478826 120218 479062 120454
rect 479146 120218 479382 120454
rect 478826 119898 479062 120134
rect 479146 119898 479382 120134
rect 478826 84218 479062 84454
rect 479146 84218 479382 84454
rect 478826 83898 479062 84134
rect 479146 83898 479382 84134
rect 478826 48218 479062 48454
rect 479146 48218 479382 48454
rect 478826 47898 479062 48134
rect 479146 47898 479382 48134
rect 478826 12218 479062 12454
rect 479146 12218 479382 12454
rect 478826 11898 479062 12134
rect 479146 11898 479382 12134
rect 478826 -2502 479062 -2266
rect 479146 -2502 479382 -2266
rect 478826 -2822 479062 -2586
rect 479146 -2822 479382 -2586
rect 483326 707482 483562 707718
rect 483646 707482 483882 707718
rect 483326 707162 483562 707398
rect 483646 707162 483882 707398
rect 483326 700718 483562 700954
rect 483646 700718 483882 700954
rect 483326 700398 483562 700634
rect 483646 700398 483882 700634
rect 483326 664718 483562 664954
rect 483646 664718 483882 664954
rect 483326 664398 483562 664634
rect 483646 664398 483882 664634
rect 483326 628718 483562 628954
rect 483646 628718 483882 628954
rect 483326 628398 483562 628634
rect 483646 628398 483882 628634
rect 483326 592718 483562 592954
rect 483646 592718 483882 592954
rect 483326 592398 483562 592634
rect 483646 592398 483882 592634
rect 483326 556718 483562 556954
rect 483646 556718 483882 556954
rect 483326 556398 483562 556634
rect 483646 556398 483882 556634
rect 483326 520718 483562 520954
rect 483646 520718 483882 520954
rect 483326 520398 483562 520634
rect 483646 520398 483882 520634
rect 483326 484718 483562 484954
rect 483646 484718 483882 484954
rect 483326 484398 483562 484634
rect 483646 484398 483882 484634
rect 483326 448718 483562 448954
rect 483646 448718 483882 448954
rect 483326 448398 483562 448634
rect 483646 448398 483882 448634
rect 483326 412718 483562 412954
rect 483646 412718 483882 412954
rect 483326 412398 483562 412634
rect 483646 412398 483882 412634
rect 483326 376718 483562 376954
rect 483646 376718 483882 376954
rect 483326 376398 483562 376634
rect 483646 376398 483882 376634
rect 483326 340718 483562 340954
rect 483646 340718 483882 340954
rect 483326 340398 483562 340634
rect 483646 340398 483882 340634
rect 483326 304718 483562 304954
rect 483646 304718 483882 304954
rect 483326 304398 483562 304634
rect 483646 304398 483882 304634
rect 483326 268718 483562 268954
rect 483646 268718 483882 268954
rect 483326 268398 483562 268634
rect 483646 268398 483882 268634
rect 483326 232718 483562 232954
rect 483646 232718 483882 232954
rect 483326 232398 483562 232634
rect 483646 232398 483882 232634
rect 483326 196718 483562 196954
rect 483646 196718 483882 196954
rect 483326 196398 483562 196634
rect 483646 196398 483882 196634
rect 483326 160718 483562 160954
rect 483646 160718 483882 160954
rect 483326 160398 483562 160634
rect 483646 160398 483882 160634
rect 483326 124718 483562 124954
rect 483646 124718 483882 124954
rect 483326 124398 483562 124634
rect 483646 124398 483882 124634
rect 483326 88718 483562 88954
rect 483646 88718 483882 88954
rect 483326 88398 483562 88634
rect 483646 88398 483882 88634
rect 483326 52718 483562 52954
rect 483646 52718 483882 52954
rect 483326 52398 483562 52634
rect 483646 52398 483882 52634
rect 483326 16718 483562 16954
rect 483646 16718 483882 16954
rect 483326 16398 483562 16634
rect 483646 16398 483882 16634
rect 483326 -3462 483562 -3226
rect 483646 -3462 483882 -3226
rect 483326 -3782 483562 -3546
rect 483646 -3782 483882 -3546
rect 487826 708442 488062 708678
rect 488146 708442 488382 708678
rect 487826 708122 488062 708358
rect 488146 708122 488382 708358
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -4422 488062 -4186
rect 488146 -4422 488382 -4186
rect 487826 -4742 488062 -4506
rect 488146 -4742 488382 -4506
rect 492326 709402 492562 709638
rect 492646 709402 492882 709638
rect 492326 709082 492562 709318
rect 492646 709082 492882 709318
rect 492326 673718 492562 673954
rect 492646 673718 492882 673954
rect 492326 673398 492562 673634
rect 492646 673398 492882 673634
rect 492326 637718 492562 637954
rect 492646 637718 492882 637954
rect 492326 637398 492562 637634
rect 492646 637398 492882 637634
rect 492326 601718 492562 601954
rect 492646 601718 492882 601954
rect 492326 601398 492562 601634
rect 492646 601398 492882 601634
rect 492326 565718 492562 565954
rect 492646 565718 492882 565954
rect 492326 565398 492562 565634
rect 492646 565398 492882 565634
rect 492326 529718 492562 529954
rect 492646 529718 492882 529954
rect 492326 529398 492562 529634
rect 492646 529398 492882 529634
rect 492326 493718 492562 493954
rect 492646 493718 492882 493954
rect 492326 493398 492562 493634
rect 492646 493398 492882 493634
rect 492326 457718 492562 457954
rect 492646 457718 492882 457954
rect 492326 457398 492562 457634
rect 492646 457398 492882 457634
rect 492326 421718 492562 421954
rect 492646 421718 492882 421954
rect 492326 421398 492562 421634
rect 492646 421398 492882 421634
rect 492326 385718 492562 385954
rect 492646 385718 492882 385954
rect 492326 385398 492562 385634
rect 492646 385398 492882 385634
rect 492326 349718 492562 349954
rect 492646 349718 492882 349954
rect 492326 349398 492562 349634
rect 492646 349398 492882 349634
rect 492326 313718 492562 313954
rect 492646 313718 492882 313954
rect 492326 313398 492562 313634
rect 492646 313398 492882 313634
rect 492326 277718 492562 277954
rect 492646 277718 492882 277954
rect 492326 277398 492562 277634
rect 492646 277398 492882 277634
rect 492326 241718 492562 241954
rect 492646 241718 492882 241954
rect 492326 241398 492562 241634
rect 492646 241398 492882 241634
rect 492326 205718 492562 205954
rect 492646 205718 492882 205954
rect 492326 205398 492562 205634
rect 492646 205398 492882 205634
rect 492326 169718 492562 169954
rect 492646 169718 492882 169954
rect 492326 169398 492562 169634
rect 492646 169398 492882 169634
rect 492326 133718 492562 133954
rect 492646 133718 492882 133954
rect 492326 133398 492562 133634
rect 492646 133398 492882 133634
rect 492326 97718 492562 97954
rect 492646 97718 492882 97954
rect 492326 97398 492562 97634
rect 492646 97398 492882 97634
rect 492326 61718 492562 61954
rect 492646 61718 492882 61954
rect 492326 61398 492562 61634
rect 492646 61398 492882 61634
rect 492326 25718 492562 25954
rect 492646 25718 492882 25954
rect 492326 25398 492562 25634
rect 492646 25398 492882 25634
rect 492326 -5382 492562 -5146
rect 492646 -5382 492882 -5146
rect 492326 -5702 492562 -5466
rect 492646 -5702 492882 -5466
rect 496826 710362 497062 710598
rect 497146 710362 497382 710598
rect 496826 710042 497062 710278
rect 497146 710042 497382 710278
rect 496826 678218 497062 678454
rect 497146 678218 497382 678454
rect 496826 677898 497062 678134
rect 497146 677898 497382 678134
rect 496826 642218 497062 642454
rect 497146 642218 497382 642454
rect 496826 641898 497062 642134
rect 497146 641898 497382 642134
rect 496826 606218 497062 606454
rect 497146 606218 497382 606454
rect 496826 605898 497062 606134
rect 497146 605898 497382 606134
rect 496826 570218 497062 570454
rect 497146 570218 497382 570454
rect 496826 569898 497062 570134
rect 497146 569898 497382 570134
rect 496826 534218 497062 534454
rect 497146 534218 497382 534454
rect 496826 533898 497062 534134
rect 497146 533898 497382 534134
rect 496826 498218 497062 498454
rect 497146 498218 497382 498454
rect 496826 497898 497062 498134
rect 497146 497898 497382 498134
rect 496826 462218 497062 462454
rect 497146 462218 497382 462454
rect 496826 461898 497062 462134
rect 497146 461898 497382 462134
rect 496826 426218 497062 426454
rect 497146 426218 497382 426454
rect 496826 425898 497062 426134
rect 497146 425898 497382 426134
rect 496826 390218 497062 390454
rect 497146 390218 497382 390454
rect 496826 389898 497062 390134
rect 497146 389898 497382 390134
rect 496826 354218 497062 354454
rect 497146 354218 497382 354454
rect 496826 353898 497062 354134
rect 497146 353898 497382 354134
rect 496826 318218 497062 318454
rect 497146 318218 497382 318454
rect 496826 317898 497062 318134
rect 497146 317898 497382 318134
rect 496826 282218 497062 282454
rect 497146 282218 497382 282454
rect 496826 281898 497062 282134
rect 497146 281898 497382 282134
rect 496826 246218 497062 246454
rect 497146 246218 497382 246454
rect 496826 245898 497062 246134
rect 497146 245898 497382 246134
rect 496826 210218 497062 210454
rect 497146 210218 497382 210454
rect 496826 209898 497062 210134
rect 497146 209898 497382 210134
rect 496826 174218 497062 174454
rect 497146 174218 497382 174454
rect 496826 173898 497062 174134
rect 497146 173898 497382 174134
rect 496826 138218 497062 138454
rect 497146 138218 497382 138454
rect 496826 137898 497062 138134
rect 497146 137898 497382 138134
rect 496826 102218 497062 102454
rect 497146 102218 497382 102454
rect 496826 101898 497062 102134
rect 497146 101898 497382 102134
rect 496826 66218 497062 66454
rect 497146 66218 497382 66454
rect 496826 65898 497062 66134
rect 497146 65898 497382 66134
rect 496826 30218 497062 30454
rect 497146 30218 497382 30454
rect 496826 29898 497062 30134
rect 497146 29898 497382 30134
rect 496826 -6342 497062 -6106
rect 497146 -6342 497382 -6106
rect 496826 -6662 497062 -6426
rect 497146 -6662 497382 -6426
rect 501326 711322 501562 711558
rect 501646 711322 501882 711558
rect 501326 711002 501562 711238
rect 501646 711002 501882 711238
rect 501326 682718 501562 682954
rect 501646 682718 501882 682954
rect 501326 682398 501562 682634
rect 501646 682398 501882 682634
rect 501326 646718 501562 646954
rect 501646 646718 501882 646954
rect 501326 646398 501562 646634
rect 501646 646398 501882 646634
rect 501326 610718 501562 610954
rect 501646 610718 501882 610954
rect 501326 610398 501562 610634
rect 501646 610398 501882 610634
rect 501326 574718 501562 574954
rect 501646 574718 501882 574954
rect 501326 574398 501562 574634
rect 501646 574398 501882 574634
rect 501326 538718 501562 538954
rect 501646 538718 501882 538954
rect 501326 538398 501562 538634
rect 501646 538398 501882 538634
rect 501326 502718 501562 502954
rect 501646 502718 501882 502954
rect 501326 502398 501562 502634
rect 501646 502398 501882 502634
rect 501326 466718 501562 466954
rect 501646 466718 501882 466954
rect 501326 466398 501562 466634
rect 501646 466398 501882 466634
rect 501326 430718 501562 430954
rect 501646 430718 501882 430954
rect 501326 430398 501562 430634
rect 501646 430398 501882 430634
rect 501326 394718 501562 394954
rect 501646 394718 501882 394954
rect 501326 394398 501562 394634
rect 501646 394398 501882 394634
rect 501326 358718 501562 358954
rect 501646 358718 501882 358954
rect 501326 358398 501562 358634
rect 501646 358398 501882 358634
rect 501326 322718 501562 322954
rect 501646 322718 501882 322954
rect 501326 322398 501562 322634
rect 501646 322398 501882 322634
rect 501326 286718 501562 286954
rect 501646 286718 501882 286954
rect 501326 286398 501562 286634
rect 501646 286398 501882 286634
rect 501326 250718 501562 250954
rect 501646 250718 501882 250954
rect 501326 250398 501562 250634
rect 501646 250398 501882 250634
rect 501326 214718 501562 214954
rect 501646 214718 501882 214954
rect 501326 214398 501562 214634
rect 501646 214398 501882 214634
rect 501326 178718 501562 178954
rect 501646 178718 501882 178954
rect 501326 178398 501562 178634
rect 501646 178398 501882 178634
rect 501326 142718 501562 142954
rect 501646 142718 501882 142954
rect 501326 142398 501562 142634
rect 501646 142398 501882 142634
rect 501326 106718 501562 106954
rect 501646 106718 501882 106954
rect 501326 106398 501562 106634
rect 501646 106398 501882 106634
rect 501326 70718 501562 70954
rect 501646 70718 501882 70954
rect 501326 70398 501562 70634
rect 501646 70398 501882 70634
rect 501326 34718 501562 34954
rect 501646 34718 501882 34954
rect 501326 34398 501562 34634
rect 501646 34398 501882 34634
rect 501326 -7302 501562 -7066
rect 501646 -7302 501882 -7066
rect 501326 -7622 501562 -7386
rect 501646 -7622 501882 -7386
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 510326 705562 510562 705798
rect 510646 705562 510882 705798
rect 510326 705242 510562 705478
rect 510646 705242 510882 705478
rect 510326 691718 510562 691954
rect 510646 691718 510882 691954
rect 510326 691398 510562 691634
rect 510646 691398 510882 691634
rect 510326 655718 510562 655954
rect 510646 655718 510882 655954
rect 510326 655398 510562 655634
rect 510646 655398 510882 655634
rect 510326 619718 510562 619954
rect 510646 619718 510882 619954
rect 510326 619398 510562 619634
rect 510646 619398 510882 619634
rect 510326 583718 510562 583954
rect 510646 583718 510882 583954
rect 510326 583398 510562 583634
rect 510646 583398 510882 583634
rect 510326 547718 510562 547954
rect 510646 547718 510882 547954
rect 510326 547398 510562 547634
rect 510646 547398 510882 547634
rect 510326 511718 510562 511954
rect 510646 511718 510882 511954
rect 510326 511398 510562 511634
rect 510646 511398 510882 511634
rect 510326 475718 510562 475954
rect 510646 475718 510882 475954
rect 510326 475398 510562 475634
rect 510646 475398 510882 475634
rect 510326 439718 510562 439954
rect 510646 439718 510882 439954
rect 510326 439398 510562 439634
rect 510646 439398 510882 439634
rect 510326 403718 510562 403954
rect 510646 403718 510882 403954
rect 510326 403398 510562 403634
rect 510646 403398 510882 403634
rect 510326 367718 510562 367954
rect 510646 367718 510882 367954
rect 510326 367398 510562 367634
rect 510646 367398 510882 367634
rect 510326 331718 510562 331954
rect 510646 331718 510882 331954
rect 510326 331398 510562 331634
rect 510646 331398 510882 331634
rect 510326 295718 510562 295954
rect 510646 295718 510882 295954
rect 510326 295398 510562 295634
rect 510646 295398 510882 295634
rect 510326 259718 510562 259954
rect 510646 259718 510882 259954
rect 510326 259398 510562 259634
rect 510646 259398 510882 259634
rect 510326 223718 510562 223954
rect 510646 223718 510882 223954
rect 510326 223398 510562 223634
rect 510646 223398 510882 223634
rect 510326 187718 510562 187954
rect 510646 187718 510882 187954
rect 510326 187398 510562 187634
rect 510646 187398 510882 187634
rect 510326 151718 510562 151954
rect 510646 151718 510882 151954
rect 510326 151398 510562 151634
rect 510646 151398 510882 151634
rect 510326 115718 510562 115954
rect 510646 115718 510882 115954
rect 510326 115398 510562 115634
rect 510646 115398 510882 115634
rect 510326 79718 510562 79954
rect 510646 79718 510882 79954
rect 510326 79398 510562 79634
rect 510646 79398 510882 79634
rect 510326 43718 510562 43954
rect 510646 43718 510882 43954
rect 510326 43398 510562 43634
rect 510646 43398 510882 43634
rect 510326 7718 510562 7954
rect 510646 7718 510882 7954
rect 510326 7398 510562 7634
rect 510646 7398 510882 7634
rect 510326 -1542 510562 -1306
rect 510646 -1542 510882 -1306
rect 510326 -1862 510562 -1626
rect 510646 -1862 510882 -1626
rect 514826 706522 515062 706758
rect 515146 706522 515382 706758
rect 514826 706202 515062 706438
rect 515146 706202 515382 706438
rect 514826 696218 515062 696454
rect 515146 696218 515382 696454
rect 514826 695898 515062 696134
rect 515146 695898 515382 696134
rect 514826 660218 515062 660454
rect 515146 660218 515382 660454
rect 514826 659898 515062 660134
rect 515146 659898 515382 660134
rect 514826 624218 515062 624454
rect 515146 624218 515382 624454
rect 514826 623898 515062 624134
rect 515146 623898 515382 624134
rect 514826 588218 515062 588454
rect 515146 588218 515382 588454
rect 514826 587898 515062 588134
rect 515146 587898 515382 588134
rect 514826 552218 515062 552454
rect 515146 552218 515382 552454
rect 514826 551898 515062 552134
rect 515146 551898 515382 552134
rect 514826 516218 515062 516454
rect 515146 516218 515382 516454
rect 514826 515898 515062 516134
rect 515146 515898 515382 516134
rect 514826 480218 515062 480454
rect 515146 480218 515382 480454
rect 514826 479898 515062 480134
rect 515146 479898 515382 480134
rect 514826 444218 515062 444454
rect 515146 444218 515382 444454
rect 514826 443898 515062 444134
rect 515146 443898 515382 444134
rect 514826 408218 515062 408454
rect 515146 408218 515382 408454
rect 514826 407898 515062 408134
rect 515146 407898 515382 408134
rect 514826 372218 515062 372454
rect 515146 372218 515382 372454
rect 514826 371898 515062 372134
rect 515146 371898 515382 372134
rect 514826 336218 515062 336454
rect 515146 336218 515382 336454
rect 514826 335898 515062 336134
rect 515146 335898 515382 336134
rect 514826 300218 515062 300454
rect 515146 300218 515382 300454
rect 514826 299898 515062 300134
rect 515146 299898 515382 300134
rect 514826 264218 515062 264454
rect 515146 264218 515382 264454
rect 514826 263898 515062 264134
rect 515146 263898 515382 264134
rect 514826 228218 515062 228454
rect 515146 228218 515382 228454
rect 514826 227898 515062 228134
rect 515146 227898 515382 228134
rect 514826 192218 515062 192454
rect 515146 192218 515382 192454
rect 514826 191898 515062 192134
rect 515146 191898 515382 192134
rect 514826 156218 515062 156454
rect 515146 156218 515382 156454
rect 514826 155898 515062 156134
rect 515146 155898 515382 156134
rect 514826 120218 515062 120454
rect 515146 120218 515382 120454
rect 514826 119898 515062 120134
rect 515146 119898 515382 120134
rect 514826 84218 515062 84454
rect 515146 84218 515382 84454
rect 514826 83898 515062 84134
rect 515146 83898 515382 84134
rect 514826 48218 515062 48454
rect 515146 48218 515382 48454
rect 514826 47898 515062 48134
rect 515146 47898 515382 48134
rect 514826 12218 515062 12454
rect 515146 12218 515382 12454
rect 514826 11898 515062 12134
rect 515146 11898 515382 12134
rect 514826 -2502 515062 -2266
rect 515146 -2502 515382 -2266
rect 514826 -2822 515062 -2586
rect 515146 -2822 515382 -2586
rect 519326 707482 519562 707718
rect 519646 707482 519882 707718
rect 519326 707162 519562 707398
rect 519646 707162 519882 707398
rect 519326 700718 519562 700954
rect 519646 700718 519882 700954
rect 519326 700398 519562 700634
rect 519646 700398 519882 700634
rect 519326 664718 519562 664954
rect 519646 664718 519882 664954
rect 519326 664398 519562 664634
rect 519646 664398 519882 664634
rect 519326 628718 519562 628954
rect 519646 628718 519882 628954
rect 519326 628398 519562 628634
rect 519646 628398 519882 628634
rect 519326 592718 519562 592954
rect 519646 592718 519882 592954
rect 519326 592398 519562 592634
rect 519646 592398 519882 592634
rect 519326 556718 519562 556954
rect 519646 556718 519882 556954
rect 519326 556398 519562 556634
rect 519646 556398 519882 556634
rect 519326 520718 519562 520954
rect 519646 520718 519882 520954
rect 519326 520398 519562 520634
rect 519646 520398 519882 520634
rect 519326 484718 519562 484954
rect 519646 484718 519882 484954
rect 519326 484398 519562 484634
rect 519646 484398 519882 484634
rect 519326 448718 519562 448954
rect 519646 448718 519882 448954
rect 519326 448398 519562 448634
rect 519646 448398 519882 448634
rect 519326 412718 519562 412954
rect 519646 412718 519882 412954
rect 519326 412398 519562 412634
rect 519646 412398 519882 412634
rect 519326 376718 519562 376954
rect 519646 376718 519882 376954
rect 519326 376398 519562 376634
rect 519646 376398 519882 376634
rect 519326 340718 519562 340954
rect 519646 340718 519882 340954
rect 519326 340398 519562 340634
rect 519646 340398 519882 340634
rect 519326 304718 519562 304954
rect 519646 304718 519882 304954
rect 519326 304398 519562 304634
rect 519646 304398 519882 304634
rect 519326 268718 519562 268954
rect 519646 268718 519882 268954
rect 519326 268398 519562 268634
rect 519646 268398 519882 268634
rect 519326 232718 519562 232954
rect 519646 232718 519882 232954
rect 519326 232398 519562 232634
rect 519646 232398 519882 232634
rect 519326 196718 519562 196954
rect 519646 196718 519882 196954
rect 519326 196398 519562 196634
rect 519646 196398 519882 196634
rect 519326 160718 519562 160954
rect 519646 160718 519882 160954
rect 519326 160398 519562 160634
rect 519646 160398 519882 160634
rect 519326 124718 519562 124954
rect 519646 124718 519882 124954
rect 519326 124398 519562 124634
rect 519646 124398 519882 124634
rect 519326 88718 519562 88954
rect 519646 88718 519882 88954
rect 519326 88398 519562 88634
rect 519646 88398 519882 88634
rect 519326 52718 519562 52954
rect 519646 52718 519882 52954
rect 519326 52398 519562 52634
rect 519646 52398 519882 52634
rect 519326 16718 519562 16954
rect 519646 16718 519882 16954
rect 519326 16398 519562 16634
rect 519646 16398 519882 16634
rect 519326 -3462 519562 -3226
rect 519646 -3462 519882 -3226
rect 519326 -3782 519562 -3546
rect 519646 -3782 519882 -3546
rect 523826 708442 524062 708678
rect 524146 708442 524382 708678
rect 523826 708122 524062 708358
rect 524146 708122 524382 708358
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -4422 524062 -4186
rect 524146 -4422 524382 -4186
rect 523826 -4742 524062 -4506
rect 524146 -4742 524382 -4506
rect 528326 709402 528562 709638
rect 528646 709402 528882 709638
rect 528326 709082 528562 709318
rect 528646 709082 528882 709318
rect 528326 673718 528562 673954
rect 528646 673718 528882 673954
rect 528326 673398 528562 673634
rect 528646 673398 528882 673634
rect 528326 637718 528562 637954
rect 528646 637718 528882 637954
rect 528326 637398 528562 637634
rect 528646 637398 528882 637634
rect 528326 601718 528562 601954
rect 528646 601718 528882 601954
rect 528326 601398 528562 601634
rect 528646 601398 528882 601634
rect 528326 565718 528562 565954
rect 528646 565718 528882 565954
rect 528326 565398 528562 565634
rect 528646 565398 528882 565634
rect 528326 529718 528562 529954
rect 528646 529718 528882 529954
rect 528326 529398 528562 529634
rect 528646 529398 528882 529634
rect 528326 493718 528562 493954
rect 528646 493718 528882 493954
rect 528326 493398 528562 493634
rect 528646 493398 528882 493634
rect 528326 457718 528562 457954
rect 528646 457718 528882 457954
rect 528326 457398 528562 457634
rect 528646 457398 528882 457634
rect 528326 421718 528562 421954
rect 528646 421718 528882 421954
rect 528326 421398 528562 421634
rect 528646 421398 528882 421634
rect 528326 385718 528562 385954
rect 528646 385718 528882 385954
rect 528326 385398 528562 385634
rect 528646 385398 528882 385634
rect 528326 349718 528562 349954
rect 528646 349718 528882 349954
rect 528326 349398 528562 349634
rect 528646 349398 528882 349634
rect 528326 313718 528562 313954
rect 528646 313718 528882 313954
rect 528326 313398 528562 313634
rect 528646 313398 528882 313634
rect 528326 277718 528562 277954
rect 528646 277718 528882 277954
rect 528326 277398 528562 277634
rect 528646 277398 528882 277634
rect 528326 241718 528562 241954
rect 528646 241718 528882 241954
rect 528326 241398 528562 241634
rect 528646 241398 528882 241634
rect 528326 205718 528562 205954
rect 528646 205718 528882 205954
rect 528326 205398 528562 205634
rect 528646 205398 528882 205634
rect 528326 169718 528562 169954
rect 528646 169718 528882 169954
rect 528326 169398 528562 169634
rect 528646 169398 528882 169634
rect 528326 133718 528562 133954
rect 528646 133718 528882 133954
rect 528326 133398 528562 133634
rect 528646 133398 528882 133634
rect 528326 97718 528562 97954
rect 528646 97718 528882 97954
rect 528326 97398 528562 97634
rect 528646 97398 528882 97634
rect 528326 61718 528562 61954
rect 528646 61718 528882 61954
rect 528326 61398 528562 61634
rect 528646 61398 528882 61634
rect 528326 25718 528562 25954
rect 528646 25718 528882 25954
rect 528326 25398 528562 25634
rect 528646 25398 528882 25634
rect 528326 -5382 528562 -5146
rect 528646 -5382 528882 -5146
rect 528326 -5702 528562 -5466
rect 528646 -5702 528882 -5466
rect 532826 710362 533062 710598
rect 533146 710362 533382 710598
rect 532826 710042 533062 710278
rect 533146 710042 533382 710278
rect 532826 678218 533062 678454
rect 533146 678218 533382 678454
rect 532826 677898 533062 678134
rect 533146 677898 533382 678134
rect 532826 642218 533062 642454
rect 533146 642218 533382 642454
rect 532826 641898 533062 642134
rect 533146 641898 533382 642134
rect 532826 606218 533062 606454
rect 533146 606218 533382 606454
rect 532826 605898 533062 606134
rect 533146 605898 533382 606134
rect 532826 570218 533062 570454
rect 533146 570218 533382 570454
rect 532826 569898 533062 570134
rect 533146 569898 533382 570134
rect 532826 534218 533062 534454
rect 533146 534218 533382 534454
rect 532826 533898 533062 534134
rect 533146 533898 533382 534134
rect 532826 498218 533062 498454
rect 533146 498218 533382 498454
rect 532826 497898 533062 498134
rect 533146 497898 533382 498134
rect 532826 462218 533062 462454
rect 533146 462218 533382 462454
rect 532826 461898 533062 462134
rect 533146 461898 533382 462134
rect 532826 426218 533062 426454
rect 533146 426218 533382 426454
rect 532826 425898 533062 426134
rect 533146 425898 533382 426134
rect 532826 390218 533062 390454
rect 533146 390218 533382 390454
rect 532826 389898 533062 390134
rect 533146 389898 533382 390134
rect 532826 354218 533062 354454
rect 533146 354218 533382 354454
rect 532826 353898 533062 354134
rect 533146 353898 533382 354134
rect 532826 318218 533062 318454
rect 533146 318218 533382 318454
rect 532826 317898 533062 318134
rect 533146 317898 533382 318134
rect 532826 282218 533062 282454
rect 533146 282218 533382 282454
rect 532826 281898 533062 282134
rect 533146 281898 533382 282134
rect 532826 246218 533062 246454
rect 533146 246218 533382 246454
rect 532826 245898 533062 246134
rect 533146 245898 533382 246134
rect 532826 210218 533062 210454
rect 533146 210218 533382 210454
rect 532826 209898 533062 210134
rect 533146 209898 533382 210134
rect 532826 174218 533062 174454
rect 533146 174218 533382 174454
rect 532826 173898 533062 174134
rect 533146 173898 533382 174134
rect 532826 138218 533062 138454
rect 533146 138218 533382 138454
rect 532826 137898 533062 138134
rect 533146 137898 533382 138134
rect 532826 102218 533062 102454
rect 533146 102218 533382 102454
rect 532826 101898 533062 102134
rect 533146 101898 533382 102134
rect 532826 66218 533062 66454
rect 533146 66218 533382 66454
rect 532826 65898 533062 66134
rect 533146 65898 533382 66134
rect 532826 30218 533062 30454
rect 533146 30218 533382 30454
rect 532826 29898 533062 30134
rect 533146 29898 533382 30134
rect 532826 -6342 533062 -6106
rect 533146 -6342 533382 -6106
rect 532826 -6662 533062 -6426
rect 533146 -6662 533382 -6426
rect 537326 711322 537562 711558
rect 537646 711322 537882 711558
rect 537326 711002 537562 711238
rect 537646 711002 537882 711238
rect 537326 682718 537562 682954
rect 537646 682718 537882 682954
rect 537326 682398 537562 682634
rect 537646 682398 537882 682634
rect 537326 646718 537562 646954
rect 537646 646718 537882 646954
rect 537326 646398 537562 646634
rect 537646 646398 537882 646634
rect 537326 610718 537562 610954
rect 537646 610718 537882 610954
rect 537326 610398 537562 610634
rect 537646 610398 537882 610634
rect 537326 574718 537562 574954
rect 537646 574718 537882 574954
rect 537326 574398 537562 574634
rect 537646 574398 537882 574634
rect 537326 538718 537562 538954
rect 537646 538718 537882 538954
rect 537326 538398 537562 538634
rect 537646 538398 537882 538634
rect 537326 502718 537562 502954
rect 537646 502718 537882 502954
rect 537326 502398 537562 502634
rect 537646 502398 537882 502634
rect 537326 466718 537562 466954
rect 537646 466718 537882 466954
rect 537326 466398 537562 466634
rect 537646 466398 537882 466634
rect 537326 430718 537562 430954
rect 537646 430718 537882 430954
rect 537326 430398 537562 430634
rect 537646 430398 537882 430634
rect 537326 394718 537562 394954
rect 537646 394718 537882 394954
rect 537326 394398 537562 394634
rect 537646 394398 537882 394634
rect 537326 358718 537562 358954
rect 537646 358718 537882 358954
rect 537326 358398 537562 358634
rect 537646 358398 537882 358634
rect 537326 322718 537562 322954
rect 537646 322718 537882 322954
rect 537326 322398 537562 322634
rect 537646 322398 537882 322634
rect 537326 286718 537562 286954
rect 537646 286718 537882 286954
rect 537326 286398 537562 286634
rect 537646 286398 537882 286634
rect 537326 250718 537562 250954
rect 537646 250718 537882 250954
rect 537326 250398 537562 250634
rect 537646 250398 537882 250634
rect 537326 214718 537562 214954
rect 537646 214718 537882 214954
rect 537326 214398 537562 214634
rect 537646 214398 537882 214634
rect 537326 178718 537562 178954
rect 537646 178718 537882 178954
rect 537326 178398 537562 178634
rect 537646 178398 537882 178634
rect 537326 142718 537562 142954
rect 537646 142718 537882 142954
rect 537326 142398 537562 142634
rect 537646 142398 537882 142634
rect 537326 106718 537562 106954
rect 537646 106718 537882 106954
rect 537326 106398 537562 106634
rect 537646 106398 537882 106634
rect 537326 70718 537562 70954
rect 537646 70718 537882 70954
rect 537326 70398 537562 70634
rect 537646 70398 537882 70634
rect 537326 34718 537562 34954
rect 537646 34718 537882 34954
rect 537326 34398 537562 34634
rect 537646 34398 537882 34634
rect 537326 -7302 537562 -7066
rect 537646 -7302 537882 -7066
rect 537326 -7622 537562 -7386
rect 537646 -7622 537882 -7386
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 546326 705562 546562 705798
rect 546646 705562 546882 705798
rect 546326 705242 546562 705478
rect 546646 705242 546882 705478
rect 546326 691718 546562 691954
rect 546646 691718 546882 691954
rect 546326 691398 546562 691634
rect 546646 691398 546882 691634
rect 546326 655718 546562 655954
rect 546646 655718 546882 655954
rect 546326 655398 546562 655634
rect 546646 655398 546882 655634
rect 546326 619718 546562 619954
rect 546646 619718 546882 619954
rect 546326 619398 546562 619634
rect 546646 619398 546882 619634
rect 546326 583718 546562 583954
rect 546646 583718 546882 583954
rect 546326 583398 546562 583634
rect 546646 583398 546882 583634
rect 546326 547718 546562 547954
rect 546646 547718 546882 547954
rect 546326 547398 546562 547634
rect 546646 547398 546882 547634
rect 546326 511718 546562 511954
rect 546646 511718 546882 511954
rect 546326 511398 546562 511634
rect 546646 511398 546882 511634
rect 546326 475718 546562 475954
rect 546646 475718 546882 475954
rect 546326 475398 546562 475634
rect 546646 475398 546882 475634
rect 546326 439718 546562 439954
rect 546646 439718 546882 439954
rect 546326 439398 546562 439634
rect 546646 439398 546882 439634
rect 546326 403718 546562 403954
rect 546646 403718 546882 403954
rect 546326 403398 546562 403634
rect 546646 403398 546882 403634
rect 546326 367718 546562 367954
rect 546646 367718 546882 367954
rect 546326 367398 546562 367634
rect 546646 367398 546882 367634
rect 546326 331718 546562 331954
rect 546646 331718 546882 331954
rect 546326 331398 546562 331634
rect 546646 331398 546882 331634
rect 546326 295718 546562 295954
rect 546646 295718 546882 295954
rect 546326 295398 546562 295634
rect 546646 295398 546882 295634
rect 546326 259718 546562 259954
rect 546646 259718 546882 259954
rect 546326 259398 546562 259634
rect 546646 259398 546882 259634
rect 546326 223718 546562 223954
rect 546646 223718 546882 223954
rect 546326 223398 546562 223634
rect 546646 223398 546882 223634
rect 546326 187718 546562 187954
rect 546646 187718 546882 187954
rect 546326 187398 546562 187634
rect 546646 187398 546882 187634
rect 546326 151718 546562 151954
rect 546646 151718 546882 151954
rect 546326 151398 546562 151634
rect 546646 151398 546882 151634
rect 546326 115718 546562 115954
rect 546646 115718 546882 115954
rect 546326 115398 546562 115634
rect 546646 115398 546882 115634
rect 546326 79718 546562 79954
rect 546646 79718 546882 79954
rect 546326 79398 546562 79634
rect 546646 79398 546882 79634
rect 546326 43718 546562 43954
rect 546646 43718 546882 43954
rect 546326 43398 546562 43634
rect 546646 43398 546882 43634
rect 546326 7718 546562 7954
rect 546646 7718 546882 7954
rect 546326 7398 546562 7634
rect 546646 7398 546882 7634
rect 546326 -1542 546562 -1306
rect 546646 -1542 546882 -1306
rect 546326 -1862 546562 -1626
rect 546646 -1862 546882 -1626
rect 550826 706522 551062 706758
rect 551146 706522 551382 706758
rect 550826 706202 551062 706438
rect 551146 706202 551382 706438
rect 550826 696218 551062 696454
rect 551146 696218 551382 696454
rect 550826 695898 551062 696134
rect 551146 695898 551382 696134
rect 550826 660218 551062 660454
rect 551146 660218 551382 660454
rect 550826 659898 551062 660134
rect 551146 659898 551382 660134
rect 550826 624218 551062 624454
rect 551146 624218 551382 624454
rect 550826 623898 551062 624134
rect 551146 623898 551382 624134
rect 550826 588218 551062 588454
rect 551146 588218 551382 588454
rect 550826 587898 551062 588134
rect 551146 587898 551382 588134
rect 550826 552218 551062 552454
rect 551146 552218 551382 552454
rect 550826 551898 551062 552134
rect 551146 551898 551382 552134
rect 550826 516218 551062 516454
rect 551146 516218 551382 516454
rect 550826 515898 551062 516134
rect 551146 515898 551382 516134
rect 550826 480218 551062 480454
rect 551146 480218 551382 480454
rect 550826 479898 551062 480134
rect 551146 479898 551382 480134
rect 550826 444218 551062 444454
rect 551146 444218 551382 444454
rect 550826 443898 551062 444134
rect 551146 443898 551382 444134
rect 550826 408218 551062 408454
rect 551146 408218 551382 408454
rect 550826 407898 551062 408134
rect 551146 407898 551382 408134
rect 550826 372218 551062 372454
rect 551146 372218 551382 372454
rect 550826 371898 551062 372134
rect 551146 371898 551382 372134
rect 550826 336218 551062 336454
rect 551146 336218 551382 336454
rect 550826 335898 551062 336134
rect 551146 335898 551382 336134
rect 550826 300218 551062 300454
rect 551146 300218 551382 300454
rect 550826 299898 551062 300134
rect 551146 299898 551382 300134
rect 550826 264218 551062 264454
rect 551146 264218 551382 264454
rect 550826 263898 551062 264134
rect 551146 263898 551382 264134
rect 550826 228218 551062 228454
rect 551146 228218 551382 228454
rect 550826 227898 551062 228134
rect 551146 227898 551382 228134
rect 550826 192218 551062 192454
rect 551146 192218 551382 192454
rect 550826 191898 551062 192134
rect 551146 191898 551382 192134
rect 550826 156218 551062 156454
rect 551146 156218 551382 156454
rect 550826 155898 551062 156134
rect 551146 155898 551382 156134
rect 550826 120218 551062 120454
rect 551146 120218 551382 120454
rect 550826 119898 551062 120134
rect 551146 119898 551382 120134
rect 550826 84218 551062 84454
rect 551146 84218 551382 84454
rect 550826 83898 551062 84134
rect 551146 83898 551382 84134
rect 550826 48218 551062 48454
rect 551146 48218 551382 48454
rect 550826 47898 551062 48134
rect 551146 47898 551382 48134
rect 550826 12218 551062 12454
rect 551146 12218 551382 12454
rect 550826 11898 551062 12134
rect 551146 11898 551382 12134
rect 550826 -2502 551062 -2266
rect 551146 -2502 551382 -2266
rect 550826 -2822 551062 -2586
rect 551146 -2822 551382 -2586
rect 555326 707482 555562 707718
rect 555646 707482 555882 707718
rect 555326 707162 555562 707398
rect 555646 707162 555882 707398
rect 555326 700718 555562 700954
rect 555646 700718 555882 700954
rect 555326 700398 555562 700634
rect 555646 700398 555882 700634
rect 555326 664718 555562 664954
rect 555646 664718 555882 664954
rect 555326 664398 555562 664634
rect 555646 664398 555882 664634
rect 555326 628718 555562 628954
rect 555646 628718 555882 628954
rect 555326 628398 555562 628634
rect 555646 628398 555882 628634
rect 555326 592718 555562 592954
rect 555646 592718 555882 592954
rect 555326 592398 555562 592634
rect 555646 592398 555882 592634
rect 555326 556718 555562 556954
rect 555646 556718 555882 556954
rect 555326 556398 555562 556634
rect 555646 556398 555882 556634
rect 555326 520718 555562 520954
rect 555646 520718 555882 520954
rect 555326 520398 555562 520634
rect 555646 520398 555882 520634
rect 555326 484718 555562 484954
rect 555646 484718 555882 484954
rect 555326 484398 555562 484634
rect 555646 484398 555882 484634
rect 555326 448718 555562 448954
rect 555646 448718 555882 448954
rect 555326 448398 555562 448634
rect 555646 448398 555882 448634
rect 555326 412718 555562 412954
rect 555646 412718 555882 412954
rect 555326 412398 555562 412634
rect 555646 412398 555882 412634
rect 555326 376718 555562 376954
rect 555646 376718 555882 376954
rect 555326 376398 555562 376634
rect 555646 376398 555882 376634
rect 555326 340718 555562 340954
rect 555646 340718 555882 340954
rect 555326 340398 555562 340634
rect 555646 340398 555882 340634
rect 555326 304718 555562 304954
rect 555646 304718 555882 304954
rect 555326 304398 555562 304634
rect 555646 304398 555882 304634
rect 555326 268718 555562 268954
rect 555646 268718 555882 268954
rect 555326 268398 555562 268634
rect 555646 268398 555882 268634
rect 555326 232718 555562 232954
rect 555646 232718 555882 232954
rect 555326 232398 555562 232634
rect 555646 232398 555882 232634
rect 555326 196718 555562 196954
rect 555646 196718 555882 196954
rect 555326 196398 555562 196634
rect 555646 196398 555882 196634
rect 555326 160718 555562 160954
rect 555646 160718 555882 160954
rect 555326 160398 555562 160634
rect 555646 160398 555882 160634
rect 555326 124718 555562 124954
rect 555646 124718 555882 124954
rect 555326 124398 555562 124634
rect 555646 124398 555882 124634
rect 555326 88718 555562 88954
rect 555646 88718 555882 88954
rect 555326 88398 555562 88634
rect 555646 88398 555882 88634
rect 555326 52718 555562 52954
rect 555646 52718 555882 52954
rect 555326 52398 555562 52634
rect 555646 52398 555882 52634
rect 555326 16718 555562 16954
rect 555646 16718 555882 16954
rect 555326 16398 555562 16634
rect 555646 16398 555882 16634
rect 555326 -3462 555562 -3226
rect 555646 -3462 555882 -3226
rect 555326 -3782 555562 -3546
rect 555646 -3782 555882 -3546
rect 559826 708442 560062 708678
rect 560146 708442 560382 708678
rect 559826 708122 560062 708358
rect 560146 708122 560382 708358
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -4422 560062 -4186
rect 560146 -4422 560382 -4186
rect 559826 -4742 560062 -4506
rect 560146 -4742 560382 -4506
rect 564326 709402 564562 709638
rect 564646 709402 564882 709638
rect 564326 709082 564562 709318
rect 564646 709082 564882 709318
rect 564326 673718 564562 673954
rect 564646 673718 564882 673954
rect 564326 673398 564562 673634
rect 564646 673398 564882 673634
rect 564326 637718 564562 637954
rect 564646 637718 564882 637954
rect 564326 637398 564562 637634
rect 564646 637398 564882 637634
rect 564326 601718 564562 601954
rect 564646 601718 564882 601954
rect 564326 601398 564562 601634
rect 564646 601398 564882 601634
rect 564326 565718 564562 565954
rect 564646 565718 564882 565954
rect 564326 565398 564562 565634
rect 564646 565398 564882 565634
rect 564326 529718 564562 529954
rect 564646 529718 564882 529954
rect 564326 529398 564562 529634
rect 564646 529398 564882 529634
rect 564326 493718 564562 493954
rect 564646 493718 564882 493954
rect 564326 493398 564562 493634
rect 564646 493398 564882 493634
rect 564326 457718 564562 457954
rect 564646 457718 564882 457954
rect 564326 457398 564562 457634
rect 564646 457398 564882 457634
rect 564326 421718 564562 421954
rect 564646 421718 564882 421954
rect 564326 421398 564562 421634
rect 564646 421398 564882 421634
rect 564326 385718 564562 385954
rect 564646 385718 564882 385954
rect 564326 385398 564562 385634
rect 564646 385398 564882 385634
rect 564326 349718 564562 349954
rect 564646 349718 564882 349954
rect 564326 349398 564562 349634
rect 564646 349398 564882 349634
rect 564326 313718 564562 313954
rect 564646 313718 564882 313954
rect 564326 313398 564562 313634
rect 564646 313398 564882 313634
rect 564326 277718 564562 277954
rect 564646 277718 564882 277954
rect 564326 277398 564562 277634
rect 564646 277398 564882 277634
rect 564326 241718 564562 241954
rect 564646 241718 564882 241954
rect 564326 241398 564562 241634
rect 564646 241398 564882 241634
rect 564326 205718 564562 205954
rect 564646 205718 564882 205954
rect 564326 205398 564562 205634
rect 564646 205398 564882 205634
rect 564326 169718 564562 169954
rect 564646 169718 564882 169954
rect 564326 169398 564562 169634
rect 564646 169398 564882 169634
rect 564326 133718 564562 133954
rect 564646 133718 564882 133954
rect 564326 133398 564562 133634
rect 564646 133398 564882 133634
rect 564326 97718 564562 97954
rect 564646 97718 564882 97954
rect 564326 97398 564562 97634
rect 564646 97398 564882 97634
rect 564326 61718 564562 61954
rect 564646 61718 564882 61954
rect 564326 61398 564562 61634
rect 564646 61398 564882 61634
rect 564326 25718 564562 25954
rect 564646 25718 564882 25954
rect 564326 25398 564562 25634
rect 564646 25398 564882 25634
rect 564326 -5382 564562 -5146
rect 564646 -5382 564882 -5146
rect 564326 -5702 564562 -5466
rect 564646 -5702 564882 -5466
rect 568826 710362 569062 710598
rect 569146 710362 569382 710598
rect 568826 710042 569062 710278
rect 569146 710042 569382 710278
rect 568826 678218 569062 678454
rect 569146 678218 569382 678454
rect 568826 677898 569062 678134
rect 569146 677898 569382 678134
rect 568826 642218 569062 642454
rect 569146 642218 569382 642454
rect 568826 641898 569062 642134
rect 569146 641898 569382 642134
rect 568826 606218 569062 606454
rect 569146 606218 569382 606454
rect 568826 605898 569062 606134
rect 569146 605898 569382 606134
rect 568826 570218 569062 570454
rect 569146 570218 569382 570454
rect 568826 569898 569062 570134
rect 569146 569898 569382 570134
rect 568826 534218 569062 534454
rect 569146 534218 569382 534454
rect 568826 533898 569062 534134
rect 569146 533898 569382 534134
rect 568826 498218 569062 498454
rect 569146 498218 569382 498454
rect 568826 497898 569062 498134
rect 569146 497898 569382 498134
rect 568826 462218 569062 462454
rect 569146 462218 569382 462454
rect 568826 461898 569062 462134
rect 569146 461898 569382 462134
rect 568826 426218 569062 426454
rect 569146 426218 569382 426454
rect 568826 425898 569062 426134
rect 569146 425898 569382 426134
rect 568826 390218 569062 390454
rect 569146 390218 569382 390454
rect 568826 389898 569062 390134
rect 569146 389898 569382 390134
rect 568826 354218 569062 354454
rect 569146 354218 569382 354454
rect 568826 353898 569062 354134
rect 569146 353898 569382 354134
rect 568826 318218 569062 318454
rect 569146 318218 569382 318454
rect 568826 317898 569062 318134
rect 569146 317898 569382 318134
rect 568826 282218 569062 282454
rect 569146 282218 569382 282454
rect 568826 281898 569062 282134
rect 569146 281898 569382 282134
rect 568826 246218 569062 246454
rect 569146 246218 569382 246454
rect 568826 245898 569062 246134
rect 569146 245898 569382 246134
rect 568826 210218 569062 210454
rect 569146 210218 569382 210454
rect 568826 209898 569062 210134
rect 569146 209898 569382 210134
rect 568826 174218 569062 174454
rect 569146 174218 569382 174454
rect 568826 173898 569062 174134
rect 569146 173898 569382 174134
rect 568826 138218 569062 138454
rect 569146 138218 569382 138454
rect 568826 137898 569062 138134
rect 569146 137898 569382 138134
rect 568826 102218 569062 102454
rect 569146 102218 569382 102454
rect 568826 101898 569062 102134
rect 569146 101898 569382 102134
rect 568826 66218 569062 66454
rect 569146 66218 569382 66454
rect 568826 65898 569062 66134
rect 569146 65898 569382 66134
rect 568826 30218 569062 30454
rect 569146 30218 569382 30454
rect 568826 29898 569062 30134
rect 569146 29898 569382 30134
rect 568826 -6342 569062 -6106
rect 569146 -6342 569382 -6106
rect 568826 -6662 569062 -6426
rect 569146 -6662 569382 -6426
rect 573326 711322 573562 711558
rect 573646 711322 573882 711558
rect 573326 711002 573562 711238
rect 573646 711002 573882 711238
rect 573326 682718 573562 682954
rect 573646 682718 573882 682954
rect 573326 682398 573562 682634
rect 573646 682398 573882 682634
rect 573326 646718 573562 646954
rect 573646 646718 573882 646954
rect 573326 646398 573562 646634
rect 573646 646398 573882 646634
rect 573326 610718 573562 610954
rect 573646 610718 573882 610954
rect 573326 610398 573562 610634
rect 573646 610398 573882 610634
rect 573326 574718 573562 574954
rect 573646 574718 573882 574954
rect 573326 574398 573562 574634
rect 573646 574398 573882 574634
rect 573326 538718 573562 538954
rect 573646 538718 573882 538954
rect 573326 538398 573562 538634
rect 573646 538398 573882 538634
rect 573326 502718 573562 502954
rect 573646 502718 573882 502954
rect 573326 502398 573562 502634
rect 573646 502398 573882 502634
rect 573326 466718 573562 466954
rect 573646 466718 573882 466954
rect 573326 466398 573562 466634
rect 573646 466398 573882 466634
rect 573326 430718 573562 430954
rect 573646 430718 573882 430954
rect 573326 430398 573562 430634
rect 573646 430398 573882 430634
rect 573326 394718 573562 394954
rect 573646 394718 573882 394954
rect 573326 394398 573562 394634
rect 573646 394398 573882 394634
rect 573326 358718 573562 358954
rect 573646 358718 573882 358954
rect 573326 358398 573562 358634
rect 573646 358398 573882 358634
rect 573326 322718 573562 322954
rect 573646 322718 573882 322954
rect 573326 322398 573562 322634
rect 573646 322398 573882 322634
rect 573326 286718 573562 286954
rect 573646 286718 573882 286954
rect 573326 286398 573562 286634
rect 573646 286398 573882 286634
rect 573326 250718 573562 250954
rect 573646 250718 573882 250954
rect 573326 250398 573562 250634
rect 573646 250398 573882 250634
rect 573326 214718 573562 214954
rect 573646 214718 573882 214954
rect 573326 214398 573562 214634
rect 573646 214398 573882 214634
rect 573326 178718 573562 178954
rect 573646 178718 573882 178954
rect 573326 178398 573562 178634
rect 573646 178398 573882 178634
rect 573326 142718 573562 142954
rect 573646 142718 573882 142954
rect 573326 142398 573562 142634
rect 573646 142398 573882 142634
rect 573326 106718 573562 106954
rect 573646 106718 573882 106954
rect 573326 106398 573562 106634
rect 573646 106398 573882 106634
rect 573326 70718 573562 70954
rect 573646 70718 573882 70954
rect 573326 70398 573562 70634
rect 573646 70398 573882 70634
rect 573326 34718 573562 34954
rect 573646 34718 573882 34954
rect 573326 34398 573562 34634
rect 573646 34398 573882 34634
rect 573326 -7302 573562 -7066
rect 573646 -7302 573882 -7066
rect 573326 -7622 573562 -7386
rect 573646 -7622 573882 -7386
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 582326 705562 582562 705798
rect 582646 705562 582882 705798
rect 582326 705242 582562 705478
rect 582646 705242 582882 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 582326 691718 582562 691954
rect 582646 691718 582882 691954
rect 582326 691398 582562 691634
rect 582646 691398 582882 691634
rect 582326 655718 582562 655954
rect 582646 655718 582882 655954
rect 582326 655398 582562 655634
rect 582646 655398 582882 655634
rect 582326 619718 582562 619954
rect 582646 619718 582882 619954
rect 582326 619398 582562 619634
rect 582646 619398 582882 619634
rect 582326 583718 582562 583954
rect 582646 583718 582882 583954
rect 582326 583398 582562 583634
rect 582646 583398 582882 583634
rect 582326 547718 582562 547954
rect 582646 547718 582882 547954
rect 582326 547398 582562 547634
rect 582646 547398 582882 547634
rect 582326 511718 582562 511954
rect 582646 511718 582882 511954
rect 582326 511398 582562 511634
rect 582646 511398 582882 511634
rect 582326 475718 582562 475954
rect 582646 475718 582882 475954
rect 582326 475398 582562 475634
rect 582646 475398 582882 475634
rect 582326 439718 582562 439954
rect 582646 439718 582882 439954
rect 582326 439398 582562 439634
rect 582646 439398 582882 439634
rect 582326 403718 582562 403954
rect 582646 403718 582882 403954
rect 582326 403398 582562 403634
rect 582646 403398 582882 403634
rect 582326 367718 582562 367954
rect 582646 367718 582882 367954
rect 582326 367398 582562 367634
rect 582646 367398 582882 367634
rect 582326 331718 582562 331954
rect 582646 331718 582882 331954
rect 582326 331398 582562 331634
rect 582646 331398 582882 331634
rect 582326 295718 582562 295954
rect 582646 295718 582882 295954
rect 582326 295398 582562 295634
rect 582646 295398 582882 295634
rect 582326 259718 582562 259954
rect 582646 259718 582882 259954
rect 582326 259398 582562 259634
rect 582646 259398 582882 259634
rect 582326 223718 582562 223954
rect 582646 223718 582882 223954
rect 582326 223398 582562 223634
rect 582646 223398 582882 223634
rect 582326 187718 582562 187954
rect 582646 187718 582882 187954
rect 582326 187398 582562 187634
rect 582646 187398 582882 187634
rect 582326 151718 582562 151954
rect 582646 151718 582882 151954
rect 582326 151398 582562 151634
rect 582646 151398 582882 151634
rect 582326 115718 582562 115954
rect 582646 115718 582882 115954
rect 582326 115398 582562 115634
rect 582646 115398 582882 115634
rect 582326 79718 582562 79954
rect 582646 79718 582882 79954
rect 582326 79398 582562 79634
rect 582646 79398 582882 79634
rect 582326 43718 582562 43954
rect 582646 43718 582882 43954
rect 582326 43398 582562 43634
rect 582646 43398 582882 43634
rect 582326 7718 582562 7954
rect 582646 7718 582882 7954
rect 582326 7398 582562 7634
rect 582646 7398 582882 7634
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 691718 586538 691954
rect 586622 691718 586858 691954
rect 586302 691398 586538 691634
rect 586622 691398 586858 691634
rect 586302 655718 586538 655954
rect 586622 655718 586858 655954
rect 586302 655398 586538 655634
rect 586622 655398 586858 655634
rect 586302 619718 586538 619954
rect 586622 619718 586858 619954
rect 586302 619398 586538 619634
rect 586622 619398 586858 619634
rect 586302 583718 586538 583954
rect 586622 583718 586858 583954
rect 586302 583398 586538 583634
rect 586622 583398 586858 583634
rect 586302 547718 586538 547954
rect 586622 547718 586858 547954
rect 586302 547398 586538 547634
rect 586622 547398 586858 547634
rect 586302 511718 586538 511954
rect 586622 511718 586858 511954
rect 586302 511398 586538 511634
rect 586622 511398 586858 511634
rect 586302 475718 586538 475954
rect 586622 475718 586858 475954
rect 586302 475398 586538 475634
rect 586622 475398 586858 475634
rect 586302 439718 586538 439954
rect 586622 439718 586858 439954
rect 586302 439398 586538 439634
rect 586622 439398 586858 439634
rect 586302 403718 586538 403954
rect 586622 403718 586858 403954
rect 586302 403398 586538 403634
rect 586622 403398 586858 403634
rect 586302 367718 586538 367954
rect 586622 367718 586858 367954
rect 586302 367398 586538 367634
rect 586622 367398 586858 367634
rect 586302 331718 586538 331954
rect 586622 331718 586858 331954
rect 586302 331398 586538 331634
rect 586622 331398 586858 331634
rect 586302 295718 586538 295954
rect 586622 295718 586858 295954
rect 586302 295398 586538 295634
rect 586622 295398 586858 295634
rect 586302 259718 586538 259954
rect 586622 259718 586858 259954
rect 586302 259398 586538 259634
rect 586622 259398 586858 259634
rect 586302 223718 586538 223954
rect 586622 223718 586858 223954
rect 586302 223398 586538 223634
rect 586622 223398 586858 223634
rect 586302 187718 586538 187954
rect 586622 187718 586858 187954
rect 586302 187398 586538 187634
rect 586622 187398 586858 187634
rect 586302 151718 586538 151954
rect 586622 151718 586858 151954
rect 586302 151398 586538 151634
rect 586622 151398 586858 151634
rect 586302 115718 586538 115954
rect 586622 115718 586858 115954
rect 586302 115398 586538 115634
rect 586622 115398 586858 115634
rect 586302 79718 586538 79954
rect 586622 79718 586858 79954
rect 586302 79398 586538 79634
rect 586622 79398 586858 79634
rect 586302 43718 586538 43954
rect 586622 43718 586858 43954
rect 586302 43398 586538 43634
rect 586622 43398 586858 43634
rect 586302 7718 586538 7954
rect 586622 7718 586858 7954
rect 586302 7398 586538 7634
rect 586622 7398 586858 7634
rect 582326 -1542 582562 -1306
rect 582646 -1542 582882 -1306
rect 582326 -1862 582562 -1626
rect 582646 -1862 582882 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 696218 587498 696454
rect 587582 696218 587818 696454
rect 587262 695898 587498 696134
rect 587582 695898 587818 696134
rect 587262 660218 587498 660454
rect 587582 660218 587818 660454
rect 587262 659898 587498 660134
rect 587582 659898 587818 660134
rect 587262 624218 587498 624454
rect 587582 624218 587818 624454
rect 587262 623898 587498 624134
rect 587582 623898 587818 624134
rect 587262 588218 587498 588454
rect 587582 588218 587818 588454
rect 587262 587898 587498 588134
rect 587582 587898 587818 588134
rect 587262 552218 587498 552454
rect 587582 552218 587818 552454
rect 587262 551898 587498 552134
rect 587582 551898 587818 552134
rect 587262 516218 587498 516454
rect 587582 516218 587818 516454
rect 587262 515898 587498 516134
rect 587582 515898 587818 516134
rect 587262 480218 587498 480454
rect 587582 480218 587818 480454
rect 587262 479898 587498 480134
rect 587582 479898 587818 480134
rect 587262 444218 587498 444454
rect 587582 444218 587818 444454
rect 587262 443898 587498 444134
rect 587582 443898 587818 444134
rect 587262 408218 587498 408454
rect 587582 408218 587818 408454
rect 587262 407898 587498 408134
rect 587582 407898 587818 408134
rect 587262 372218 587498 372454
rect 587582 372218 587818 372454
rect 587262 371898 587498 372134
rect 587582 371898 587818 372134
rect 587262 336218 587498 336454
rect 587582 336218 587818 336454
rect 587262 335898 587498 336134
rect 587582 335898 587818 336134
rect 587262 300218 587498 300454
rect 587582 300218 587818 300454
rect 587262 299898 587498 300134
rect 587582 299898 587818 300134
rect 587262 264218 587498 264454
rect 587582 264218 587818 264454
rect 587262 263898 587498 264134
rect 587582 263898 587818 264134
rect 587262 228218 587498 228454
rect 587582 228218 587818 228454
rect 587262 227898 587498 228134
rect 587582 227898 587818 228134
rect 587262 192218 587498 192454
rect 587582 192218 587818 192454
rect 587262 191898 587498 192134
rect 587582 191898 587818 192134
rect 587262 156218 587498 156454
rect 587582 156218 587818 156454
rect 587262 155898 587498 156134
rect 587582 155898 587818 156134
rect 587262 120218 587498 120454
rect 587582 120218 587818 120454
rect 587262 119898 587498 120134
rect 587582 119898 587818 120134
rect 587262 84218 587498 84454
rect 587582 84218 587818 84454
rect 587262 83898 587498 84134
rect 587582 83898 587818 84134
rect 587262 48218 587498 48454
rect 587582 48218 587818 48454
rect 587262 47898 587498 48134
rect 587582 47898 587818 48134
rect 587262 12218 587498 12454
rect 587582 12218 587818 12454
rect 587262 11898 587498 12134
rect 587582 11898 587818 12134
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 700718 588458 700954
rect 588542 700718 588778 700954
rect 588222 700398 588458 700634
rect 588542 700398 588778 700634
rect 588222 664718 588458 664954
rect 588542 664718 588778 664954
rect 588222 664398 588458 664634
rect 588542 664398 588778 664634
rect 588222 628718 588458 628954
rect 588542 628718 588778 628954
rect 588222 628398 588458 628634
rect 588542 628398 588778 628634
rect 588222 592718 588458 592954
rect 588542 592718 588778 592954
rect 588222 592398 588458 592634
rect 588542 592398 588778 592634
rect 588222 556718 588458 556954
rect 588542 556718 588778 556954
rect 588222 556398 588458 556634
rect 588542 556398 588778 556634
rect 588222 520718 588458 520954
rect 588542 520718 588778 520954
rect 588222 520398 588458 520634
rect 588542 520398 588778 520634
rect 588222 484718 588458 484954
rect 588542 484718 588778 484954
rect 588222 484398 588458 484634
rect 588542 484398 588778 484634
rect 588222 448718 588458 448954
rect 588542 448718 588778 448954
rect 588222 448398 588458 448634
rect 588542 448398 588778 448634
rect 588222 412718 588458 412954
rect 588542 412718 588778 412954
rect 588222 412398 588458 412634
rect 588542 412398 588778 412634
rect 588222 376718 588458 376954
rect 588542 376718 588778 376954
rect 588222 376398 588458 376634
rect 588542 376398 588778 376634
rect 588222 340718 588458 340954
rect 588542 340718 588778 340954
rect 588222 340398 588458 340634
rect 588542 340398 588778 340634
rect 588222 304718 588458 304954
rect 588542 304718 588778 304954
rect 588222 304398 588458 304634
rect 588542 304398 588778 304634
rect 588222 268718 588458 268954
rect 588542 268718 588778 268954
rect 588222 268398 588458 268634
rect 588542 268398 588778 268634
rect 588222 232718 588458 232954
rect 588542 232718 588778 232954
rect 588222 232398 588458 232634
rect 588542 232398 588778 232634
rect 588222 196718 588458 196954
rect 588542 196718 588778 196954
rect 588222 196398 588458 196634
rect 588542 196398 588778 196634
rect 588222 160718 588458 160954
rect 588542 160718 588778 160954
rect 588222 160398 588458 160634
rect 588542 160398 588778 160634
rect 588222 124718 588458 124954
rect 588542 124718 588778 124954
rect 588222 124398 588458 124634
rect 588542 124398 588778 124634
rect 588222 88718 588458 88954
rect 588542 88718 588778 88954
rect 588222 88398 588458 88634
rect 588542 88398 588778 88634
rect 588222 52718 588458 52954
rect 588542 52718 588778 52954
rect 588222 52398 588458 52634
rect 588542 52398 588778 52634
rect 588222 16718 588458 16954
rect 588542 16718 588778 16954
rect 588222 16398 588458 16634
rect 588542 16398 588778 16634
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 669218 589418 669454
rect 589502 669218 589738 669454
rect 589182 668898 589418 669134
rect 589502 668898 589738 669134
rect 589182 633218 589418 633454
rect 589502 633218 589738 633454
rect 589182 632898 589418 633134
rect 589502 632898 589738 633134
rect 589182 597218 589418 597454
rect 589502 597218 589738 597454
rect 589182 596898 589418 597134
rect 589502 596898 589738 597134
rect 589182 561218 589418 561454
rect 589502 561218 589738 561454
rect 589182 560898 589418 561134
rect 589502 560898 589738 561134
rect 589182 525218 589418 525454
rect 589502 525218 589738 525454
rect 589182 524898 589418 525134
rect 589502 524898 589738 525134
rect 589182 489218 589418 489454
rect 589502 489218 589738 489454
rect 589182 488898 589418 489134
rect 589502 488898 589738 489134
rect 589182 453218 589418 453454
rect 589502 453218 589738 453454
rect 589182 452898 589418 453134
rect 589502 452898 589738 453134
rect 589182 417218 589418 417454
rect 589502 417218 589738 417454
rect 589182 416898 589418 417134
rect 589502 416898 589738 417134
rect 589182 381218 589418 381454
rect 589502 381218 589738 381454
rect 589182 380898 589418 381134
rect 589502 380898 589738 381134
rect 589182 345218 589418 345454
rect 589502 345218 589738 345454
rect 589182 344898 589418 345134
rect 589502 344898 589738 345134
rect 589182 309218 589418 309454
rect 589502 309218 589738 309454
rect 589182 308898 589418 309134
rect 589502 308898 589738 309134
rect 589182 273218 589418 273454
rect 589502 273218 589738 273454
rect 589182 272898 589418 273134
rect 589502 272898 589738 273134
rect 589182 237218 589418 237454
rect 589502 237218 589738 237454
rect 589182 236898 589418 237134
rect 589502 236898 589738 237134
rect 589182 201218 589418 201454
rect 589502 201218 589738 201454
rect 589182 200898 589418 201134
rect 589502 200898 589738 201134
rect 589182 165218 589418 165454
rect 589502 165218 589738 165454
rect 589182 164898 589418 165134
rect 589502 164898 589738 165134
rect 589182 129218 589418 129454
rect 589502 129218 589738 129454
rect 589182 128898 589418 129134
rect 589502 128898 589738 129134
rect 589182 93218 589418 93454
rect 589502 93218 589738 93454
rect 589182 92898 589418 93134
rect 589502 92898 589738 93134
rect 589182 57218 589418 57454
rect 589502 57218 589738 57454
rect 589182 56898 589418 57134
rect 589502 56898 589738 57134
rect 589182 21218 589418 21454
rect 589502 21218 589738 21454
rect 589182 20898 589418 21134
rect 589502 20898 589738 21134
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 673718 590378 673954
rect 590462 673718 590698 673954
rect 590142 673398 590378 673634
rect 590462 673398 590698 673634
rect 590142 637718 590378 637954
rect 590462 637718 590698 637954
rect 590142 637398 590378 637634
rect 590462 637398 590698 637634
rect 590142 601718 590378 601954
rect 590462 601718 590698 601954
rect 590142 601398 590378 601634
rect 590462 601398 590698 601634
rect 590142 565718 590378 565954
rect 590462 565718 590698 565954
rect 590142 565398 590378 565634
rect 590462 565398 590698 565634
rect 590142 529718 590378 529954
rect 590462 529718 590698 529954
rect 590142 529398 590378 529634
rect 590462 529398 590698 529634
rect 590142 493718 590378 493954
rect 590462 493718 590698 493954
rect 590142 493398 590378 493634
rect 590462 493398 590698 493634
rect 590142 457718 590378 457954
rect 590462 457718 590698 457954
rect 590142 457398 590378 457634
rect 590462 457398 590698 457634
rect 590142 421718 590378 421954
rect 590462 421718 590698 421954
rect 590142 421398 590378 421634
rect 590462 421398 590698 421634
rect 590142 385718 590378 385954
rect 590462 385718 590698 385954
rect 590142 385398 590378 385634
rect 590462 385398 590698 385634
rect 590142 349718 590378 349954
rect 590462 349718 590698 349954
rect 590142 349398 590378 349634
rect 590462 349398 590698 349634
rect 590142 313718 590378 313954
rect 590462 313718 590698 313954
rect 590142 313398 590378 313634
rect 590462 313398 590698 313634
rect 590142 277718 590378 277954
rect 590462 277718 590698 277954
rect 590142 277398 590378 277634
rect 590462 277398 590698 277634
rect 590142 241718 590378 241954
rect 590462 241718 590698 241954
rect 590142 241398 590378 241634
rect 590462 241398 590698 241634
rect 590142 205718 590378 205954
rect 590462 205718 590698 205954
rect 590142 205398 590378 205634
rect 590462 205398 590698 205634
rect 590142 169718 590378 169954
rect 590462 169718 590698 169954
rect 590142 169398 590378 169634
rect 590462 169398 590698 169634
rect 590142 133718 590378 133954
rect 590462 133718 590698 133954
rect 590142 133398 590378 133634
rect 590462 133398 590698 133634
rect 590142 97718 590378 97954
rect 590462 97718 590698 97954
rect 590142 97398 590378 97634
rect 590462 97398 590698 97634
rect 590142 61718 590378 61954
rect 590462 61718 590698 61954
rect 590142 61398 590378 61634
rect 590462 61398 590698 61634
rect 590142 25718 590378 25954
rect 590462 25718 590698 25954
rect 590142 25398 590378 25634
rect 590462 25398 590698 25634
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 678218 591338 678454
rect 591422 678218 591658 678454
rect 591102 677898 591338 678134
rect 591422 677898 591658 678134
rect 591102 642218 591338 642454
rect 591422 642218 591658 642454
rect 591102 641898 591338 642134
rect 591422 641898 591658 642134
rect 591102 606218 591338 606454
rect 591422 606218 591658 606454
rect 591102 605898 591338 606134
rect 591422 605898 591658 606134
rect 591102 570218 591338 570454
rect 591422 570218 591658 570454
rect 591102 569898 591338 570134
rect 591422 569898 591658 570134
rect 591102 534218 591338 534454
rect 591422 534218 591658 534454
rect 591102 533898 591338 534134
rect 591422 533898 591658 534134
rect 591102 498218 591338 498454
rect 591422 498218 591658 498454
rect 591102 497898 591338 498134
rect 591422 497898 591658 498134
rect 591102 462218 591338 462454
rect 591422 462218 591658 462454
rect 591102 461898 591338 462134
rect 591422 461898 591658 462134
rect 591102 426218 591338 426454
rect 591422 426218 591658 426454
rect 591102 425898 591338 426134
rect 591422 425898 591658 426134
rect 591102 390218 591338 390454
rect 591422 390218 591658 390454
rect 591102 389898 591338 390134
rect 591422 389898 591658 390134
rect 591102 354218 591338 354454
rect 591422 354218 591658 354454
rect 591102 353898 591338 354134
rect 591422 353898 591658 354134
rect 591102 318218 591338 318454
rect 591422 318218 591658 318454
rect 591102 317898 591338 318134
rect 591422 317898 591658 318134
rect 591102 282218 591338 282454
rect 591422 282218 591658 282454
rect 591102 281898 591338 282134
rect 591422 281898 591658 282134
rect 591102 246218 591338 246454
rect 591422 246218 591658 246454
rect 591102 245898 591338 246134
rect 591422 245898 591658 246134
rect 591102 210218 591338 210454
rect 591422 210218 591658 210454
rect 591102 209898 591338 210134
rect 591422 209898 591658 210134
rect 591102 174218 591338 174454
rect 591422 174218 591658 174454
rect 591102 173898 591338 174134
rect 591422 173898 591658 174134
rect 591102 138218 591338 138454
rect 591422 138218 591658 138454
rect 591102 137898 591338 138134
rect 591422 137898 591658 138134
rect 591102 102218 591338 102454
rect 591422 102218 591658 102454
rect 591102 101898 591338 102134
rect 591422 101898 591658 102134
rect 591102 66218 591338 66454
rect 591422 66218 591658 66454
rect 591102 65898 591338 66134
rect 591422 65898 591658 66134
rect 591102 30218 591338 30454
rect 591422 30218 591658 30454
rect 591102 29898 591338 30134
rect 591422 29898 591658 30134
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 682718 592298 682954
rect 592382 682718 592618 682954
rect 592062 682398 592298 682634
rect 592382 682398 592618 682634
rect 592062 646718 592298 646954
rect 592382 646718 592618 646954
rect 592062 646398 592298 646634
rect 592382 646398 592618 646634
rect 592062 610718 592298 610954
rect 592382 610718 592618 610954
rect 592062 610398 592298 610634
rect 592382 610398 592618 610634
rect 592062 574718 592298 574954
rect 592382 574718 592618 574954
rect 592062 574398 592298 574634
rect 592382 574398 592618 574634
rect 592062 538718 592298 538954
rect 592382 538718 592618 538954
rect 592062 538398 592298 538634
rect 592382 538398 592618 538634
rect 592062 502718 592298 502954
rect 592382 502718 592618 502954
rect 592062 502398 592298 502634
rect 592382 502398 592618 502634
rect 592062 466718 592298 466954
rect 592382 466718 592618 466954
rect 592062 466398 592298 466634
rect 592382 466398 592618 466634
rect 592062 430718 592298 430954
rect 592382 430718 592618 430954
rect 592062 430398 592298 430634
rect 592382 430398 592618 430634
rect 592062 394718 592298 394954
rect 592382 394718 592618 394954
rect 592062 394398 592298 394634
rect 592382 394398 592618 394634
rect 592062 358718 592298 358954
rect 592382 358718 592618 358954
rect 592062 358398 592298 358634
rect 592382 358398 592618 358634
rect 592062 322718 592298 322954
rect 592382 322718 592618 322954
rect 592062 322398 592298 322634
rect 592382 322398 592618 322634
rect 592062 286718 592298 286954
rect 592382 286718 592618 286954
rect 592062 286398 592298 286634
rect 592382 286398 592618 286634
rect 592062 250718 592298 250954
rect 592382 250718 592618 250954
rect 592062 250398 592298 250634
rect 592382 250398 592618 250634
rect 592062 214718 592298 214954
rect 592382 214718 592618 214954
rect 592062 214398 592298 214634
rect 592382 214398 592618 214634
rect 592062 178718 592298 178954
rect 592382 178718 592618 178954
rect 592062 178398 592298 178634
rect 592382 178398 592618 178634
rect 592062 142718 592298 142954
rect 592382 142718 592618 142954
rect 592062 142398 592298 142634
rect 592382 142398 592618 142634
rect 592062 106718 592298 106954
rect 592382 106718 592618 106954
rect 592062 106398 592298 106634
rect 592382 106398 592618 106634
rect 592062 70718 592298 70954
rect 592382 70718 592618 70954
rect 592062 70398 592298 70634
rect 592382 70398 592618 70634
rect 592062 34718 592298 34954
rect 592382 34718 592618 34954
rect 592062 34398 592298 34634
rect 592382 34398 592618 34634
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 700954 592650 700986
rect -8726 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 592650 700954
rect -8726 700634 592650 700718
rect -8726 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 592650 700634
rect -8726 700366 592650 700398
rect -8726 696454 592650 696486
rect -8726 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 592650 696454
rect -8726 696134 592650 696218
rect -8726 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 592650 696134
rect -8726 695866 592650 695898
rect -8726 691954 592650 691986
rect -8726 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 592650 691954
rect -8726 691634 592650 691718
rect -8726 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 592650 691634
rect -8726 691366 592650 691398
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 682954 592650 682986
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect -8726 682634 592650 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect -8726 682366 592650 682398
rect -8726 678454 592650 678486
rect -8726 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 592650 678454
rect -8726 678134 592650 678218
rect -8726 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 592650 678134
rect -8726 677866 592650 677898
rect -8726 673954 592650 673986
rect -8726 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 592650 673954
rect -8726 673634 592650 673718
rect -8726 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 592650 673634
rect -8726 673366 592650 673398
rect -8726 669454 592650 669486
rect -8726 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 592650 669454
rect -8726 669134 592650 669218
rect -8726 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 592650 669134
rect -8726 668866 592650 668898
rect -8726 664954 592650 664986
rect -8726 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 592650 664954
rect -8726 664634 592650 664718
rect -8726 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 592650 664634
rect -8726 664366 592650 664398
rect -8726 660454 592650 660486
rect -8726 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 592650 660454
rect -8726 660134 592650 660218
rect -8726 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 592650 660134
rect -8726 659866 592650 659898
rect -8726 655954 592650 655986
rect -8726 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 592650 655954
rect -8726 655634 592650 655718
rect -8726 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 592650 655634
rect -8726 655366 592650 655398
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 646954 592650 646986
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect -8726 646634 592650 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect -8726 646366 592650 646398
rect -8726 642454 592650 642486
rect -8726 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 592650 642454
rect -8726 642134 592650 642218
rect -8726 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 592650 642134
rect -8726 641866 592650 641898
rect -8726 637954 592650 637986
rect -8726 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 592650 637954
rect -8726 637634 592650 637718
rect -8726 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 592650 637634
rect -8726 637366 592650 637398
rect -8726 633454 592650 633486
rect -8726 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 592650 633454
rect -8726 633134 592650 633218
rect -8726 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 592650 633134
rect -8726 632866 592650 632898
rect -8726 628954 592650 628986
rect -8726 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 592650 628954
rect -8726 628634 592650 628718
rect -8726 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 592650 628634
rect -8726 628366 592650 628398
rect -8726 624454 592650 624486
rect -8726 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 592650 624454
rect -8726 624134 592650 624218
rect -8726 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 592650 624134
rect -8726 623866 592650 623898
rect -8726 619954 592650 619986
rect -8726 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 592650 619954
rect -8726 619634 592650 619718
rect -8726 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 592650 619634
rect -8726 619366 592650 619398
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 610954 592650 610986
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect -8726 610634 592650 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect -8726 610366 592650 610398
rect -8726 606454 592650 606486
rect -8726 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 592650 606454
rect -8726 606134 592650 606218
rect -8726 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 592650 606134
rect -8726 605866 592650 605898
rect -8726 601954 592650 601986
rect -8726 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 592650 601954
rect -8726 601634 592650 601718
rect -8726 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 592650 601634
rect -8726 601366 592650 601398
rect -8726 597454 592650 597486
rect -8726 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 592650 597454
rect -8726 597134 592650 597218
rect -8726 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 592650 597134
rect -8726 596866 592650 596898
rect -8726 592954 592650 592986
rect -8726 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 592650 592954
rect -8726 592634 592650 592718
rect -8726 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 592650 592634
rect -8726 592366 592650 592398
rect -8726 588454 592650 588486
rect -8726 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 592650 588454
rect -8726 588134 592650 588218
rect -8726 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 592650 588134
rect -8726 587866 592650 587898
rect -8726 583954 592650 583986
rect -8726 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 592650 583954
rect -8726 583634 592650 583718
rect -8726 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 592650 583634
rect -8726 583366 592650 583398
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 574954 592650 574986
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect -8726 574634 592650 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect -8726 574366 592650 574398
rect -8726 570454 592650 570486
rect -8726 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 592650 570454
rect -8726 570134 592650 570218
rect -8726 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 592650 570134
rect -8726 569866 592650 569898
rect -8726 565954 592650 565986
rect -8726 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 592650 565954
rect -8726 565634 592650 565718
rect -8726 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 592650 565634
rect -8726 565366 592650 565398
rect -8726 561454 592650 561486
rect -8726 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 592650 561454
rect -8726 561134 592650 561218
rect -8726 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 592650 561134
rect -8726 560866 592650 560898
rect -8726 556954 592650 556986
rect -8726 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 592650 556954
rect -8726 556634 592650 556718
rect -8726 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 592650 556634
rect -8726 556366 592650 556398
rect -8726 552454 592650 552486
rect -8726 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 592650 552454
rect -8726 552134 592650 552218
rect -8726 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 592650 552134
rect -8726 551866 592650 551898
rect -8726 547954 592650 547986
rect -8726 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 592650 547954
rect -8726 547634 592650 547718
rect -8726 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 592650 547634
rect -8726 547366 592650 547398
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 538954 592650 538986
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect -8726 538634 592650 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect -8726 538366 592650 538398
rect -8726 534454 592650 534486
rect -8726 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 592650 534454
rect -8726 534134 592650 534218
rect -8726 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 592650 534134
rect -8726 533866 592650 533898
rect -8726 529954 592650 529986
rect -8726 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 592650 529954
rect -8726 529634 592650 529718
rect -8726 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 592650 529634
rect -8726 529366 592650 529398
rect -8726 525454 592650 525486
rect -8726 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 592650 525454
rect -8726 525134 592650 525218
rect -8726 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 592650 525134
rect -8726 524866 592650 524898
rect -8726 520954 592650 520986
rect -8726 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 592650 520954
rect -8726 520634 592650 520718
rect -8726 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 592650 520634
rect -8726 520366 592650 520398
rect -8726 516454 592650 516486
rect -8726 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 592650 516454
rect -8726 516134 592650 516218
rect -8726 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 592650 516134
rect -8726 515866 592650 515898
rect -8726 511954 592650 511986
rect -8726 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 592650 511954
rect -8726 511634 592650 511718
rect -8726 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 592650 511634
rect -8726 511366 592650 511398
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 502954 592650 502986
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect -8726 502634 592650 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect -8726 502366 592650 502398
rect -8726 498454 592650 498486
rect -8726 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 592650 498454
rect -8726 498134 592650 498218
rect -8726 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 592650 498134
rect -8726 497866 592650 497898
rect -8726 493954 592650 493986
rect -8726 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 592650 493954
rect -8726 493634 592650 493718
rect -8726 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 592650 493634
rect -8726 493366 592650 493398
rect -8726 489454 592650 489486
rect -8726 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 592650 489454
rect -8726 489134 592650 489218
rect -8726 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 592650 489134
rect -8726 488866 592650 488898
rect -8726 484954 592650 484986
rect -8726 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 592650 484954
rect -8726 484634 592650 484718
rect -8726 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 592650 484634
rect -8726 484366 592650 484398
rect -8726 480454 592650 480486
rect -8726 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 592650 480454
rect -8726 480134 592650 480218
rect -8726 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 592650 480134
rect -8726 479866 592650 479898
rect -8726 475954 592650 475986
rect -8726 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 592650 475954
rect -8726 475634 592650 475718
rect -8726 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 592650 475634
rect -8726 475366 592650 475398
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 466954 592650 466986
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect -8726 466634 592650 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect -8726 466366 592650 466398
rect -8726 462454 592650 462486
rect -8726 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 592650 462454
rect -8726 462134 592650 462218
rect -8726 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 592650 462134
rect -8726 461866 592650 461898
rect -8726 457954 592650 457986
rect -8726 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 592650 457954
rect -8726 457634 592650 457718
rect -8726 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 592650 457634
rect -8726 457366 592650 457398
rect -8726 453454 592650 453486
rect -8726 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 592650 453454
rect -8726 453134 592650 453218
rect -8726 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 592650 453134
rect -8726 452866 592650 452898
rect -8726 448954 592650 448986
rect -8726 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 592650 448954
rect -8726 448634 592650 448718
rect -8726 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 592650 448634
rect -8726 448366 592650 448398
rect -8726 444454 592650 444486
rect -8726 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 592650 444454
rect -8726 444134 592650 444218
rect -8726 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 592650 444134
rect -8726 443866 592650 443898
rect -8726 439954 592650 439986
rect -8726 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 592650 439954
rect -8726 439634 592650 439718
rect -8726 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 592650 439634
rect -8726 439366 592650 439398
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 430954 592650 430986
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect -8726 430634 592650 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect -8726 430366 592650 430398
rect -8726 426454 592650 426486
rect -8726 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 592650 426454
rect -8726 426134 592650 426218
rect -8726 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 592650 426134
rect -8726 425866 592650 425898
rect -8726 421954 592650 421986
rect -8726 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 592650 421954
rect -8726 421634 592650 421718
rect -8726 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 592650 421634
rect -8726 421366 592650 421398
rect -8726 417454 592650 417486
rect -8726 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 592650 417454
rect -8726 417134 592650 417218
rect -8726 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 592650 417134
rect -8726 416866 592650 416898
rect -8726 412954 592650 412986
rect -8726 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 592650 412954
rect -8726 412634 592650 412718
rect -8726 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 592650 412634
rect -8726 412366 592650 412398
rect -8726 408454 592650 408486
rect -8726 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 592650 408454
rect -8726 408134 592650 408218
rect -8726 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 592650 408134
rect -8726 407866 592650 407898
rect -8726 403954 592650 403986
rect -8726 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 592650 403954
rect -8726 403634 592650 403718
rect -8726 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 592650 403634
rect -8726 403366 592650 403398
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 394954 592650 394986
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect -8726 394634 592650 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect -8726 394366 592650 394398
rect -8726 390454 592650 390486
rect -8726 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 592650 390454
rect -8726 390134 592650 390218
rect -8726 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 592650 390134
rect -8726 389866 592650 389898
rect -8726 385954 592650 385986
rect -8726 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 592650 385954
rect -8726 385634 592650 385718
rect -8726 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 592650 385634
rect -8726 385366 592650 385398
rect -8726 381454 592650 381486
rect -8726 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 592650 381454
rect -8726 381134 592650 381218
rect -8726 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 592650 381134
rect -8726 380866 592650 380898
rect -8726 376954 592650 376986
rect -8726 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 592650 376954
rect -8726 376634 592650 376718
rect -8726 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 592650 376634
rect -8726 376366 592650 376398
rect -8726 372454 592650 372486
rect -8726 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 592650 372454
rect -8726 372134 592650 372218
rect -8726 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 592650 372134
rect -8726 371866 592650 371898
rect -8726 367954 592650 367986
rect -8726 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 592650 367954
rect -8726 367634 592650 367718
rect -8726 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 592650 367634
rect -8726 367366 592650 367398
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 358954 592650 358986
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect -8726 358634 592650 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect -8726 358366 592650 358398
rect -8726 354454 592650 354486
rect -8726 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 244826 354454
rect 245062 354218 245146 354454
rect 245382 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 592650 354454
rect -8726 354134 592650 354218
rect -8726 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 244826 354134
rect 245062 353898 245146 354134
rect 245382 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 592650 354134
rect -8726 353866 592650 353898
rect -8726 349954 592650 349986
rect -8726 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 240326 349954
rect 240562 349718 240646 349954
rect 240882 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 592650 349954
rect -8726 349634 592650 349718
rect -8726 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 240326 349634
rect 240562 349398 240646 349634
rect 240882 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 592650 349634
rect -8726 349366 592650 349398
rect -8726 345454 592650 345486
rect -8726 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 592650 345454
rect -8726 345134 592650 345218
rect -8726 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 592650 345134
rect -8726 344866 592650 344898
rect -8726 340954 592650 340986
rect -8726 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 592650 340954
rect -8726 340634 592650 340718
rect -8726 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 592650 340634
rect -8726 340366 592650 340398
rect -8726 336454 592650 336486
rect -8726 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 592650 336454
rect -8726 336134 592650 336218
rect -8726 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 592650 336134
rect -8726 335866 592650 335898
rect -8726 331954 592650 331986
rect -8726 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 592650 331954
rect -8726 331634 592650 331718
rect -8726 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 592650 331634
rect -8726 331366 592650 331398
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 322954 592650 322986
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect -8726 322634 592650 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect -8726 322366 592650 322398
rect -8726 318454 592650 318486
rect -8726 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 592650 318454
rect -8726 318134 592650 318218
rect -8726 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 592650 318134
rect -8726 317866 592650 317898
rect -8726 313954 592650 313986
rect -8726 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 592650 313954
rect -8726 313634 592650 313718
rect -8726 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 592650 313634
rect -8726 313366 592650 313398
rect -8726 309454 592650 309486
rect -8726 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 592650 309454
rect -8726 309134 592650 309218
rect -8726 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 592650 309134
rect -8726 308866 592650 308898
rect -8726 304954 592650 304986
rect -8726 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 592650 304954
rect -8726 304634 592650 304718
rect -8726 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 592650 304634
rect -8726 304366 592650 304398
rect -8726 300454 592650 300486
rect -8726 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 592650 300454
rect -8726 300134 592650 300218
rect -8726 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 592650 300134
rect -8726 299866 592650 299898
rect -8726 295954 592650 295986
rect -8726 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 592650 295954
rect -8726 295634 592650 295718
rect -8726 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 592650 295634
rect -8726 295366 592650 295398
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 286954 592650 286986
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect -8726 286634 592650 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect -8726 286366 592650 286398
rect -8726 282454 592650 282486
rect -8726 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 592650 282454
rect -8726 282134 592650 282218
rect -8726 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 592650 282134
rect -8726 281866 592650 281898
rect -8726 277954 592650 277986
rect -8726 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 592650 277954
rect -8726 277634 592650 277718
rect -8726 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 592650 277634
rect -8726 277366 592650 277398
rect -8726 273454 592650 273486
rect -8726 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 592650 273454
rect -8726 273134 592650 273218
rect -8726 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 592650 273134
rect -8726 272866 592650 272898
rect -8726 268954 592650 268986
rect -8726 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 592650 268954
rect -8726 268634 592650 268718
rect -8726 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 592650 268634
rect -8726 268366 592650 268398
rect -8726 264454 592650 264486
rect -8726 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 592650 264454
rect -8726 264134 592650 264218
rect -8726 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 592650 264134
rect -8726 263866 592650 263898
rect -8726 259954 592650 259986
rect -8726 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 592650 259954
rect -8726 259634 592650 259718
rect -8726 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 592650 259634
rect -8726 259366 592650 259398
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 250954 592650 250986
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect -8726 250634 592650 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect -8726 250366 592650 250398
rect -8726 246454 592650 246486
rect -8726 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 136826 246454
rect 137062 246218 137146 246454
rect 137382 246218 172826 246454
rect 173062 246218 173146 246454
rect 173382 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 592650 246454
rect -8726 246134 592650 246218
rect -8726 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 136826 246134
rect 137062 245898 137146 246134
rect 137382 245898 172826 246134
rect 173062 245898 173146 246134
rect 173382 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 592650 246134
rect -8726 245866 592650 245898
rect -8726 241954 592650 241986
rect -8726 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 132326 241954
rect 132562 241718 132646 241954
rect 132882 241718 168326 241954
rect 168562 241718 168646 241954
rect 168882 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 240326 241954
rect 240562 241718 240646 241954
rect 240882 241718 276326 241954
rect 276562 241718 276646 241954
rect 276882 241718 312326 241954
rect 312562 241718 312646 241954
rect 312882 241718 348326 241954
rect 348562 241718 348646 241954
rect 348882 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 592650 241954
rect -8726 241634 592650 241718
rect -8726 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 132326 241634
rect 132562 241398 132646 241634
rect 132882 241398 168326 241634
rect 168562 241398 168646 241634
rect 168882 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 240326 241634
rect 240562 241398 240646 241634
rect 240882 241398 276326 241634
rect 276562 241398 276646 241634
rect 276882 241398 312326 241634
rect 312562 241398 312646 241634
rect 312882 241398 348326 241634
rect 348562 241398 348646 241634
rect 348882 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 592650 241634
rect -8726 241366 592650 241398
rect -8726 237454 592650 237486
rect -8726 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 592650 237454
rect -8726 237134 592650 237218
rect -8726 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 592650 237134
rect -8726 236866 592650 236898
rect -8726 232954 592650 232986
rect -8726 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 123326 232954
rect 123562 232718 123646 232954
rect 123882 232718 159326 232954
rect 159562 232718 159646 232954
rect 159882 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 231326 232954
rect 231562 232718 231646 232954
rect 231882 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 303326 232954
rect 303562 232718 303646 232954
rect 303882 232718 339326 232954
rect 339562 232718 339646 232954
rect 339882 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 592650 232954
rect -8726 232634 592650 232718
rect -8726 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 123326 232634
rect 123562 232398 123646 232634
rect 123882 232398 159326 232634
rect 159562 232398 159646 232634
rect 159882 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 231326 232634
rect 231562 232398 231646 232634
rect 231882 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 303326 232634
rect 303562 232398 303646 232634
rect 303882 232398 339326 232634
rect 339562 232398 339646 232634
rect 339882 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 592650 232634
rect -8726 232366 592650 232398
rect -8726 228454 592650 228486
rect -8726 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 118826 228454
rect 119062 228218 119146 228454
rect 119382 228218 154826 228454
rect 155062 228218 155146 228454
rect 155382 228218 190826 228454
rect 191062 228218 191146 228454
rect 191382 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 298826 228454
rect 299062 228218 299146 228454
rect 299382 228218 334826 228454
rect 335062 228218 335146 228454
rect 335382 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 592650 228454
rect -8726 228134 592650 228218
rect -8726 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 118826 228134
rect 119062 227898 119146 228134
rect 119382 227898 154826 228134
rect 155062 227898 155146 228134
rect 155382 227898 190826 228134
rect 191062 227898 191146 228134
rect 191382 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 298826 228134
rect 299062 227898 299146 228134
rect 299382 227898 334826 228134
rect 335062 227898 335146 228134
rect 335382 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 592650 228134
rect -8726 227866 592650 227898
rect -8726 223954 592650 223986
rect -8726 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 150326 223954
rect 150562 223718 150646 223954
rect 150882 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 592650 223954
rect -8726 223634 592650 223718
rect -8726 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 150326 223634
rect 150562 223398 150646 223634
rect 150882 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 592650 223634
rect -8726 223366 592650 223398
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 214954 592650 214986
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 141326 214954
rect 141562 214718 141646 214954
rect 141882 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect -8726 214634 592650 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 141326 214634
rect 141562 214398 141646 214634
rect 141882 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect -8726 214366 592650 214398
rect -8726 210454 592650 210486
rect -8726 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 136826 210454
rect 137062 210218 137146 210454
rect 137382 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 592650 210454
rect -8726 210134 592650 210218
rect -8726 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 136826 210134
rect 137062 209898 137146 210134
rect 137382 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 592650 210134
rect -8726 209866 592650 209898
rect -8726 205954 592650 205986
rect -8726 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205718 168326 205954
rect 168562 205718 168646 205954
rect 168882 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 592650 205954
rect -8726 205634 592650 205718
rect -8726 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205398 168326 205634
rect 168562 205398 168646 205634
rect 168882 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 592650 205634
rect -8726 205366 592650 205398
rect -8726 201454 592650 201486
rect -8726 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 592650 201454
rect -8726 201134 592650 201218
rect -8726 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 592650 201134
rect -8726 200866 592650 200898
rect -8726 196954 592650 196986
rect -8726 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 592650 196954
rect -8726 196634 592650 196718
rect -8726 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 592650 196634
rect -8726 196366 592650 196398
rect -8726 192454 592650 192486
rect -8726 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 592650 192454
rect -8726 192134 592650 192218
rect -8726 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 592650 192134
rect -8726 191866 592650 191898
rect -8726 187954 592650 187986
rect -8726 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 592650 187954
rect -8726 187634 592650 187718
rect -8726 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 592650 187634
rect -8726 187366 592650 187398
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 178954 592650 178986
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect -8726 178634 592650 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect -8726 178366 592650 178398
rect -8726 174454 592650 174486
rect -8726 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 136826 174454
rect 137062 174218 137146 174454
rect 137382 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 316826 174454
rect 317062 174218 317146 174454
rect 317382 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 592650 174454
rect -8726 174134 592650 174218
rect -8726 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 136826 174134
rect 137062 173898 137146 174134
rect 137382 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 316826 174134
rect 317062 173898 317146 174134
rect 317382 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 592650 174134
rect -8726 173866 592650 173898
rect -8726 169954 592650 169986
rect -8726 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 132326 169954
rect 132562 169718 132646 169954
rect 132882 169718 168326 169954
rect 168562 169718 168646 169954
rect 168882 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 312326 169954
rect 312562 169718 312646 169954
rect 312882 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 592650 169954
rect -8726 169634 592650 169718
rect -8726 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 132326 169634
rect 132562 169398 132646 169634
rect 132882 169398 168326 169634
rect 168562 169398 168646 169634
rect 168882 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 312326 169634
rect 312562 169398 312646 169634
rect 312882 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 592650 169634
rect -8726 169366 592650 169398
rect -8726 165454 592650 165486
rect -8726 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 592650 165454
rect -8726 165134 592650 165218
rect -8726 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 592650 165134
rect -8726 164866 592650 164898
rect -8726 160954 592650 160986
rect -8726 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 159326 160954
rect 159562 160718 159646 160954
rect 159882 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 592650 160954
rect -8726 160634 592650 160718
rect -8726 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 159326 160634
rect 159562 160398 159646 160634
rect 159882 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 592650 160634
rect -8726 160366 592650 160398
rect -8726 156454 592650 156486
rect -8726 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 592650 156454
rect -8726 156134 592650 156218
rect -8726 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 592650 156134
rect -8726 155866 592650 155898
rect -8726 151954 592650 151986
rect -8726 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 150326 151954
rect 150562 151718 150646 151954
rect 150882 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 592650 151954
rect -8726 151634 592650 151718
rect -8726 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 150326 151634
rect 150562 151398 150646 151634
rect 150882 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 592650 151634
rect -8726 151366 592650 151398
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 142954 592650 142986
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 141326 142954
rect 141562 142718 141646 142954
rect 141882 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect -8726 142634 592650 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 141326 142634
rect 141562 142398 141646 142634
rect 141882 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect -8726 142366 592650 142398
rect -8726 138454 592650 138486
rect -8726 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 592650 138454
rect -8726 138134 592650 138218
rect -8726 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 592650 138134
rect -8726 137866 592650 137898
rect -8726 133954 592650 133986
rect -8726 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 592650 133954
rect -8726 133634 592650 133718
rect -8726 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 592650 133634
rect -8726 133366 592650 133398
rect -8726 129454 592650 129486
rect -8726 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 592650 129454
rect -8726 129134 592650 129218
rect -8726 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 592650 129134
rect -8726 128866 592650 128898
rect -8726 124954 592650 124986
rect -8726 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 592650 124954
rect -8726 124634 592650 124718
rect -8726 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 592650 124634
rect -8726 124366 592650 124398
rect -8726 120454 592650 120486
rect -8726 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 592650 120454
rect -8726 120134 592650 120218
rect -8726 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 592650 120134
rect -8726 119866 592650 119898
rect -8726 115954 592650 115986
rect -8726 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 139610 115954
rect 139846 115718 170330 115954
rect 170566 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 592650 115954
rect -8726 115634 592650 115718
rect -8726 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 139610 115634
rect 139846 115398 170330 115634
rect 170566 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 592650 115634
rect -8726 115366 592650 115398
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 124250 111454
rect 124486 111218 154970 111454
rect 155206 111218 185690 111454
rect 185926 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 124250 111134
rect 124486 110898 154970 111134
rect 155206 110898 185690 111134
rect 185926 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 106954 592650 106986
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect -8726 106634 592650 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect -8726 106366 592650 106398
rect -8726 102454 592650 102486
rect -8726 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 592650 102454
rect -8726 102134 592650 102218
rect -8726 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 592650 102134
rect -8726 101866 592650 101898
rect -8726 97954 592650 97986
rect -8726 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 592650 97954
rect -8726 97634 592650 97718
rect -8726 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 592650 97634
rect -8726 97366 592650 97398
rect -8726 93454 592650 93486
rect -8726 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 592650 93454
rect -8726 93134 592650 93218
rect -8726 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 592650 93134
rect -8726 92866 592650 92898
rect -8726 88954 592650 88986
rect -8726 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 592650 88954
rect -8726 88634 592650 88718
rect -8726 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 592650 88634
rect -8726 88366 592650 88398
rect -8726 84454 592650 84486
rect -8726 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 592650 84454
rect -8726 84134 592650 84218
rect -8726 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 592650 84134
rect -8726 83866 592650 83898
rect -8726 79954 592650 79986
rect -8726 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 592650 79954
rect -8726 79634 592650 79718
rect -8726 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 592650 79634
rect -8726 79366 592650 79398
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 70954 592650 70986
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect -8726 70634 592650 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect -8726 70366 592650 70398
rect -8726 66454 592650 66486
rect -8726 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 592650 66454
rect -8726 66134 592650 66218
rect -8726 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 592650 66134
rect -8726 65866 592650 65898
rect -8726 61954 592650 61986
rect -8726 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 592650 61954
rect -8726 61634 592650 61718
rect -8726 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 592650 61634
rect -8726 61366 592650 61398
rect -8726 57454 592650 57486
rect -8726 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 592650 57454
rect -8726 57134 592650 57218
rect -8726 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 592650 57134
rect -8726 56866 592650 56898
rect -8726 52954 592650 52986
rect -8726 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 592650 52954
rect -8726 52634 592650 52718
rect -8726 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 592650 52634
rect -8726 52366 592650 52398
rect -8726 48454 592650 48486
rect -8726 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 592650 48454
rect -8726 48134 592650 48218
rect -8726 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 592650 48134
rect -8726 47866 592650 47898
rect -8726 43954 592650 43986
rect -8726 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 592650 43954
rect -8726 43634 592650 43718
rect -8726 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 592650 43634
rect -8726 43366 592650 43398
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 34954 592650 34986
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect -8726 34634 592650 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect -8726 34366 592650 34398
rect -8726 30454 592650 30486
rect -8726 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 592650 30454
rect -8726 30134 592650 30218
rect -8726 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 592650 30134
rect -8726 29866 592650 29898
rect -8726 25954 592650 25986
rect -8726 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 592650 25954
rect -8726 25634 592650 25718
rect -8726 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 592650 25634
rect -8726 25366 592650 25398
rect -8726 21454 592650 21486
rect -8726 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 592650 21454
rect -8726 21134 592650 21218
rect -8726 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 592650 21134
rect -8726 20866 592650 20898
rect -8726 16954 592650 16986
rect -8726 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 592650 16954
rect -8726 16634 592650 16718
rect -8726 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 592650 16634
rect -8726 16366 592650 16398
rect -8726 12454 592650 12486
rect -8726 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 592650 12454
rect -8726 12134 592650 12218
rect -8726 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 592650 12134
rect -8726 11866 592650 11898
rect -8726 7954 592650 7986
rect -8726 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 592650 7954
rect -8726 7634 592650 7718
rect -8726 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 592650 7634
rect -8726 7366 592650 7398
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use rlbp_macro  rlbp_macro0
timestamp 0
transform 1 0 120000 0 1 80000
box 0 0 70000 60000
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 78000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 142000 146414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 78000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 142000 182414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 10794 -7654 11414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 46794 -7654 47414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 -7654 83414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 -7654 119414 78000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 142000 119414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 -7654 155414 78000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 142000 155414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 -7654 191414 78000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 142000 191414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 -7654 227414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 -7654 263414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 -7654 299414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 -7654 335414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 -7654 371414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 406794 -7654 407414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 442794 -7654 443414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 478794 -7654 479414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 514794 -7654 515414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 550794 -7654 551414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 11866 592650 12486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 47866 592650 48486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 83866 592650 84486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 119866 592650 120486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 155866 592650 156486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 191866 592650 192486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 227866 592650 228486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 263866 592650 264486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 299866 592650 300486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 335866 592650 336486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 371866 592650 372486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 407866 592650 408486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 443866 592650 444486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 479866 592650 480486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 515866 592650 516486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 551866 592650 552486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 587866 592650 588486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 623866 592650 624486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 659866 592650 660486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 695866 592650 696486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 19794 -7654 20414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 55794 -7654 56414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 -7654 92414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 -7654 128414 78000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 142000 128414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 -7654 164414 78000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 142000 164414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 -7654 200414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 -7654 236414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 271794 -7654 272414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 -7654 308414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 343794 -7654 344414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 -7654 380414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 415794 -7654 416414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 451794 -7654 452414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 487794 -7654 488414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 523794 -7654 524414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 559794 -7654 560414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 20866 592650 21486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 56866 592650 57486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 92866 592650 93486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 128866 592650 129486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 164866 592650 165486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 200866 592650 201486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 236866 592650 237486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 272866 592650 273486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 308866 592650 309486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 344866 592650 345486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 380866 592650 381486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 416866 592650 417486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 452866 592650 453486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 488866 592650 489486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 524866 592650 525486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 560866 592650 561486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 596866 592650 597486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 632866 592650 633486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 668866 592650 669486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 28794 -7654 29414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 64794 -7654 65414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 100794 -7654 101414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 -7654 137414 78000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 142000 137414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 -7654 173414 78000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 142000 173414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 208794 -7654 209414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 244794 -7654 245414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 280794 -7654 281414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 316794 -7654 317414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 352794 -7654 353414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 388794 -7654 389414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 424794 -7654 425414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 460794 -7654 461414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 496794 -7654 497414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 532794 -7654 533414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 568794 -7654 569414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 29866 592650 30486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 65866 592650 66486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 101866 592650 102486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 137866 592650 138486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 173866 592650 174486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 209866 592650 210486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 245866 592650 246486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 281866 592650 282486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 317866 592650 318486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 353866 592650 354486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 389866 592650 390486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 425866 592650 426486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 461866 592650 462486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 497866 592650 498486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 533866 592650 534486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 569866 592650 570486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 605866 592650 606486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 641866 592650 642486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 677866 592650 678486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 24294 -7654 24914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 60294 -7654 60914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 96294 -7654 96914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 -7654 132914 78000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 142000 132914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 -7654 168914 78000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 142000 168914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 204294 -7654 204914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 240294 -7654 240914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 276294 -7654 276914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 -7654 312914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 348294 -7654 348914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 384294 -7654 384914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 420294 -7654 420914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 456294 -7654 456914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 492294 -7654 492914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 528294 -7654 528914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 564294 -7654 564914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 25366 592650 25986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 61366 592650 61986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 97366 592650 97986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 133366 592650 133986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 169366 592650 169986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 205366 592650 205986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 241366 592650 241986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 277366 592650 277986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 313366 592650 313986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 349366 592650 349986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 385366 592650 385986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 421366 592650 421986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 457366 592650 457986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 493366 592650 493986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 529366 592650 529986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 565366 592650 565986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 601366 592650 601986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 637366 592650 637986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 673366 592650 673986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 33294 -7654 33914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 69294 -7654 69914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 -7654 105914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 -7654 141914 78000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 142000 141914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 -7654 177914 78000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 142000 177914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 213294 -7654 213914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 -7654 249914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 285294 -7654 285914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 321294 -7654 321914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 357294 -7654 357914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 393294 -7654 393914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 429294 -7654 429914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 465294 -7654 465914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 501294 -7654 501914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 537294 -7654 537914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 573294 -7654 573914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 34366 592650 34986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 70366 592650 70986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 106366 592650 106986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 142366 592650 142986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 178366 592650 178986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 214366 592650 214986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 250366 592650 250986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 286366 592650 286986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 322366 592650 322986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 358366 592650 358986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 394366 592650 394986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 430366 592650 430986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 466366 592650 466986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 502366 592650 502986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 538366 592650 538986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 574366 592650 574986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 610366 592650 610986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 646366 592650 646986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 682366 592650 682986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 6294 -7654 6914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 42294 -7654 42914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 -7654 78914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 -7654 114914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 -7654 150914 78000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 142000 150914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 -7654 186914 78000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 142000 186914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 -7654 222914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 -7654 258914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 -7654 294914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 -7654 330914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 -7654 366914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 402294 -7654 402914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 438294 -7654 438914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 474294 -7654 474914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 510294 -7654 510914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 546294 -7654 546914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 582294 -7654 582914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 7366 592650 7986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 43366 592650 43986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 79366 592650 79986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 115366 592650 115986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 151366 592650 151986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 187366 592650 187986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 223366 592650 223986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 259366 592650 259986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 295366 592650 295986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 331366 592650 331986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 367366 592650 367986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 403366 592650 403986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 439366 592650 439986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 475366 592650 475986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 511366 592650 511986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 547366 592650 547986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 583366 592650 583986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 619366 592650 619986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 655366 592650 655986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 691366 592650 691986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 15294 -7654 15914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 51294 -7654 51914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 -7654 87914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 -7654 123914 78000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 142000 123914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 -7654 159914 78000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 142000 159914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 -7654 195914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 -7654 231914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 -7654 267914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 -7654 303914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 -7654 339914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 -7654 375914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 411294 -7654 411914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 447294 -7654 447914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 483294 -7654 483914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 519294 -7654 519914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 555294 -7654 555914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 16366 592650 16986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 52366 592650 52986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 88366 592650 88986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 124366 592650 124986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 160366 592650 160986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 196366 592650 196986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 232366 592650 232986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 268366 592650 268986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 304366 592650 304986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 340366 592650 340986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 376366 592650 376986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 412366 592650 412986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 448366 592650 448986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 484366 592650 484986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 520366 592650 520986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 556366 592650 556986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 592366 592650 592986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 628366 592650 628986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 664366 592650 664986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 700366 592650 700986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
