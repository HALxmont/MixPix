VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO res
  CLASS BLOCK ;
  FOREIGN res ;
  ORIGIN 17.500 14.000 ;
  SIZE 58.500 BY 34.500 ;
  PIN in1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT -2.000 -14.000 5.500 -2.000 ;
    END
  END in1
  PIN in2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.000 -14.000 18.500 -2.000 ;
    END
  END in2
  PIN out1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.000 8.500 11.500 20.500 ;
    END
  END out1
  PIN out2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.500 8.500 25.000 20.500 ;
    END
  END out2
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT -17.500 1.000 -5.500 8.500 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 29.000 -2.000 41.000 5.500 ;
    END
  END VSS
  OBS
      LAYER li1 ;
        RECT -1.820 -0.320 24.830 6.300 ;
      LAYER met1 ;
        RECT -2.780 0.360 26.000 5.620 ;
      LAYER met2 ;
        RECT -5.220 8.220 3.720 8.500 ;
        RECT 11.780 8.220 17.220 8.500 ;
        RECT 25.280 8.220 29.000 8.500 ;
        RECT -5.220 5.780 29.000 8.220 ;
        RECT -5.220 0.720 28.720 5.780 ;
        RECT -5.500 -1.720 28.720 0.720 ;
        RECT -5.500 -2.000 -2.280 -1.720 ;
        RECT 5.780 -2.000 10.720 -1.720 ;
        RECT 18.780 -2.000 28.720 -1.720 ;
  END
END res
END LIBRARY

