magic
tech sky130B
magscale 1 2
timestamp 1668186310
<< metal1 >>
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 201494 702992 201500 703044
rect 201552 703032 201558 703044
rect 202782 703032 202788 703044
rect 201552 703004 202788 703032
rect 201552 702992 201558 703004
rect 202782 702992 202788 703004
rect 202840 702992 202846 703044
rect 331214 702992 331220 703044
rect 331272 703032 331278 703044
rect 332502 703032 332508 703044
rect 331272 703004 332508 703032
rect 331272 702992 331278 703004
rect 332502 702992 332508 703004
rect 332560 702992 332566 703044
rect 196618 700612 196624 700664
rect 196676 700652 196682 700664
rect 218974 700652 218980 700664
rect 196676 700624 218980 700652
rect 196676 700612 196682 700624
rect 218974 700612 218980 700624
rect 219032 700612 219038 700664
rect 193858 700544 193864 700596
rect 193916 700584 193922 700596
rect 283834 700584 283840 700596
rect 193916 700556 283840 700584
rect 193916 700544 193922 700556
rect 283834 700544 283840 700556
rect 283892 700544 283898 700596
rect 192478 700476 192484 700528
rect 192536 700516 192542 700528
rect 348786 700516 348792 700528
rect 192536 700488 348792 700516
rect 192536 700476 192542 700488
rect 348786 700476 348792 700488
rect 348844 700476 348850 700528
rect 189718 700408 189724 700460
rect 189776 700448 189782 700460
rect 413646 700448 413652 700460
rect 189776 700420 413652 700448
rect 189776 700408 189782 700420
rect 413646 700408 413652 700420
rect 413704 700408 413710 700460
rect 89162 700340 89168 700392
rect 89220 700380 89226 700392
rect 182542 700380 182548 700392
rect 89220 700352 182548 700380
rect 89220 700340 89226 700352
rect 182542 700340 182548 700352
rect 182600 700340 182606 700392
rect 188338 700340 188344 700392
rect 188396 700380 188402 700392
rect 478506 700380 478512 700392
rect 188396 700352 478512 700380
rect 188396 700340 188402 700352
rect 478506 700340 478512 700352
rect 478564 700340 478570 700392
rect 8110 700272 8116 700324
rect 8168 700312 8174 700324
rect 119338 700312 119344 700324
rect 8168 700284 119344 700312
rect 8168 700272 8174 700284
rect 119338 700272 119344 700284
rect 119396 700272 119402 700324
rect 137830 700272 137836 700324
rect 137888 700312 137894 700324
rect 180794 700312 180800 700324
rect 137888 700284 180800 700312
rect 137888 700272 137894 700284
rect 180794 700272 180800 700284
rect 180852 700272 180858 700324
rect 185578 700272 185584 700324
rect 185636 700312 185642 700324
rect 543458 700312 543464 700324
rect 185636 700284 543464 700312
rect 185636 700272 185642 700284
rect 543458 700272 543464 700284
rect 543516 700272 543522 700324
rect 105446 699660 105452 699712
rect 105504 699700 105510 699712
rect 106918 699700 106924 699712
rect 105504 699672 106924 699700
rect 105504 699660 105510 699672
rect 106918 699660 106924 699672
rect 106976 699660 106982 699712
rect 266354 697552 266360 697604
rect 266412 697592 266418 697604
rect 267642 697592 267648 697604
rect 266412 697564 267648 697592
rect 266412 697552 266418 697564
rect 267642 697552 267648 697564
rect 267700 697552 267706 697604
rect 2774 683680 2780 683732
rect 2832 683720 2838 683732
rect 4798 683720 4804 683732
rect 2832 683692 4804 683720
rect 2832 683680 2838 683692
rect 4798 683680 4804 683692
rect 4856 683680 4862 683732
rect 184198 683136 184204 683188
rect 184256 683176 184262 683188
rect 579614 683176 579620 683188
rect 184256 683148 579620 683176
rect 184256 683136 184262 683148
rect 579614 683136 579620 683148
rect 579672 683136 579678 683188
rect 3326 632068 3332 632120
rect 3384 632108 3390 632120
rect 7558 632108 7564 632120
rect 3384 632080 7564 632108
rect 3384 632068 3390 632080
rect 7558 632068 7564 632080
rect 7616 632068 7622 632120
rect 184290 630640 184296 630692
rect 184348 630680 184354 630692
rect 580166 630680 580172 630692
rect 184348 630652 580172 630680
rect 184348 630640 184354 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 120718 616836 120724 616888
rect 120776 616876 120782 616888
rect 579982 616876 579988 616888
rect 120776 616848 579988 616876
rect 120776 616836 120782 616848
rect 579982 616836 579988 616848
rect 580040 616836 580046 616888
rect 3142 579640 3148 579692
rect 3200 579680 3206 579692
rect 17218 579680 17224 579692
rect 3200 579652 17224 579680
rect 3200 579640 3206 579652
rect 17218 579640 17224 579652
rect 17276 579640 17282 579692
rect 184382 576852 184388 576904
rect 184440 576892 184446 576904
rect 579982 576892 579988 576904
rect 184440 576864 579988 576892
rect 184440 576852 184446 576864
rect 579982 576852 579988 576864
rect 580040 576852 580046 576904
rect 120810 563048 120816 563100
rect 120868 563088 120874 563100
rect 580166 563088 580172 563100
rect 120868 563060 580172 563088
rect 120868 563048 120874 563060
rect 580166 563048 580172 563060
rect 580224 563048 580230 563100
rect 3142 553392 3148 553444
rect 3200 553432 3206 553444
rect 115198 553432 115204 553444
rect 3200 553404 115204 553432
rect 3200 553392 3206 553404
rect 115198 553392 115204 553404
rect 115256 553392 115262 553444
rect 182358 536800 182364 536852
rect 182416 536840 182422 536852
rect 579614 536840 579620 536852
rect 182416 536812 579620 536840
rect 182416 536800 182422 536812
rect 579614 536800 579620 536812
rect 579672 536800 579678 536852
rect 3326 527824 3332 527876
rect 3384 527864 3390 527876
rect 8938 527864 8944 527876
rect 3384 527836 8944 527864
rect 3384 527824 3390 527836
rect 8938 527824 8944 527836
rect 8996 527824 9002 527876
rect 214558 524424 214564 524476
rect 214616 524464 214622 524476
rect 580166 524464 580172 524476
rect 214616 524436 580172 524464
rect 214616 524424 214622 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 3326 514768 3332 514820
rect 3384 514808 3390 514820
rect 180886 514808 180892 514820
rect 3384 514780 180892 514808
rect 3384 514768 3390 514780
rect 180886 514768 180892 514780
rect 180944 514768 180950 514820
rect 120902 510620 120908 510672
rect 120960 510660 120966 510672
rect 579614 510660 579620 510672
rect 120960 510632 579620 510660
rect 120960 510620 120966 510632
rect 579614 510620 579620 510632
rect 579672 510620 579678 510672
rect 2774 501032 2780 501084
rect 2832 501072 2838 501084
rect 4890 501072 4896 501084
rect 2832 501044 4896 501072
rect 2832 501032 2838 501044
rect 4890 501032 4896 501044
rect 4948 501032 4954 501084
rect 182266 484372 182272 484424
rect 182324 484412 182330 484424
rect 580166 484412 580172 484424
rect 182324 484384 580172 484412
rect 182324 484372 182330 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 211798 470568 211804 470620
rect 211856 470608 211862 470620
rect 579982 470608 579988 470620
rect 211856 470580 579988 470608
rect 211856 470568 211862 470580
rect 579982 470568 579988 470580
rect 580040 470568 580046 470620
rect 3050 462340 3056 462392
rect 3108 462380 3114 462392
rect 179414 462380 179420 462392
rect 3108 462352 179420 462380
rect 3108 462340 3114 462352
rect 179414 462340 179420 462352
rect 179472 462340 179478 462392
rect 3878 461592 3884 461644
rect 3936 461632 3942 461644
rect 53098 461632 53104 461644
rect 3936 461604 53104 461632
rect 3936 461592 3942 461604
rect 53098 461592 53104 461604
rect 53156 461592 53162 461644
rect 120994 456764 121000 456816
rect 121052 456804 121058 456816
rect 580166 456804 580172 456816
rect 121052 456776 580172 456804
rect 121052 456764 121058 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 2958 448536 2964 448588
rect 3016 448576 3022 448588
rect 44818 448576 44824 448588
rect 3016 448548 44824 448576
rect 3016 448536 3022 448548
rect 44818 448536 44824 448548
rect 44876 448536 44882 448588
rect 118694 429836 118700 429888
rect 118752 429876 118758 429888
rect 580626 429876 580632 429888
rect 118752 429848 580632 429876
rect 118752 429836 118758 429848
rect 580626 429836 580632 429848
rect 580684 429836 580690 429888
rect 3326 422288 3332 422340
rect 3384 422328 3390 422340
rect 10318 422328 10324 422340
rect 3384 422300 10324 422328
rect 3384 422288 3390 422300
rect 10318 422288 10324 422300
rect 10376 422288 10382 422340
rect 182818 418140 182824 418192
rect 182876 418180 182882 418192
rect 579706 418180 579712 418192
rect 182876 418152 579712 418180
rect 182876 418140 182882 418152
rect 579706 418140 579712 418152
rect 579764 418140 579770 418192
rect 118602 404336 118608 404388
rect 118660 404376 118666 404388
rect 580166 404376 580172 404388
rect 118660 404348 580172 404376
rect 118660 404336 118666 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 3326 397468 3332 397520
rect 3384 397508 3390 397520
rect 86218 397508 86224 397520
rect 3384 397480 86224 397508
rect 3384 397468 3390 397480
rect 86218 397468 86224 397480
rect 86276 397468 86282 397520
rect 3326 371220 3332 371272
rect 3384 371260 3390 371272
rect 84838 371260 84844 371272
rect 3384 371232 84844 371260
rect 3384 371220 3390 371232
rect 84838 371220 84844 371232
rect 84896 371220 84902 371272
rect 224218 364352 224224 364404
rect 224276 364392 224282 364404
rect 580166 364392 580172 364404
rect 224276 364364 580172 364392
rect 224276 364352 224282 364364
rect 580166 364352 580172 364364
rect 580224 364352 580230 364404
rect 3326 357416 3332 357468
rect 3384 357456 3390 357468
rect 180978 357456 180984 357468
rect 3384 357428 180984 357456
rect 3384 357416 3390 357428
rect 180978 357416 180984 357428
rect 181036 357416 181042 357468
rect 118510 351908 118516 351960
rect 118568 351948 118574 351960
rect 580166 351948 580172 351960
rect 118568 351920 580172 351948
rect 118568 351908 118574 351920
rect 580166 351908 580172 351920
rect 580224 351908 580230 351960
rect 3326 345040 3332 345092
rect 3384 345080 3390 345092
rect 116578 345080 116584 345092
rect 3384 345052 116584 345080
rect 3384 345040 3390 345052
rect 116578 345040 116584 345052
rect 116636 345040 116642 345092
rect 3142 318792 3148 318844
rect 3200 318832 3206 318844
rect 13078 318832 13084 318844
rect 3200 318804 13084 318832
rect 3200 318792 3206 318804
rect 13078 318792 13084 318804
rect 13136 318792 13142 318844
rect 221458 311856 221464 311908
rect 221516 311896 221522 311908
rect 580166 311896 580172 311908
rect 221516 311868 580172 311896
rect 221516 311856 221522 311868
rect 580166 311856 580172 311868
rect 580224 311856 580230 311908
rect 3326 304988 3332 305040
rect 3384 305028 3390 305040
rect 178678 305028 178684 305040
rect 3384 305000 178684 305028
rect 3384 304988 3390 305000
rect 178678 304988 178684 305000
rect 178736 304988 178742 305040
rect 124858 298120 124864 298172
rect 124916 298160 124922 298172
rect 580166 298160 580172 298172
rect 124916 298132 580172 298160
rect 124916 298120 124922 298132
rect 580166 298120 580172 298132
rect 580224 298120 580230 298172
rect 3326 292544 3332 292596
rect 3384 292584 3390 292596
rect 121086 292584 121092 292596
rect 3384 292556 121092 292584
rect 3384 292544 3390 292556
rect 121086 292544 121092 292556
rect 121144 292544 121150 292596
rect 180058 271872 180064 271924
rect 180116 271912 180122 271924
rect 579614 271912 579620 271924
rect 180116 271884 579620 271912
rect 180116 271872 180122 271884
rect 579614 271872 579620 271884
rect 579672 271872 579678 271924
rect 3234 266364 3240 266416
rect 3292 266404 3298 266416
rect 18598 266404 18604 266416
rect 3292 266376 18604 266404
rect 3292 266364 3298 266376
rect 18598 266364 18604 266376
rect 18656 266364 18662 266416
rect 220078 258068 220084 258120
rect 220136 258108 220142 258120
rect 580166 258108 580172 258120
rect 220136 258080 580172 258108
rect 220136 258068 220142 258080
rect 580166 258068 580172 258080
rect 580224 258068 580230 258120
rect 2958 253920 2964 253972
rect 3016 253960 3022 253972
rect 178770 253960 178776 253972
rect 3016 253932 178776 253960
rect 3016 253920 3022 253932
rect 178770 253920 178776 253932
rect 178828 253920 178834 253972
rect 128998 244264 129004 244316
rect 129056 244304 129062 244316
rect 579614 244304 579620 244316
rect 129056 244276 579620 244304
rect 129056 244264 129062 244276
rect 579614 244264 579620 244276
rect 579672 244264 579678 244316
rect 182174 233792 182180 233844
rect 182232 233832 182238 233844
rect 182542 233832 182548 233844
rect 182232 233804 182548 233832
rect 182232 233792 182238 233804
rect 182542 233792 182548 233804
rect 182600 233792 182606 233844
rect 182818 231548 182824 231600
rect 182876 231548 182882 231600
rect 182836 230376 182864 231548
rect 182818 230324 182824 230376
rect 182876 230324 182882 230376
rect 207658 229780 207664 229832
rect 207716 229820 207722 229832
rect 212534 229820 212540 229832
rect 207716 229792 212540 229820
rect 207716 229780 207722 229792
rect 212534 229780 212540 229792
rect 212592 229780 212598 229832
rect 161382 229712 161388 229764
rect 161440 229752 161446 229764
rect 392486 229752 392492 229764
rect 161440 229724 392492 229752
rect 161440 229712 161446 229724
rect 392486 229712 392492 229724
rect 392544 229712 392550 229764
rect 180150 229100 180156 229152
rect 180208 229140 180214 229152
rect 182542 229140 182548 229152
rect 180208 229112 182548 229140
rect 180208 229100 180214 229112
rect 182542 229100 182548 229112
rect 182600 229100 182606 229152
rect 123662 228352 123668 228404
rect 123720 228392 123726 228404
rect 143534 228392 143540 228404
rect 123720 228364 143540 228392
rect 123720 228352 123726 228364
rect 143534 228352 143540 228364
rect 143592 228352 143598 228404
rect 166258 228352 166264 228404
rect 166316 228392 166322 228404
rect 272518 228392 272524 228404
rect 166316 228364 272524 228392
rect 166316 228352 166322 228364
rect 272518 228352 272524 228364
rect 272576 228352 272582 228404
rect 2866 227740 2872 227792
rect 2924 227780 2930 227792
rect 138658 227780 138664 227792
rect 2924 227752 138664 227780
rect 2924 227740 2930 227752
rect 138658 227740 138664 227752
rect 138716 227740 138722 227792
rect 182174 224204 182180 224256
rect 182232 224244 182238 224256
rect 182542 224244 182548 224256
rect 182232 224216 182548 224244
rect 182232 224204 182238 224216
rect 182542 224204 182548 224216
rect 182600 224204 182606 224256
rect 217318 218016 217324 218068
rect 217376 218056 217382 218068
rect 579982 218056 579988 218068
rect 217376 218028 579988 218056
rect 217376 218016 217382 218028
rect 579982 218016 579988 218028
rect 580040 218016 580046 218068
rect 3326 213936 3332 213988
rect 3384 213976 3390 213988
rect 31018 213976 31024 213988
rect 3384 213948 31024 213976
rect 3384 213936 3390 213948
rect 31018 213936 31024 213948
rect 31076 213936 31082 213988
rect 144914 208360 144920 208412
rect 144972 208400 144978 208412
rect 151814 208400 151820 208412
rect 144972 208372 151820 208400
rect 144972 208360 144978 208372
rect 151814 208360 151820 208372
rect 151872 208360 151878 208412
rect 126238 205640 126244 205692
rect 126296 205680 126302 205692
rect 580166 205680 580172 205692
rect 126296 205652 580172 205680
rect 126296 205640 126302 205652
rect 580166 205640 580172 205652
rect 580224 205640 580230 205692
rect 154114 204892 154120 204944
rect 154172 204932 154178 204944
rect 242894 204932 242900 204944
rect 154172 204904 242900 204932
rect 154172 204892 154178 204904
rect 242894 204892 242900 204904
rect 242952 204892 242958 204944
rect 146202 203532 146208 203584
rect 146260 203572 146266 203584
rect 207658 203572 207664 203584
rect 146260 203544 207664 203572
rect 146260 203532 146266 203544
rect 207658 203532 207664 203544
rect 207716 203532 207722 203584
rect 147398 202104 147404 202156
rect 147456 202144 147462 202156
rect 180150 202144 180156 202156
rect 147456 202116 180156 202144
rect 147456 202104 147462 202116
rect 180150 202104 180156 202116
rect 180208 202104 180214 202156
rect 3326 201492 3332 201544
rect 3384 201532 3390 201544
rect 179598 201532 179604 201544
rect 3384 201504 179604 201532
rect 3384 201492 3390 201504
rect 179598 201492 179604 201504
rect 179656 201492 179662 201544
rect 159174 199384 159180 199436
rect 159232 199424 159238 199436
rect 362954 199424 362960 199436
rect 159232 199396 362960 199424
rect 159232 199384 159238 199396
rect 362954 199384 362960 199396
rect 363012 199384 363018 199436
rect 154574 198024 154580 198076
rect 154632 198064 154638 198076
rect 166258 198064 166264 198076
rect 154632 198036 166264 198064
rect 154632 198024 154638 198036
rect 166258 198024 166264 198036
rect 166316 198024 166322 198076
rect 157334 197956 157340 198008
rect 157392 197996 157398 198008
rect 332594 197996 332600 198008
rect 157392 197968 332600 197996
rect 157392 197956 157398 197968
rect 332594 197956 332600 197968
rect 332652 197956 332658 198008
rect 138658 196732 138664 196784
rect 138716 196772 138722 196784
rect 164234 196772 164240 196784
rect 138716 196744 164240 196772
rect 138716 196732 138722 196744
rect 164234 196732 164240 196744
rect 164292 196732 164298 196784
rect 153838 196664 153844 196716
rect 153896 196704 153902 196716
rect 181070 196704 181076 196716
rect 153896 196676 181076 196704
rect 153896 196664 153902 196676
rect 181070 196664 181076 196676
rect 181128 196664 181134 196716
rect 157242 196596 157248 196648
rect 157300 196636 157306 196648
rect 302234 196636 302240 196648
rect 157300 196608 302240 196636
rect 157300 196596 157306 196608
rect 302234 196596 302240 196608
rect 302292 196596 302298 196648
rect 152458 196460 152464 196512
rect 152516 196500 152522 196512
rect 154574 196500 154580 196512
rect 152516 196472 154580 196500
rect 152516 196460 152522 196472
rect 154574 196460 154580 196472
rect 154632 196460 154638 196512
rect 62114 195916 62120 195968
rect 62172 195956 62178 195968
rect 138106 195956 138112 195968
rect 62172 195928 138112 195956
rect 62172 195916 62178 195928
rect 138106 195916 138112 195928
rect 138164 195916 138170 195968
rect 153470 195916 153476 195968
rect 153528 195956 153534 195968
rect 154114 195956 154120 195968
rect 153528 195928 154120 195956
rect 153528 195916 153534 195928
rect 154114 195916 154120 195928
rect 154172 195916 154178 195968
rect 92474 195848 92480 195900
rect 92532 195888 92538 195900
rect 139394 195888 139400 195900
rect 92532 195860 139400 195888
rect 92532 195848 92538 195860
rect 139394 195848 139400 195860
rect 139452 195848 139458 195900
rect 148778 195644 148784 195696
rect 148836 195684 148842 195696
rect 165522 195684 165528 195696
rect 148836 195656 165528 195684
rect 148836 195644 148842 195656
rect 165522 195644 165528 195656
rect 165580 195644 165586 195696
rect 151446 191088 151452 191140
rect 151504 191088 151510 191140
rect 3326 187688 3332 187740
rect 3384 187728 3390 187740
rect 121178 187728 121184 187740
rect 3384 187700 121184 187728
rect 3384 187688 3390 187700
rect 121178 187688 121184 187700
rect 121236 187688 121242 187740
rect 162118 180928 162124 180940
rect 161676 180900 162124 180928
rect 144454 180684 144460 180736
rect 144512 180724 144518 180736
rect 146110 180724 146116 180736
rect 144512 180696 146116 180724
rect 144512 180684 144518 180696
rect 146110 180684 146116 180696
rect 146168 180684 146174 180736
rect 161474 180548 161480 180600
rect 161532 180588 161538 180600
rect 161676 180588 161704 180900
rect 162118 180888 162124 180900
rect 162176 180888 162182 180940
rect 161532 180560 161704 180588
rect 161532 180548 161538 180560
rect 136818 180316 136824 180328
rect 122806 180288 136824 180316
rect 17862 180072 17868 180124
rect 17920 180112 17926 180124
rect 122806 180112 122834 180288
rect 136818 180276 136824 180288
rect 136876 180276 136882 180328
rect 17920 180084 122834 180112
rect 17920 180072 17926 180084
rect 136634 180072 136640 180124
rect 136692 180112 136698 180124
rect 141234 180112 141240 180124
rect 136692 180084 141240 180112
rect 136692 180072 136698 180084
rect 141234 180072 141240 180084
rect 141292 180072 141298 180124
rect 143534 179596 143540 179648
rect 143592 179596 143598 179648
rect 122834 178780 122840 178832
rect 122892 178820 122898 178832
rect 136634 178820 136640 178832
rect 122892 178792 136640 178820
rect 122892 178780 122898 178792
rect 136634 178780 136640 178792
rect 136692 178780 136698 178832
rect 121454 178644 121460 178696
rect 121512 178684 121518 178696
rect 137002 178684 137008 178696
rect 121512 178656 137008 178684
rect 121512 178644 121518 178656
rect 137002 178644 137008 178656
rect 137060 178644 137066 178696
rect 143552 178684 143580 179596
rect 144178 178684 144184 178696
rect 143552 178656 144184 178684
rect 144178 178644 144184 178656
rect 144236 178644 144242 178696
rect 215938 178032 215944 178084
rect 215996 178072 216002 178084
rect 580166 178072 580172 178084
rect 215996 178044 580172 178072
rect 215996 178032 216002 178044
rect 580166 178032 580172 178044
rect 580224 178032 580230 178084
rect 140774 177828 140780 177880
rect 140832 177868 140838 177880
rect 141602 177868 141608 177880
rect 140832 177840 141608 177868
rect 140832 177828 140838 177840
rect 141602 177828 141608 177840
rect 141660 177828 141666 177880
rect 124214 177284 124220 177336
rect 124272 177324 124278 177336
rect 137094 177324 137100 177336
rect 124272 177296 137100 177324
rect 124272 177284 124278 177296
rect 137094 177284 137100 177296
rect 137152 177284 137158 177336
rect 3326 176604 3332 176656
rect 3384 176644 3390 176656
rect 17862 176644 17868 176656
rect 3384 176616 17868 176644
rect 3384 176604 3390 176616
rect 17862 176604 17868 176616
rect 17920 176604 17926 176656
rect 161382 176196 161388 176248
rect 161440 176196 161446 176248
rect 125594 175992 125600 176044
rect 125652 176032 125658 176044
rect 137186 176032 137192 176044
rect 125652 176004 137192 176032
rect 125652 175992 125658 176004
rect 137186 175992 137192 176004
rect 137244 175992 137250 176044
rect 128354 175924 128360 175976
rect 128412 175964 128418 175976
rect 137278 175964 137284 175976
rect 128412 175936 137284 175964
rect 128412 175924 128418 175936
rect 137278 175924 137284 175936
rect 137336 175924 137342 175976
rect 159082 175584 159088 175636
rect 159140 175624 159146 175636
rect 161400 175624 161428 176196
rect 159140 175596 161428 175624
rect 159140 175584 159146 175596
rect 165430 174972 165436 175024
rect 165488 174972 165494 175024
rect 165522 174972 165528 175024
rect 165580 174972 165586 175024
rect 163148 174752 163176 174866
rect 165448 174752 165476 174972
rect 165540 174752 165568 174972
rect 163130 174700 163136 174752
rect 163188 174700 163194 174752
rect 165430 174700 165436 174752
rect 165488 174700 165494 174752
rect 165522 174700 165528 174752
rect 165580 174700 165586 174752
rect 133874 173884 133880 173936
rect 133932 173924 133938 173936
rect 135254 173924 135260 173936
rect 133932 173896 135260 173924
rect 133932 173884 133938 173896
rect 135254 173884 135260 173896
rect 135312 173884 135318 173936
rect 140774 173816 140780 173868
rect 140832 173856 140838 173868
rect 141602 173856 141608 173868
rect 140832 173828 141608 173856
rect 140832 173816 140838 173828
rect 141602 173816 141608 173828
rect 141660 173816 141666 173868
rect 131114 173272 131120 173324
rect 131172 173312 131178 173324
rect 137370 173312 137376 173324
rect 131172 173284 137376 173312
rect 131172 173272 131178 173284
rect 137370 173272 137376 173284
rect 137428 173272 137434 173324
rect 126974 173204 126980 173256
rect 127032 173244 127038 173256
rect 140774 173244 140780 173256
rect 127032 173216 140780 173244
rect 127032 173204 127038 173216
rect 140774 173204 140780 173216
rect 140832 173204 140838 173256
rect 3786 173136 3792 173188
rect 3844 173176 3850 173188
rect 179690 173176 179696 173188
rect 3844 173148 179696 173176
rect 3844 173136 3850 173148
rect 179690 173136 179696 173148
rect 179748 173136 179754 173188
rect 135254 172388 135260 172440
rect 135312 172428 135318 172440
rect 138934 172428 138940 172440
rect 135312 172400 138940 172428
rect 135312 172388 135318 172400
rect 138934 172388 138940 172400
rect 138992 172388 138998 172440
rect 132494 172184 132500 172236
rect 132552 172224 132558 172236
rect 137462 172224 137468 172236
rect 132552 172196 137468 172224
rect 132552 172184 132558 172196
rect 137462 172184 137468 172196
rect 137520 172184 137526 172236
rect 138014 171368 138020 171420
rect 138072 171408 138078 171420
rect 140958 171408 140964 171420
rect 138072 171380 140964 171408
rect 138072 171368 138078 171380
rect 140958 171368 140964 171380
rect 141016 171368 141022 171420
rect 122098 165588 122104 165640
rect 122156 165628 122162 165640
rect 579798 165628 579804 165640
rect 122156 165600 579804 165628
rect 122156 165588 122162 165600
rect 579798 165588 579804 165600
rect 579856 165588 579862 165640
rect 162854 164704 162860 164756
rect 162912 164744 162918 164756
rect 163590 164744 163596 164756
rect 162912 164716 163596 164744
rect 162912 164704 162918 164716
rect 163590 164704 163596 164716
rect 163648 164704 163654 164756
rect 165522 164160 165528 164212
rect 165580 164200 165586 164212
rect 168374 164200 168380 164212
rect 165580 164172 168380 164200
rect 165580 164160 165586 164172
rect 168374 164160 168380 164172
rect 168432 164160 168438 164212
rect 3326 162868 3332 162920
rect 3384 162908 3390 162920
rect 14458 162908 14464 162920
rect 3384 162880 14464 162908
rect 3384 162868 3390 162880
rect 14458 162868 14464 162880
rect 14516 162868 14522 162920
rect 165430 162800 165436 162852
rect 165488 162840 165494 162852
rect 169846 162840 169852 162852
rect 165488 162812 169852 162840
rect 165488 162800 165494 162812
rect 169846 162800 169852 162812
rect 169904 162800 169910 162852
rect 182910 151784 182916 151836
rect 182968 151824 182974 151836
rect 579982 151824 579988 151836
rect 182968 151796 579988 151824
rect 182968 151784 182974 151796
rect 579982 151784 579988 151796
rect 580040 151784 580046 151836
rect 3694 151036 3700 151088
rect 3752 151076 3758 151088
rect 181254 151076 181260 151088
rect 3752 151048 181260 151076
rect 3752 151036 3758 151048
rect 181254 151036 181260 151048
rect 181312 151036 181318 151088
rect 3510 150016 3516 150068
rect 3568 150056 3574 150068
rect 3694 150056 3700 150068
rect 3568 150028 3700 150056
rect 3568 150016 3574 150028
rect 3694 150016 3700 150028
rect 3752 150016 3758 150068
rect 3510 149064 3516 149116
rect 3568 149104 3574 149116
rect 181162 149104 181168 149116
rect 3568 149076 181168 149104
rect 3568 149064 3574 149076
rect 181162 149064 181168 149076
rect 181220 149064 181226 149116
rect 3694 148316 3700 148368
rect 3752 148356 3758 148368
rect 181346 148356 181352 148368
rect 3752 148328 181352 148356
rect 3752 148316 3758 148328
rect 181346 148316 181352 148328
rect 181404 148316 181410 148368
rect 119062 146956 119068 147008
rect 119120 146996 119126 147008
rect 234614 146996 234620 147008
rect 119120 146968 234620 146996
rect 119120 146956 119126 146968
rect 234614 146956 234620 146968
rect 234672 146956 234678 147008
rect 23474 146888 23480 146940
rect 23532 146928 23538 146940
rect 179782 146928 179788 146940
rect 23532 146900 179788 146928
rect 23532 146888 23538 146900
rect 179782 146888 179788 146900
rect 179840 146888 179846 146940
rect 119154 145528 119160 145580
rect 119212 145568 119218 145580
rect 299474 145568 299480 145580
rect 119212 145540 299480 145568
rect 119212 145528 119218 145540
rect 299474 145528 299480 145540
rect 299532 145528 299538 145580
rect 118878 144168 118884 144220
rect 118936 144208 118942 144220
rect 429194 144208 429200 144220
rect 118936 144180 429200 144208
rect 118936 144168 118942 144180
rect 429194 144168 429200 144180
rect 429252 144168 429258 144220
rect 151814 143488 151820 143540
rect 151872 143528 151878 143540
rect 157426 143528 157432 143540
rect 151872 143500 157432 143528
rect 151872 143488 151878 143500
rect 157426 143488 157432 143500
rect 157484 143488 157490 143540
rect 164050 143488 164056 143540
rect 164108 143528 164114 143540
rect 166166 143528 166172 143540
rect 164108 143500 166172 143528
rect 164108 143488 164114 143500
rect 166166 143488 166172 143500
rect 166224 143488 166230 143540
rect 162762 143216 162768 143268
rect 162820 143256 162826 143268
rect 166074 143256 166080 143268
rect 162820 143228 166080 143256
rect 162820 143216 162826 143228
rect 166074 143216 166080 143228
rect 166132 143216 166138 143268
rect 137738 143148 137744 143200
rect 137796 143188 137802 143200
rect 139394 143188 139400 143200
rect 137796 143160 139400 143188
rect 137796 143148 137802 143160
rect 139394 143148 139400 143160
rect 139452 143148 139458 143200
rect 164234 142944 164240 142996
rect 164292 142984 164298 142996
rect 176194 142984 176200 142996
rect 164292 142956 176200 142984
rect 164292 142944 164298 142956
rect 176194 142944 176200 142956
rect 176252 142944 176258 142996
rect 150434 142876 150440 142928
rect 150492 142916 150498 142928
rect 154574 142916 154580 142928
rect 150492 142888 154580 142916
rect 150492 142876 150498 142888
rect 154574 142876 154580 142888
rect 154632 142876 154638 142928
rect 162854 142876 162860 142928
rect 162912 142916 162918 142928
rect 174630 142916 174636 142928
rect 162912 142888 174636 142916
rect 162912 142876 162918 142888
rect 174630 142876 174636 142888
rect 174688 142876 174694 142928
rect 163130 142808 163136 142860
rect 163188 142848 163194 142860
rect 178034 142848 178040 142860
rect 163188 142820 178040 142848
rect 163188 142808 163194 142820
rect 178034 142808 178040 142820
rect 178092 142808 178098 142860
rect 118234 142128 118240 142180
rect 118292 142168 118298 142180
rect 124858 142168 124864 142180
rect 118292 142140 124864 142168
rect 118292 142128 118298 142140
rect 124858 142128 124864 142140
rect 124916 142128 124922 142180
rect 149054 142128 149060 142180
rect 149112 142168 149118 142180
rect 152734 142168 152740 142180
rect 149112 142140 152740 142168
rect 149112 142128 149118 142140
rect 152734 142128 152740 142140
rect 152792 142128 152798 142180
rect 118142 141516 118148 141568
rect 118200 141556 118206 141568
rect 128998 141556 129004 141568
rect 118200 141528 129004 141556
rect 118200 141516 118206 141528
rect 128998 141516 129004 141528
rect 129056 141516 129062 141568
rect 118050 141448 118056 141500
rect 118108 141488 118114 141500
rect 169754 141488 169760 141500
rect 118108 141460 169760 141488
rect 118108 141448 118114 141460
rect 169754 141448 169760 141460
rect 169812 141448 169818 141500
rect 118970 141380 118976 141432
rect 119028 141420 119034 141432
rect 494054 141420 494060 141432
rect 119028 141392 494060 141420
rect 119028 141380 119034 141392
rect 494054 141380 494060 141392
rect 494112 141380 494118 141432
rect 118326 140224 118332 140276
rect 118384 140264 118390 140276
rect 126238 140264 126244 140276
rect 118384 140236 126244 140264
rect 118384 140224 118390 140236
rect 126238 140224 126244 140236
rect 126296 140224 126302 140276
rect 3878 140156 3884 140208
rect 3936 140196 3942 140208
rect 181438 140196 181444 140208
rect 3936 140168 181444 140196
rect 3936 140156 3942 140168
rect 181438 140156 181444 140168
rect 181496 140156 181502 140208
rect 119246 140088 119252 140140
rect 119304 140128 119310 140140
rect 364334 140128 364340 140140
rect 119304 140100 364340 140128
rect 119304 140088 119310 140100
rect 364334 140088 364340 140100
rect 364392 140088 364398 140140
rect 118786 140020 118792 140072
rect 118844 140060 118850 140072
rect 558914 140060 558920 140072
rect 118844 140032 558920 140060
rect 118844 140020 118850 140032
rect 558914 140020 558920 140032
rect 558972 140020 558978 140072
rect 118418 139476 118424 139528
rect 118476 139516 118482 139528
rect 122098 139516 122104 139528
rect 118476 139488 122104 139516
rect 118476 139476 118482 139488
rect 122098 139476 122104 139488
rect 122156 139476 122162 139528
rect 3510 139408 3516 139460
rect 3568 139448 3574 139460
rect 179506 139448 179512 139460
rect 3568 139420 179512 139448
rect 3568 139408 3574 139420
rect 179506 139408 179512 139420
rect 179564 139408 179570 139460
rect 178770 139340 178776 139392
rect 178828 139380 178834 139392
rect 182174 139380 182180 139392
rect 178828 139352 182180 139380
rect 178828 139340 178834 139352
rect 182174 139340 182180 139352
rect 182232 139340 182238 139392
rect 178678 139272 178684 139324
rect 178736 139312 178742 139324
rect 182450 139312 182456 139324
rect 178736 139284 182456 139312
rect 178736 139272 178742 139284
rect 182450 139272 182456 139284
rect 182508 139272 182514 139324
rect 193950 137980 193956 138032
rect 194008 138020 194014 138032
rect 580166 138020 580172 138032
rect 194008 137992 580172 138020
rect 194008 137980 194014 137992
rect 580166 137980 580172 137992
rect 580224 137980 580230 138032
rect 7650 136688 7656 136740
rect 7708 136728 7714 136740
rect 117314 136728 117320 136740
rect 7708 136700 117320 136728
rect 7708 136688 7714 136700
rect 117314 136688 117320 136700
rect 117372 136688 117378 136740
rect 2866 136620 2872 136672
rect 2924 136660 2930 136672
rect 115290 136660 115296 136672
rect 2924 136632 115296 136660
rect 2924 136620 2930 136632
rect 115290 136620 115296 136632
rect 115348 136620 115354 136672
rect 9030 135260 9036 135312
rect 9088 135300 9094 135312
rect 117314 135300 117320 135312
rect 9088 135272 117320 135300
rect 9088 135260 9094 135272
rect 117314 135260 117320 135272
rect 117372 135260 117378 135312
rect 21358 133900 21364 133952
rect 21416 133940 21422 133952
rect 117314 133940 117320 133952
rect 21416 133912 117320 133940
rect 21416 133900 21422 133912
rect 117314 133900 117320 133912
rect 117372 133900 117378 133952
rect 14458 133832 14464 133884
rect 14516 133872 14522 133884
rect 117406 133872 117412 133884
rect 14516 133844 117412 133872
rect 14516 133832 14522 133844
rect 117406 133832 117412 133844
rect 117464 133832 117470 133884
rect 31018 132404 31024 132456
rect 31076 132444 31082 132456
rect 117314 132444 117320 132456
rect 31076 132416 117320 132444
rect 31076 132404 31082 132416
rect 117314 132404 117320 132416
rect 117372 132404 117378 132456
rect 18598 131044 18604 131096
rect 18656 131084 18662 131096
rect 117314 131084 117320 131096
rect 18656 131056 117320 131084
rect 18656 131044 18662 131056
rect 117314 131044 117320 131056
rect 117372 131044 117378 131096
rect 13078 129684 13084 129736
rect 13136 129724 13142 129736
rect 117314 129724 117320 129736
rect 13136 129696 117320 129724
rect 13136 129684 13142 129696
rect 117314 129684 117320 129696
rect 117372 129684 117378 129736
rect 84838 128256 84844 128308
rect 84896 128296 84902 128308
rect 117314 128296 117320 128308
rect 84896 128268 117320 128296
rect 84896 128256 84902 128268
rect 117314 128256 117320 128268
rect 117372 128256 117378 128308
rect 10318 126896 10324 126948
rect 10376 126936 10382 126948
rect 117314 126936 117320 126948
rect 10376 126908 117320 126936
rect 10376 126896 10382 126908
rect 117314 126896 117320 126908
rect 117372 126896 117378 126948
rect 53098 124108 53104 124160
rect 53156 124148 53162 124160
rect 117314 124148 117320 124160
rect 53156 124120 117320 124148
rect 53156 124108 53162 124120
rect 117314 124108 117320 124120
rect 117372 124108 117378 124160
rect 8938 122748 8944 122800
rect 8996 122788 9002 122800
rect 117314 122788 117320 122800
rect 8996 122760 117320 122788
rect 8996 122748 9002 122760
rect 117314 122748 117320 122760
rect 117372 122748 117378 122800
rect 17218 121388 17224 121440
rect 17276 121428 17282 121440
rect 117314 121428 117320 121440
rect 17276 121400 117320 121428
rect 17276 121388 17282 121400
rect 117314 121388 117320 121400
rect 117372 121388 117378 121440
rect 7558 120028 7564 120080
rect 7616 120068 7622 120080
rect 117314 120068 117320 120080
rect 7616 120040 117320 120068
rect 7616 120028 7622 120040
rect 117314 120028 117320 120040
rect 117372 120028 117378 120080
rect 4798 118600 4804 118652
rect 4856 118640 4862 118652
rect 117314 118640 117320 118652
rect 4856 118612 117320 118640
rect 4856 118600 4862 118612
rect 117314 118600 117320 118612
rect 117372 118600 117378 118652
rect 40034 117240 40040 117292
rect 40092 117280 40098 117292
rect 117314 117280 117320 117292
rect 40092 117252 117320 117280
rect 40092 117240 40098 117252
rect 117314 117240 117320 117252
rect 117372 117240 117378 117292
rect 106918 115880 106924 115932
rect 106976 115920 106982 115932
rect 117314 115920 117320 115932
rect 106976 115892 117320 115920
rect 106976 115880 106982 115892
rect 117314 115880 117320 115892
rect 117372 115880 117378 115932
rect 180150 111800 180156 111852
rect 180208 111840 180214 111852
rect 580074 111840 580080 111852
rect 180208 111812 580080 111840
rect 180208 111800 180214 111812
rect 580074 111800 580080 111812
rect 580132 111800 580138 111852
rect 3326 111732 3332 111784
rect 3384 111772 3390 111784
rect 21358 111772 21364 111784
rect 3384 111744 21364 111772
rect 3384 111732 3390 111744
rect 21358 111732 21364 111744
rect 21416 111732 21422 111784
rect 183278 108944 183284 108996
rect 183336 108984 183342 108996
rect 196618 108984 196624 108996
rect 183336 108956 196624 108984
rect 183336 108944 183342 108956
rect 196618 108944 196624 108956
rect 196676 108944 196682 108996
rect 183278 107584 183284 107636
rect 183336 107624 183342 107636
rect 193858 107624 193864 107636
rect 183336 107596 193864 107624
rect 183336 107584 183342 107596
rect 193858 107584 193864 107596
rect 193916 107584 193922 107636
rect 183278 106224 183284 106276
rect 183336 106264 183342 106276
rect 192478 106264 192484 106276
rect 183336 106236 192484 106264
rect 183336 106224 183342 106236
rect 192478 106224 192484 106236
rect 192536 106224 192542 106276
rect 183278 104592 183284 104644
rect 183336 104632 183342 104644
rect 189718 104632 189724 104644
rect 183336 104604 189724 104632
rect 183336 104592 183342 104604
rect 189718 104592 189724 104604
rect 189776 104592 189782 104644
rect 183462 102892 183468 102944
rect 183520 102932 183526 102944
rect 188338 102932 188344 102944
rect 183520 102904 188344 102932
rect 183520 102892 183526 102904
rect 188338 102892 188344 102904
rect 188396 102892 188402 102944
rect 182634 101260 182640 101312
rect 182692 101300 182698 101312
rect 185578 101300 185584 101312
rect 182692 101272 185584 101300
rect 182692 101260 182698 101272
rect 185578 101260 185584 101272
rect 185636 101260 185642 101312
rect 182450 100444 182456 100496
rect 182508 100484 182514 100496
rect 184198 100484 184204 100496
rect 182508 100456 184204 100484
rect 182508 100444 182514 100456
rect 184198 100444 184204 100456
rect 184256 100444 184262 100496
rect 192478 99356 192484 99408
rect 192536 99396 192542 99408
rect 580074 99396 580080 99408
rect 192536 99368 580080 99396
rect 192536 99356 192542 99368
rect 580074 99356 580080 99368
rect 580132 99356 580138 99408
rect 182174 99288 182180 99340
rect 182232 99328 182238 99340
rect 184290 99328 184296 99340
rect 182232 99300 184296 99328
rect 182232 99288 182238 99300
rect 184290 99288 184296 99300
rect 184348 99288 184354 99340
rect 182174 97384 182180 97436
rect 182232 97424 182238 97436
rect 184382 97424 184388 97436
rect 182232 97396 184388 97424
rect 182232 97384 182238 97396
rect 184382 97384 184388 97396
rect 184440 97384 184446 97436
rect 183186 96568 183192 96620
rect 183244 96608 183250 96620
rect 214558 96608 214564 96620
rect 183244 96580 214564 96608
rect 183244 96568 183250 96580
rect 214558 96568 214564 96580
rect 214616 96568 214622 96620
rect 183462 95140 183468 95192
rect 183520 95180 183526 95192
rect 211798 95180 211804 95192
rect 183520 95152 211804 95180
rect 183520 95140 183526 95152
rect 211798 95140 211804 95152
rect 211856 95140 211862 95192
rect 183370 93100 183376 93152
rect 183428 93140 183434 93152
rect 224218 93140 224224 93152
rect 183428 93112 224224 93140
rect 183428 93100 183434 93112
rect 224218 93100 224224 93112
rect 224276 93100 224282 93152
rect 183462 91740 183468 91792
rect 183520 91780 183526 91792
rect 221458 91780 221464 91792
rect 183520 91752 221464 91780
rect 183520 91740 183526 91752
rect 221458 91740 221464 91752
rect 221516 91740 221522 91792
rect 183370 90312 183376 90364
rect 183428 90352 183434 90364
rect 220078 90352 220084 90364
rect 183428 90324 220084 90352
rect 183428 90312 183434 90324
rect 220078 90312 220084 90324
rect 220136 90312 220142 90364
rect 580074 89360 580080 89412
rect 580132 89400 580138 89412
rect 580534 89400 580540 89412
rect 580132 89372 580540 89400
rect 580132 89360 580138 89372
rect 580534 89360 580540 89372
rect 580592 89360 580598 89412
rect 580534 89224 580540 89276
rect 580592 89264 580598 89276
rect 580718 89264 580724 89276
rect 580592 89236 580724 89264
rect 580592 89224 580598 89236
rect 580718 89224 580724 89236
rect 580776 89224 580782 89276
rect 183462 88952 183468 89004
rect 183520 88992 183526 89004
rect 217318 88992 217324 89004
rect 183520 88964 217324 88992
rect 183520 88952 183526 88964
rect 217318 88952 217324 88964
rect 217376 88952 217382 89004
rect 183370 87592 183376 87644
rect 183428 87632 183434 87644
rect 215938 87632 215944 87644
rect 183428 87604 215944 87632
rect 183428 87592 183434 87604
rect 215938 87592 215944 87604
rect 215996 87592 216002 87644
rect 183462 85484 183468 85536
rect 183520 85524 183526 85536
rect 193950 85524 193956 85536
rect 183520 85496 193956 85524
rect 183520 85484 183526 85496
rect 193950 85484 193956 85496
rect 194008 85484 194014 85536
rect 183462 84124 183468 84176
rect 183520 84164 183526 84176
rect 192478 84164 192484 84176
rect 183520 84136 192484 84164
rect 183520 84124 183526 84136
rect 192478 84124 192484 84136
rect 192536 84124 192542 84176
rect 118602 80724 118608 80776
rect 118660 80764 118666 80776
rect 580902 80764 580908 80776
rect 118660 80736 171318 80764
rect 118660 80724 118666 80736
rect 171290 80696 171318 80736
rect 172348 80736 580908 80764
rect 172348 80696 172376 80736
rect 580902 80724 580908 80736
rect 580960 80724 580966 80776
rect 144886 80668 147674 80696
rect 135870 80464 137416 80492
rect 135870 80356 135898 80464
rect 137388 80424 137416 80464
rect 137388 80396 142154 80424
rect 122806 80328 135898 80356
rect 142126 80356 142154 80396
rect 144886 80356 144914 80668
rect 147646 80628 147674 80668
rect 154546 80668 171134 80696
rect 171290 80668 172376 80696
rect 147646 80600 150434 80628
rect 142126 80328 144914 80356
rect 150406 80356 150434 80600
rect 151786 80532 153194 80560
rect 151786 80356 151814 80532
rect 150406 80328 151814 80356
rect 121086 79976 121092 80028
rect 121144 80016 121150 80028
rect 122806 80016 122834 80328
rect 125410 80248 125416 80300
rect 125468 80288 125474 80300
rect 125468 80260 132678 80288
rect 125468 80248 125474 80260
rect 132650 80220 132678 80260
rect 140378 80260 142154 80288
rect 140378 80220 140406 80260
rect 132650 80192 140406 80220
rect 142126 80220 142154 80260
rect 143506 80260 144914 80288
rect 143506 80220 143534 80260
rect 142126 80192 143534 80220
rect 144886 80220 144914 80260
rect 146266 80260 147674 80288
rect 146266 80220 146294 80260
rect 144886 80192 146294 80220
rect 125226 80044 125232 80096
rect 125284 80084 125290 80096
rect 147646 80084 147674 80260
rect 153166 80220 153194 80532
rect 154546 80220 154574 80668
rect 171106 80628 171134 80668
rect 178586 80656 178592 80708
rect 178644 80696 178650 80708
rect 580810 80696 580816 80708
rect 178644 80668 580816 80696
rect 178644 80656 178650 80668
rect 580810 80656 580816 80668
rect 580868 80656 580874 80708
rect 174630 80628 174636 80640
rect 158778 80600 169754 80628
rect 171106 80600 174636 80628
rect 153166 80192 154574 80220
rect 155926 80328 158714 80356
rect 149026 80124 150434 80152
rect 149026 80084 149054 80124
rect 125284 80056 128630 80084
rect 147646 80056 149054 80084
rect 150406 80084 150434 80124
rect 150406 80056 153470 80084
rect 125284 80044 125290 80056
rect 121144 79988 122834 80016
rect 121144 79976 121150 79988
rect 123846 79976 123852 80028
rect 123904 80016 123910 80028
rect 123904 79988 127250 80016
rect 123904 79976 123910 79988
rect 127222 79960 127250 79988
rect 127498 79988 128078 80016
rect 127498 79960 127526 79988
rect 124950 79908 124956 79960
rect 125008 79948 125014 79960
rect 126100 79948 126106 79960
rect 125008 79920 126106 79948
rect 125008 79908 125014 79920
rect 126100 79908 126106 79920
rect 126158 79908 126164 79960
rect 126192 79908 126198 79960
rect 126250 79908 126256 79960
rect 126376 79908 126382 79960
rect 126434 79908 126440 79960
rect 126836 79908 126842 79960
rect 126894 79908 126900 79960
rect 127204 79908 127210 79960
rect 127262 79908 127268 79960
rect 127296 79908 127302 79960
rect 127354 79908 127360 79960
rect 127480 79908 127486 79960
rect 127538 79908 127544 79960
rect 127572 79908 127578 79960
rect 127630 79908 127636 79960
rect 127664 79908 127670 79960
rect 127722 79908 127728 79960
rect 127848 79948 127854 79960
rect 127820 79908 127854 79948
rect 127906 79908 127912 79960
rect 125824 79840 125830 79892
rect 125882 79840 125888 79892
rect 126008 79840 126014 79892
rect 126066 79840 126072 79892
rect 126210 79880 126238 79908
rect 126164 79852 126238 79880
rect 124766 79772 124772 79824
rect 124824 79812 124830 79824
rect 124824 79784 125594 79812
rect 124824 79772 124830 79784
rect 116578 79704 116584 79756
rect 116636 79744 116642 79756
rect 123570 79744 123576 79756
rect 116636 79716 123576 79744
rect 116636 79704 116642 79716
rect 123570 79704 123576 79716
rect 123628 79704 123634 79756
rect 125566 79688 125594 79784
rect 125732 79772 125738 79824
rect 125790 79772 125796 79824
rect 125750 79688 125778 79772
rect 121178 79636 121184 79688
rect 121236 79676 121242 79688
rect 125410 79676 125416 79688
rect 121236 79648 125416 79676
rect 121236 79636 121242 79648
rect 125410 79636 125416 79648
rect 125468 79636 125474 79688
rect 125566 79648 125600 79688
rect 125594 79636 125600 79648
rect 125652 79636 125658 79688
rect 125686 79636 125692 79688
rect 125744 79648 125778 79688
rect 125842 79676 125870 79840
rect 126026 79744 126054 79840
rect 126026 79716 126100 79744
rect 125962 79676 125968 79688
rect 125842 79648 125968 79676
rect 125744 79636 125750 79648
rect 125962 79636 125968 79648
rect 126020 79636 126026 79688
rect 126072 79620 126100 79716
rect 126164 79620 126192 79852
rect 126284 79840 126290 79892
rect 126342 79840 126348 79892
rect 126302 79812 126330 79840
rect 126256 79784 126330 79812
rect 126256 79756 126284 79784
rect 126394 79756 126422 79908
rect 126238 79704 126244 79756
rect 126296 79704 126302 79756
rect 126330 79704 126336 79756
rect 126388 79716 126422 79756
rect 126388 79704 126394 79716
rect 126854 79688 126882 79908
rect 127020 79772 127026 79824
rect 127078 79772 127084 79824
rect 127038 79688 127066 79772
rect 127314 79756 127342 79908
rect 127590 79824 127618 79908
rect 127572 79772 127578 79824
rect 127630 79772 127636 79824
rect 127250 79704 127256 79756
rect 127308 79716 127342 79756
rect 127308 79704 127314 79716
rect 126854 79648 126888 79688
rect 126882 79636 126888 79648
rect 126940 79636 126946 79688
rect 126974 79636 126980 79688
rect 127032 79648 127066 79688
rect 127032 79636 127038 79648
rect 127158 79636 127164 79688
rect 127216 79676 127222 79688
rect 127682 79676 127710 79908
rect 127216 79648 127710 79676
rect 127820 79676 127848 79908
rect 127940 79880 127946 79892
rect 127912 79840 127946 79880
rect 127998 79840 128004 79892
rect 127912 79756 127940 79840
rect 128050 79812 128078 79988
rect 128602 79960 128630 80056
rect 128694 79988 129274 80016
rect 128124 79908 128130 79960
rect 128182 79908 128188 79960
rect 128584 79908 128590 79960
rect 128642 79908 128648 79960
rect 128004 79784 128078 79812
rect 128004 79756 128032 79784
rect 128142 79756 128170 79908
rect 128694 79880 128722 79988
rect 129246 79960 129274 79988
rect 130350 79988 130608 80016
rect 130350 79960 130378 79988
rect 128768 79908 128774 79960
rect 128826 79908 128832 79960
rect 128860 79908 128866 79960
rect 128918 79908 128924 79960
rect 128952 79908 128958 79960
rect 129010 79908 129016 79960
rect 129228 79908 129234 79960
rect 129286 79908 129292 79960
rect 130148 79908 130154 79960
rect 130206 79908 130212 79960
rect 130240 79908 130246 79960
rect 130298 79908 130304 79960
rect 130332 79908 130338 79960
rect 130390 79908 130396 79960
rect 130424 79908 130430 79960
rect 130482 79948 130488 79960
rect 130482 79908 130516 79948
rect 128648 79852 128722 79880
rect 128648 79824 128676 79852
rect 128786 79824 128814 79908
rect 128400 79772 128406 79824
rect 128458 79772 128464 79824
rect 128630 79772 128636 79824
rect 128688 79772 128694 79824
rect 128722 79772 128728 79824
rect 128780 79784 128814 79824
rect 128780 79772 128786 79784
rect 127894 79704 127900 79756
rect 127952 79704 127958 79756
rect 127986 79704 127992 79756
rect 128044 79704 128050 79756
rect 128078 79704 128084 79756
rect 128136 79716 128170 79756
rect 128418 79744 128446 79772
rect 128878 79756 128906 79908
rect 128418 79716 128492 79744
rect 128136 79704 128142 79716
rect 128464 79688 128492 79716
rect 128814 79704 128820 79756
rect 128872 79716 128906 79756
rect 128872 79704 128878 79716
rect 128354 79676 128360 79688
rect 127820 79648 128360 79676
rect 127216 79636 127222 79648
rect 128354 79636 128360 79648
rect 128412 79636 128418 79688
rect 128446 79636 128452 79688
rect 128504 79636 128510 79688
rect 86218 79568 86224 79620
rect 86276 79608 86282 79620
rect 86276 79580 123616 79608
rect 86276 79568 86282 79580
rect 115290 79432 115296 79484
rect 115348 79472 115354 79484
rect 115348 79444 123524 79472
rect 115348 79432 115354 79444
rect 71774 79364 71780 79416
rect 71832 79404 71838 79416
rect 71832 79376 123432 79404
rect 71832 79364 71838 79376
rect 3970 79296 3976 79348
rect 4028 79336 4034 79348
rect 4028 79308 118694 79336
rect 4028 79296 4034 79308
rect 118666 79132 118694 79308
rect 123404 79200 123432 79376
rect 123496 79268 123524 79444
rect 123588 79404 123616 79580
rect 126054 79568 126060 79620
rect 126112 79568 126118 79620
rect 126146 79568 126152 79620
rect 126204 79568 126210 79620
rect 128970 79552 128998 79908
rect 129136 79840 129142 79892
rect 129194 79880 129200 79892
rect 129194 79840 129228 79880
rect 129780 79840 129786 79892
rect 129838 79840 129844 79892
rect 129200 79688 129228 79840
rect 129596 79772 129602 79824
rect 129654 79772 129660 79824
rect 129614 79688 129642 79772
rect 129182 79636 129188 79688
rect 129240 79636 129246 79688
rect 129550 79636 129556 79688
rect 129608 79648 129642 79688
rect 129608 79636 129614 79648
rect 129274 79568 129280 79620
rect 129332 79608 129338 79620
rect 129458 79608 129464 79620
rect 129332 79580 129464 79608
rect 129332 79568 129338 79580
rect 129458 79568 129464 79580
rect 129516 79568 129522 79620
rect 129798 79608 129826 79840
rect 130166 79756 130194 79908
rect 130258 79812 130286 79908
rect 130258 79784 130332 79812
rect 130304 79756 130332 79784
rect 130166 79716 130200 79756
rect 130194 79704 130200 79716
rect 130252 79704 130258 79756
rect 130286 79704 130292 79756
rect 130344 79704 130350 79756
rect 129752 79580 129826 79608
rect 129752 79552 129780 79580
rect 128906 79500 128912 79552
rect 128964 79512 128998 79552
rect 128964 79500 128970 79512
rect 129090 79500 129096 79552
rect 129148 79500 129154 79552
rect 129734 79500 129740 79552
rect 129792 79500 129798 79552
rect 125502 79432 125508 79484
rect 125560 79472 125566 79484
rect 129108 79472 129136 79500
rect 130488 79472 130516 79908
rect 130580 79620 130608 79988
rect 132420 79988 133966 80016
rect 130884 79908 130890 79960
rect 130942 79908 130948 79960
rect 131712 79908 131718 79960
rect 131770 79908 131776 79960
rect 131988 79908 131994 79960
rect 132046 79908 132052 79960
rect 132264 79908 132270 79960
rect 132322 79948 132328 79960
rect 132322 79908 132356 79948
rect 130700 79812 130706 79824
rect 130672 79772 130706 79812
rect 130758 79772 130764 79824
rect 130672 79688 130700 79772
rect 130654 79636 130660 79688
rect 130712 79636 130718 79688
rect 130562 79568 130568 79620
rect 130620 79568 130626 79620
rect 130902 79552 130930 79908
rect 131068 79880 131074 79892
rect 131040 79840 131074 79880
rect 131126 79880 131132 79892
rect 131126 79852 131173 79880
rect 131126 79840 131132 79852
rect 131040 79756 131068 79840
rect 131022 79704 131028 79756
rect 131080 79704 131086 79756
rect 131730 79676 131758 79908
rect 131850 79676 131856 79688
rect 131730 79648 131856 79676
rect 131850 79636 131856 79648
rect 131908 79636 131914 79688
rect 131298 79568 131304 79620
rect 131356 79608 131362 79620
rect 132006 79608 132034 79908
rect 132328 79756 132356 79908
rect 132310 79704 132316 79756
rect 132368 79704 132374 79756
rect 131356 79580 132034 79608
rect 131356 79568 131362 79580
rect 130838 79500 130844 79552
rect 130896 79512 130930 79552
rect 130896 79500 130902 79512
rect 132218 79500 132224 79552
rect 132276 79540 132282 79552
rect 132420 79540 132448 79988
rect 133938 79960 133966 79988
rect 134030 79988 135898 80016
rect 132908 79948 132914 79960
rect 132276 79512 132448 79540
rect 132512 79920 132914 79948
rect 132276 79500 132282 79512
rect 125560 79444 129136 79472
rect 129844 79444 130516 79472
rect 125560 79432 125566 79444
rect 129844 79416 129872 79444
rect 130930 79432 130936 79484
rect 130988 79472 130994 79484
rect 132512 79472 132540 79920
rect 132908 79908 132914 79920
rect 132966 79908 132972 79960
rect 133184 79908 133190 79960
rect 133242 79948 133248 79960
rect 133242 79908 133276 79948
rect 133920 79908 133926 79960
rect 133978 79908 133984 79960
rect 133248 79744 133276 79908
rect 133736 79880 133742 79892
rect 132880 79716 133276 79744
rect 133340 79852 133742 79880
rect 132880 79688 132908 79716
rect 132862 79636 132868 79688
rect 132920 79636 132926 79688
rect 132954 79568 132960 79620
rect 133012 79608 133018 79620
rect 133340 79608 133368 79852
rect 133736 79840 133742 79852
rect 133794 79840 133800 79892
rect 134030 79824 134058 79988
rect 134656 79908 134662 79960
rect 134714 79908 134720 79960
rect 134840 79908 134846 79960
rect 134898 79908 134904 79960
rect 135116 79908 135122 79960
rect 135174 79908 135180 79960
rect 135392 79908 135398 79960
rect 135450 79908 135456 79960
rect 135576 79908 135582 79960
rect 135634 79908 135640 79960
rect 135870 79948 135898 79988
rect 144242 79988 150112 80016
rect 144242 79960 144270 79988
rect 135944 79948 135950 79960
rect 135870 79920 135950 79948
rect 135944 79908 135950 79920
rect 136002 79908 136008 79960
rect 137232 79908 137238 79960
rect 137290 79908 137296 79960
rect 137600 79908 137606 79960
rect 137658 79908 137664 79960
rect 138520 79948 138526 79960
rect 138216 79920 138526 79948
rect 134196 79840 134202 79892
rect 134254 79840 134260 79892
rect 133966 79772 133972 79824
rect 134024 79784 134058 79824
rect 134024 79772 134030 79784
rect 134214 79676 134242 79840
rect 134674 79824 134702 79908
rect 134674 79784 134708 79824
rect 134702 79772 134708 79784
rect 134760 79772 134766 79824
rect 133524 79648 134242 79676
rect 133524 79620 133552 79648
rect 133012 79580 133368 79608
rect 133012 79568 133018 79580
rect 133506 79568 133512 79620
rect 133564 79568 133570 79620
rect 133782 79568 133788 79620
rect 133840 79608 133846 79620
rect 134858 79608 134886 79908
rect 133840 79580 134886 79608
rect 133840 79568 133846 79580
rect 133322 79500 133328 79552
rect 133380 79540 133386 79552
rect 135134 79540 135162 79908
rect 135300 79840 135306 79892
rect 135358 79840 135364 79892
rect 135318 79688 135346 79840
rect 135410 79744 135438 79908
rect 135410 79716 135484 79744
rect 135318 79648 135352 79688
rect 135346 79636 135352 79648
rect 135404 79636 135410 79688
rect 133380 79512 135162 79540
rect 133380 79500 133386 79512
rect 135254 79500 135260 79552
rect 135312 79540 135318 79552
rect 135456 79540 135484 79716
rect 135594 79552 135622 79908
rect 135760 79840 135766 79892
rect 135818 79840 135824 79892
rect 136036 79840 136042 79892
rect 136094 79880 136100 79892
rect 136094 79840 136128 79880
rect 136680 79840 136686 79892
rect 136738 79840 136744 79892
rect 136864 79840 136870 79892
rect 136922 79840 136928 79892
rect 135778 79756 135806 79840
rect 135714 79704 135720 79756
rect 135772 79716 135806 79756
rect 135772 79704 135778 79716
rect 135312 79512 135484 79540
rect 135312 79500 135318 79512
rect 135530 79500 135536 79552
rect 135588 79512 135622 79552
rect 135588 79500 135594 79512
rect 134794 79472 134800 79484
rect 130988 79444 132540 79472
rect 132696 79444 134800 79472
rect 130988 79432 130994 79444
rect 129090 79404 129096 79416
rect 123588 79376 129096 79404
rect 129090 79364 129096 79376
rect 129148 79364 129154 79416
rect 129826 79364 129832 79416
rect 129884 79364 129890 79416
rect 130102 79364 130108 79416
rect 130160 79404 130166 79416
rect 132696 79404 132724 79444
rect 134794 79432 134800 79444
rect 134852 79432 134858 79484
rect 130160 79376 132724 79404
rect 130160 79364 130166 79376
rect 132770 79364 132776 79416
rect 132828 79404 132834 79416
rect 133874 79404 133880 79416
rect 132828 79376 133880 79404
rect 132828 79364 132834 79376
rect 133874 79364 133880 79376
rect 133932 79364 133938 79416
rect 135990 79364 135996 79416
rect 136048 79404 136054 79416
rect 136100 79404 136128 79840
rect 136698 79540 136726 79840
rect 136882 79688 136910 79840
rect 136818 79636 136824 79688
rect 136876 79648 136910 79688
rect 136876 79636 136882 79648
rect 137002 79568 137008 79620
rect 137060 79608 137066 79620
rect 137250 79608 137278 79908
rect 137060 79580 137278 79608
rect 137618 79608 137646 79908
rect 138216 79620 138244 79920
rect 138520 79908 138526 79920
rect 138578 79908 138584 79960
rect 138704 79948 138710 79960
rect 138676 79908 138710 79948
rect 138762 79908 138768 79960
rect 138888 79908 138894 79960
rect 138946 79908 138952 79960
rect 139072 79908 139078 79960
rect 139130 79908 139136 79960
rect 139440 79908 139446 79960
rect 139498 79948 139504 79960
rect 139498 79920 139624 79948
rect 139498 79908 139504 79920
rect 138336 79840 138342 79892
rect 138394 79880 138400 79892
rect 138394 79852 138612 79880
rect 138394 79840 138400 79852
rect 138584 79824 138612 79852
rect 138676 79824 138704 79908
rect 138566 79772 138572 79824
rect 138624 79772 138630 79824
rect 138658 79772 138664 79824
rect 138716 79772 138722 79824
rect 138796 79772 138802 79824
rect 138854 79772 138860 79824
rect 138814 79744 138842 79772
rect 138768 79716 138842 79744
rect 138768 79688 138796 79716
rect 138906 79688 138934 79908
rect 139090 79756 139118 79908
rect 139164 79840 139170 79892
rect 139222 79840 139228 79892
rect 139026 79704 139032 79756
rect 139084 79716 139118 79756
rect 139084 79704 139090 79716
rect 138750 79636 138756 79688
rect 138808 79636 138814 79688
rect 138842 79636 138848 79688
rect 138900 79648 138934 79688
rect 138900 79636 138906 79648
rect 137830 79608 137836 79620
rect 137618 79580 137836 79608
rect 137060 79568 137066 79580
rect 137830 79568 137836 79580
rect 137888 79568 137894 79620
rect 138198 79568 138204 79620
rect 138256 79568 138262 79620
rect 138934 79568 138940 79620
rect 138992 79608 138998 79620
rect 139182 79608 139210 79840
rect 139596 79744 139624 79920
rect 139900 79908 139906 79960
rect 139958 79908 139964 79960
rect 140360 79908 140366 79960
rect 140418 79948 140424 79960
rect 141280 79948 141286 79960
rect 140418 79920 140636 79948
rect 140418 79908 140424 79920
rect 139918 79880 139946 79908
rect 139504 79716 139624 79744
rect 139688 79852 139946 79880
rect 139504 79688 139532 79716
rect 139486 79636 139492 79688
rect 139544 79636 139550 79688
rect 138992 79580 139210 79608
rect 138992 79568 138998 79580
rect 139688 79552 139716 79852
rect 140084 79840 140090 79892
rect 140142 79840 140148 79892
rect 140268 79840 140274 79892
rect 140326 79840 140332 79892
rect 137462 79540 137468 79552
rect 136698 79512 137468 79540
rect 137462 79500 137468 79512
rect 137520 79500 137526 79552
rect 139670 79500 139676 79552
rect 139728 79500 139734 79552
rect 140102 79484 140130 79840
rect 140286 79552 140314 79840
rect 140286 79512 140320 79552
rect 140314 79500 140320 79512
rect 140372 79500 140378 79552
rect 140498 79500 140504 79552
rect 140556 79540 140562 79552
rect 140608 79540 140636 79920
rect 140556 79512 140636 79540
rect 140792 79920 141286 79948
rect 140792 79540 140820 79920
rect 141280 79908 141286 79920
rect 141338 79908 141344 79960
rect 141556 79908 141562 79960
rect 141614 79948 141620 79960
rect 141614 79920 141878 79948
rect 141614 79908 141620 79920
rect 140912 79880 140918 79892
rect 140884 79840 140918 79880
rect 140970 79840 140976 79892
rect 141004 79840 141010 79892
rect 141062 79840 141068 79892
rect 141096 79840 141102 79892
rect 141154 79840 141160 79892
rect 141464 79840 141470 79892
rect 141522 79840 141528 79892
rect 141740 79840 141746 79892
rect 141798 79840 141804 79892
rect 140884 79608 140912 79840
rect 141022 79688 141050 79840
rect 140958 79636 140964 79688
rect 141016 79648 141050 79688
rect 141114 79676 141142 79840
rect 141482 79756 141510 79840
rect 141482 79716 141516 79756
rect 141510 79704 141516 79716
rect 141568 79704 141574 79756
rect 141114 79648 141280 79676
rect 141016 79636 141022 79648
rect 141142 79608 141148 79620
rect 140884 79580 141148 79608
rect 141142 79568 141148 79580
rect 141200 79568 141206 79620
rect 140958 79540 140964 79552
rect 140792 79512 140964 79540
rect 140556 79500 140562 79512
rect 140958 79500 140964 79512
rect 141016 79500 141022 79552
rect 140038 79432 140044 79484
rect 140096 79444 140130 79484
rect 141252 79472 141280 79648
rect 141326 79568 141332 79620
rect 141384 79608 141390 79620
rect 141758 79608 141786 79840
rect 141384 79580 141786 79608
rect 141384 79568 141390 79580
rect 141694 79500 141700 79552
rect 141752 79540 141758 79552
rect 141850 79540 141878 79920
rect 142476 79908 142482 79960
rect 142534 79908 142540 79960
rect 142568 79908 142574 79960
rect 142626 79908 142632 79960
rect 142752 79908 142758 79960
rect 142810 79908 142816 79960
rect 142844 79908 142850 79960
rect 142902 79908 142908 79960
rect 142936 79908 142942 79960
rect 142994 79908 143000 79960
rect 143028 79908 143034 79960
rect 143086 79908 143092 79960
rect 144132 79908 144138 79960
rect 144190 79908 144196 79960
rect 144224 79908 144230 79960
rect 144282 79908 144288 79960
rect 144316 79908 144322 79960
rect 144374 79908 144380 79960
rect 144408 79908 144414 79960
rect 144466 79908 144472 79960
rect 144592 79908 144598 79960
rect 144650 79908 144656 79960
rect 144684 79908 144690 79960
rect 144742 79908 144748 79960
rect 145696 79948 145702 79960
rect 144932 79920 145702 79948
rect 142200 79840 142206 79892
rect 142258 79840 142264 79892
rect 142218 79620 142246 79840
rect 142494 79756 142522 79908
rect 142586 79812 142614 79908
rect 142586 79784 142660 79812
rect 142494 79716 142528 79756
rect 142522 79704 142528 79716
rect 142580 79704 142586 79756
rect 142218 79580 142252 79620
rect 142246 79568 142252 79580
rect 142304 79568 142310 79620
rect 141752 79512 141878 79540
rect 141752 79500 141758 79512
rect 142338 79500 142344 79552
rect 142396 79540 142402 79552
rect 142632 79540 142660 79784
rect 142770 79620 142798 79908
rect 142706 79568 142712 79620
rect 142764 79580 142798 79620
rect 142764 79568 142770 79580
rect 142396 79512 142660 79540
rect 142396 79500 142402 79512
rect 141878 79472 141884 79484
rect 141252 79444 141884 79472
rect 140096 79432 140102 79444
rect 141878 79432 141884 79444
rect 141936 79432 141942 79484
rect 142154 79432 142160 79484
rect 142212 79472 142218 79484
rect 142862 79472 142890 79908
rect 142954 79540 142982 79908
rect 143046 79620 143074 79908
rect 143856 79840 143862 79892
rect 143914 79840 143920 79892
rect 144150 79880 144178 79908
rect 144150 79852 144224 79880
rect 143304 79772 143310 79824
rect 143362 79772 143368 79824
rect 143396 79772 143402 79824
rect 143454 79772 143460 79824
rect 143580 79772 143586 79824
rect 143638 79772 143644 79824
rect 143672 79772 143678 79824
rect 143730 79772 143736 79824
rect 143322 79688 143350 79772
rect 143258 79636 143264 79688
rect 143316 79648 143350 79688
rect 143316 79636 143322 79648
rect 143414 79620 143442 79772
rect 143598 79744 143626 79772
rect 143552 79716 143626 79744
rect 143552 79688 143580 79716
rect 143534 79636 143540 79688
rect 143592 79636 143598 79688
rect 143046 79580 143080 79620
rect 143074 79568 143080 79580
rect 143132 79568 143138 79620
rect 143414 79580 143448 79620
rect 143442 79568 143448 79580
rect 143500 79568 143506 79620
rect 143690 79608 143718 79772
rect 143874 79744 143902 79840
rect 143948 79772 143954 79824
rect 144006 79812 144012 79824
rect 144006 79772 144040 79812
rect 144012 79744 144040 79772
rect 143874 79716 143948 79744
rect 144012 79716 144132 79744
rect 143920 79676 143948 79716
rect 143994 79676 144000 79688
rect 143920 79648 144000 79676
rect 143994 79636 144000 79648
rect 144052 79636 144058 79688
rect 144104 79620 144132 79716
rect 144196 79688 144224 79852
rect 144178 79636 144184 79688
rect 144236 79636 144242 79688
rect 143644 79580 143718 79608
rect 143350 79540 143356 79552
rect 142954 79512 143356 79540
rect 143350 79500 143356 79512
rect 143408 79500 143414 79552
rect 142212 79444 142890 79472
rect 143644 79472 143672 79580
rect 144086 79568 144092 79620
rect 144144 79568 144150 79620
rect 143718 79500 143724 79552
rect 143776 79540 143782 79552
rect 144334 79540 144362 79908
rect 144426 79676 144454 79908
rect 144426 79648 144500 79676
rect 143776 79512 144362 79540
rect 143776 79500 143782 79512
rect 143810 79472 143816 79484
rect 143644 79444 143816 79472
rect 142212 79432 142218 79444
rect 143810 79432 143816 79444
rect 143868 79432 143874 79484
rect 144362 79432 144368 79484
rect 144420 79472 144426 79484
rect 144472 79472 144500 79648
rect 144420 79444 144500 79472
rect 144610 79472 144638 79908
rect 144702 79620 144730 79908
rect 144702 79580 144736 79620
rect 144730 79568 144736 79580
rect 144788 79568 144794 79620
rect 144932 79552 144960 79920
rect 145696 79908 145702 79920
rect 145754 79908 145760 79960
rect 145788 79908 145794 79960
rect 145846 79908 145852 79960
rect 146248 79908 146254 79960
rect 146306 79908 146312 79960
rect 146340 79908 146346 79960
rect 146398 79908 146404 79960
rect 147168 79948 147174 79960
rect 146726 79920 147174 79948
rect 145144 79840 145150 79892
rect 145202 79840 145208 79892
rect 145236 79840 145242 79892
rect 145294 79840 145300 79892
rect 144914 79500 144920 79552
rect 144972 79500 144978 79552
rect 145162 79540 145190 79840
rect 145254 79688 145282 79840
rect 145806 79824 145834 79908
rect 145742 79772 145748 79824
rect 145800 79784 145834 79824
rect 145800 79772 145806 79784
rect 146266 79756 146294 79908
rect 146358 79812 146386 79908
rect 146432 79840 146438 79892
rect 146490 79880 146496 79892
rect 146490 79840 146524 79880
rect 146358 79784 146432 79812
rect 146266 79716 146300 79756
rect 146294 79704 146300 79716
rect 146352 79704 146358 79756
rect 145254 79648 145288 79688
rect 145282 79636 145288 79648
rect 145340 79636 145346 79688
rect 146110 79636 146116 79688
rect 146168 79676 146174 79688
rect 146404 79676 146432 79784
rect 146168 79648 146432 79676
rect 146168 79636 146174 79648
rect 146386 79568 146392 79620
rect 146444 79608 146450 79620
rect 146496 79608 146524 79840
rect 146726 79620 146754 79920
rect 147168 79908 147174 79920
rect 147226 79908 147232 79960
rect 147352 79908 147358 79960
rect 147410 79908 147416 79960
rect 147444 79908 147450 79960
rect 147502 79908 147508 79960
rect 147536 79908 147542 79960
rect 147594 79908 147600 79960
rect 147628 79908 147634 79960
rect 147686 79948 147692 79960
rect 147686 79920 149008 79948
rect 147686 79908 147692 79920
rect 146984 79840 146990 79892
rect 147042 79840 147048 79892
rect 147370 79880 147398 79908
rect 147324 79852 147398 79880
rect 146800 79772 146806 79824
rect 146858 79772 146864 79824
rect 146818 79688 146846 79772
rect 146818 79648 146852 79688
rect 146846 79636 146852 79648
rect 146904 79636 146910 79688
rect 147002 79620 147030 79840
rect 147324 79688 147352 79852
rect 147462 79812 147490 79908
rect 147416 79784 147490 79812
rect 147416 79688 147444 79784
rect 147554 79756 147582 79908
rect 148272 79880 148278 79892
rect 147490 79704 147496 79756
rect 147548 79716 147582 79756
rect 147692 79852 148278 79880
rect 147548 79704 147554 79716
rect 147306 79636 147312 79688
rect 147364 79636 147370 79688
rect 147398 79636 147404 79688
rect 147456 79636 147462 79688
rect 146444 79580 146524 79608
rect 146444 79568 146450 79580
rect 146662 79568 146668 79620
rect 146720 79580 146754 79620
rect 146720 79568 146726 79580
rect 146938 79568 146944 79620
rect 146996 79580 147030 79620
rect 146996 79568 147002 79580
rect 147692 79552 147720 79852
rect 148272 79840 148278 79852
rect 148330 79840 148336 79892
rect 148364 79840 148370 79892
rect 148422 79840 148428 79892
rect 147904 79772 147910 79824
rect 147962 79812 147968 79824
rect 147962 79784 148180 79812
rect 147962 79772 147968 79784
rect 148152 79620 148180 79784
rect 148382 79756 148410 79840
rect 148318 79704 148324 79756
rect 148376 79716 148410 79756
rect 148376 79704 148382 79716
rect 148980 79688 149008 79920
rect 149192 79908 149198 79960
rect 149250 79908 149256 79960
rect 149284 79908 149290 79960
rect 149342 79908 149348 79960
rect 149560 79908 149566 79960
rect 149618 79948 149624 79960
rect 149618 79920 150020 79948
rect 149618 79908 149624 79920
rect 149210 79744 149238 79908
rect 149164 79716 149238 79744
rect 148962 79636 148968 79688
rect 149020 79636 149026 79688
rect 148134 79568 148140 79620
rect 148192 79568 148198 79620
rect 147214 79540 147220 79552
rect 145162 79512 147220 79540
rect 147214 79500 147220 79512
rect 147272 79500 147278 79552
rect 147674 79500 147680 79552
rect 147732 79500 147738 79552
rect 149164 79540 149192 79716
rect 149302 79620 149330 79908
rect 149376 79840 149382 79892
rect 149434 79840 149440 79892
rect 149468 79840 149474 79892
rect 149526 79840 149532 79892
rect 149836 79840 149842 79892
rect 149894 79840 149900 79892
rect 149394 79676 149422 79840
rect 149486 79744 149514 79840
rect 149486 79716 149698 79744
rect 149514 79676 149520 79688
rect 149394 79648 149520 79676
rect 149514 79636 149520 79648
rect 149572 79636 149578 79688
rect 149238 79568 149244 79620
rect 149296 79580 149330 79620
rect 149296 79568 149302 79580
rect 149422 79540 149428 79552
rect 149164 79512 149428 79540
rect 149422 79500 149428 79512
rect 149480 79500 149486 79552
rect 148502 79472 148508 79484
rect 144610 79444 148508 79472
rect 144420 79432 144426 79444
rect 148502 79432 148508 79444
rect 148560 79432 148566 79484
rect 136048 79376 136128 79404
rect 136048 79364 136054 79376
rect 149054 79364 149060 79416
rect 149112 79404 149118 79416
rect 149670 79404 149698 79716
rect 149854 79688 149882 79840
rect 149790 79636 149796 79688
rect 149848 79648 149882 79688
rect 149848 79636 149854 79648
rect 149992 79620 150020 79920
rect 149974 79568 149980 79620
rect 150032 79568 150038 79620
rect 150084 79608 150112 79988
rect 151970 79988 152366 80016
rect 151970 79960 151998 79988
rect 151124 79908 151130 79960
rect 151182 79908 151188 79960
rect 151492 79908 151498 79960
rect 151550 79908 151556 79960
rect 151584 79908 151590 79960
rect 151642 79908 151648 79960
rect 151952 79908 151958 79960
rect 152010 79908 152016 79960
rect 150664 79880 150670 79892
rect 150452 79852 150670 79880
rect 150250 79608 150256 79620
rect 150084 79580 150256 79608
rect 150250 79568 150256 79580
rect 150308 79568 150314 79620
rect 150452 79552 150480 79852
rect 150664 79840 150670 79852
rect 150722 79840 150728 79892
rect 150848 79840 150854 79892
rect 150906 79840 150912 79892
rect 150866 79812 150894 79840
rect 150636 79784 150894 79812
rect 150636 79552 150664 79784
rect 150434 79500 150440 79552
rect 150492 79500 150498 79552
rect 150618 79500 150624 79552
rect 150676 79500 150682 79552
rect 151142 79472 151170 79908
rect 151216 79840 151222 79892
rect 151274 79840 151280 79892
rect 151308 79840 151314 79892
rect 151366 79880 151372 79892
rect 151510 79880 151538 79908
rect 151366 79840 151400 79880
rect 151234 79756 151262 79840
rect 151234 79716 151268 79756
rect 151262 79704 151268 79716
rect 151320 79704 151326 79756
rect 151372 79620 151400 79840
rect 151464 79852 151538 79880
rect 151354 79568 151360 79620
rect 151412 79568 151418 79620
rect 151464 79608 151492 79852
rect 151602 79824 151630 79908
rect 152228 79880 152234 79892
rect 152200 79840 152234 79880
rect 152286 79840 152292 79892
rect 151538 79772 151544 79824
rect 151596 79784 151630 79824
rect 151596 79772 151602 79784
rect 151860 79772 151866 79824
rect 151918 79772 151924 79824
rect 151630 79704 151636 79756
rect 151688 79744 151694 79756
rect 151878 79744 151906 79772
rect 151688 79716 151814 79744
rect 151878 79716 152136 79744
rect 151688 79704 151694 79716
rect 151786 79676 151814 79716
rect 151998 79676 152004 79688
rect 151786 79648 152004 79676
rect 151998 79636 152004 79648
rect 152056 79636 152062 79688
rect 151906 79608 151912 79620
rect 151464 79580 151912 79608
rect 151906 79568 151912 79580
rect 151964 79568 151970 79620
rect 151262 79472 151268 79484
rect 151142 79444 151268 79472
rect 151262 79432 151268 79444
rect 151320 79432 151326 79484
rect 152108 79416 152136 79716
rect 149112 79376 149698 79404
rect 149112 79364 149118 79376
rect 152090 79364 152096 79416
rect 152148 79364 152154 79416
rect 123570 79296 123576 79348
rect 123628 79336 123634 79348
rect 123628 79308 150434 79336
rect 123628 79296 123634 79308
rect 123496 79240 128354 79268
rect 125594 79200 125600 79212
rect 123404 79172 125600 79200
rect 125594 79160 125600 79172
rect 125652 79160 125658 79212
rect 127618 79160 127624 79212
rect 127676 79200 127682 79212
rect 128078 79200 128084 79212
rect 127676 79172 128084 79200
rect 127676 79160 127682 79172
rect 128078 79160 128084 79172
rect 128136 79160 128142 79212
rect 128326 79200 128354 79240
rect 129642 79228 129648 79280
rect 129700 79268 129706 79280
rect 133506 79268 133512 79280
rect 129700 79240 133512 79268
rect 129700 79228 129706 79240
rect 133506 79228 133512 79240
rect 133564 79228 133570 79280
rect 133874 79228 133880 79280
rect 133932 79268 133938 79280
rect 133932 79240 145604 79268
rect 133932 79228 133938 79240
rect 145466 79200 145472 79212
rect 128326 79172 145472 79200
rect 145466 79160 145472 79172
rect 145524 79160 145530 79212
rect 145576 79132 145604 79240
rect 150406 79200 150434 79308
rect 151906 79296 151912 79348
rect 151964 79336 151970 79348
rect 152200 79336 152228 79840
rect 152338 79812 152366 79988
rect 152614 79988 153194 80016
rect 152504 79908 152510 79960
rect 152562 79908 152568 79960
rect 152292 79784 152366 79812
rect 152292 79688 152320 79784
rect 152366 79704 152372 79756
rect 152424 79704 152430 79756
rect 152274 79636 152280 79688
rect 152332 79636 152338 79688
rect 152384 79608 152412 79704
rect 152522 79688 152550 79908
rect 152614 79892 152642 79988
rect 152688 79908 152694 79960
rect 152746 79908 152752 79960
rect 153166 79948 153194 79988
rect 153166 79920 153240 79948
rect 152596 79840 152602 79892
rect 152654 79840 152660 79892
rect 152706 79756 152734 79908
rect 152964 79772 152970 79824
rect 153022 79772 153028 79824
rect 152642 79704 152648 79756
rect 152700 79716 152734 79756
rect 152700 79704 152706 79716
rect 152522 79648 152556 79688
rect 152550 79636 152556 79648
rect 152608 79636 152614 79688
rect 152384 79580 152872 79608
rect 152844 79552 152872 79580
rect 152982 79552 153010 79772
rect 153212 79744 153240 79920
rect 153332 79908 153338 79960
rect 153390 79908 153396 79960
rect 153350 79812 153378 79908
rect 153442 79880 153470 80056
rect 155926 80016 155954 80328
rect 153534 79988 155954 80016
rect 157030 79988 158392 80016
rect 153534 79960 153562 79988
rect 157030 79960 157058 79988
rect 153516 79908 153522 79960
rect 153574 79908 153580 79960
rect 153700 79908 153706 79960
rect 153758 79948 153764 79960
rect 153758 79908 153792 79948
rect 154896 79908 154902 79960
rect 154954 79908 154960 79960
rect 155448 79908 155454 79960
rect 155506 79908 155512 79960
rect 155816 79908 155822 79960
rect 155874 79908 155880 79960
rect 155908 79908 155914 79960
rect 155966 79908 155972 79960
rect 156276 79908 156282 79960
rect 156334 79908 156340 79960
rect 156368 79908 156374 79960
rect 156426 79908 156432 79960
rect 157012 79908 157018 79960
rect 157070 79908 157076 79960
rect 157564 79948 157570 79960
rect 157490 79920 157570 79948
rect 153442 79852 153608 79880
rect 153350 79784 153516 79812
rect 153212 79716 153378 79744
rect 153350 79552 153378 79716
rect 153488 79620 153516 79784
rect 153470 79568 153476 79620
rect 153528 79568 153534 79620
rect 153580 79608 153608 79852
rect 153764 79744 153792 79908
rect 153884 79840 153890 79892
rect 153942 79840 153948 79892
rect 154160 79840 154166 79892
rect 154218 79840 154224 79892
rect 154712 79840 154718 79892
rect 154770 79840 154776 79892
rect 153672 79716 153792 79744
rect 153672 79688 153700 79716
rect 153902 79688 153930 79840
rect 154178 79744 154206 79840
rect 153654 79636 153660 79688
rect 153712 79636 153718 79688
rect 153838 79636 153844 79688
rect 153896 79648 153930 79688
rect 154132 79716 154206 79744
rect 154730 79744 154758 79840
rect 154730 79716 154804 79744
rect 153896 79636 153902 79648
rect 154022 79608 154028 79620
rect 153580 79580 154028 79608
rect 154022 79568 154028 79580
rect 154080 79568 154086 79620
rect 154132 79608 154160 79716
rect 154298 79608 154304 79620
rect 154132 79580 154304 79608
rect 154298 79568 154304 79580
rect 154356 79568 154362 79620
rect 154574 79568 154580 79620
rect 154632 79608 154638 79620
rect 154776 79608 154804 79716
rect 154632 79580 154804 79608
rect 154632 79568 154638 79580
rect 152826 79500 152832 79552
rect 152884 79500 152890 79552
rect 152982 79512 153016 79552
rect 153010 79500 153016 79512
rect 153068 79500 153074 79552
rect 153286 79500 153292 79552
rect 153344 79512 153378 79552
rect 154914 79540 154942 79908
rect 155466 79552 155494 79908
rect 155834 79880 155862 79908
rect 155126 79540 155132 79552
rect 154914 79512 155132 79540
rect 153344 79500 153350 79512
rect 155126 79500 155132 79512
rect 155184 79500 155190 79552
rect 155402 79500 155408 79552
rect 155460 79512 155494 79552
rect 155788 79852 155862 79880
rect 155788 79540 155816 79852
rect 155926 79824 155954 79908
rect 155862 79772 155868 79824
rect 155920 79784 155954 79824
rect 155920 79772 155926 79784
rect 156294 79620 156322 79908
rect 156386 79676 156414 79908
rect 156460 79840 156466 79892
rect 156518 79880 156524 79892
rect 156518 79852 157104 79880
rect 156518 79840 156524 79852
rect 157076 79824 157104 79852
rect 157288 79840 157294 79892
rect 157346 79840 157352 79892
rect 157380 79840 157386 79892
rect 157438 79840 157444 79892
rect 156552 79772 156558 79824
rect 156610 79772 156616 79824
rect 156736 79772 156742 79824
rect 156794 79772 156800 79824
rect 157058 79772 157064 79824
rect 157116 79772 157122 79824
rect 156570 79744 156598 79772
rect 156570 79716 156644 79744
rect 156506 79676 156512 79688
rect 156386 79648 156512 79676
rect 156506 79636 156512 79648
rect 156564 79636 156570 79688
rect 156294 79580 156328 79620
rect 156322 79568 156328 79580
rect 156380 79568 156386 79620
rect 156414 79568 156420 79620
rect 156472 79568 156478 79620
rect 156432 79540 156460 79568
rect 155788 79512 156460 79540
rect 155460 79500 155466 79512
rect 152918 79432 152924 79484
rect 152976 79472 152982 79484
rect 152976 79444 156046 79472
rect 152976 79432 152982 79444
rect 152458 79364 152464 79416
rect 152516 79404 152522 79416
rect 155678 79404 155684 79416
rect 152516 79376 155684 79404
rect 152516 79364 152522 79376
rect 155678 79364 155684 79376
rect 155736 79364 155742 79416
rect 151964 79308 152228 79336
rect 151964 79296 151970 79308
rect 153102 79296 153108 79348
rect 153160 79336 153166 79348
rect 154942 79336 154948 79348
rect 153160 79308 154948 79336
rect 153160 79296 153166 79308
rect 154942 79296 154948 79308
rect 155000 79296 155006 79348
rect 156018 79336 156046 79444
rect 156414 79432 156420 79484
rect 156472 79472 156478 79484
rect 156616 79472 156644 79716
rect 156472 79444 156644 79472
rect 156472 79432 156478 79444
rect 156754 79404 156782 79772
rect 157306 79744 157334 79840
rect 157168 79716 157334 79744
rect 157168 79688 157196 79716
rect 157398 79688 157426 79840
rect 157150 79636 157156 79688
rect 157208 79636 157214 79688
rect 157334 79636 157340 79688
rect 157392 79648 157426 79688
rect 157392 79636 157398 79648
rect 157490 79620 157518 79920
rect 157564 79908 157570 79920
rect 157622 79908 157628 79960
rect 158208 79948 158214 79960
rect 158042 79920 158214 79948
rect 157656 79840 157662 79892
rect 157714 79840 157720 79892
rect 157748 79840 157754 79892
rect 157806 79840 157812 79892
rect 157426 79568 157432 79620
rect 157484 79580 157518 79620
rect 157484 79568 157490 79580
rect 157674 79552 157702 79840
rect 157766 79608 157794 79840
rect 158042 79744 158070 79920
rect 158208 79908 158214 79920
rect 158266 79908 158272 79960
rect 158116 79840 158122 79892
rect 158174 79840 158180 79892
rect 158134 79812 158162 79840
rect 158134 79784 158300 79812
rect 158162 79744 158168 79756
rect 158042 79716 158168 79744
rect 158162 79704 158168 79716
rect 158220 79704 158226 79756
rect 158272 79688 158300 79784
rect 158364 79688 158392 79988
rect 158484 79840 158490 79892
rect 158542 79840 158548 79892
rect 158576 79840 158582 79892
rect 158634 79840 158640 79892
rect 158502 79756 158530 79840
rect 158438 79704 158444 79756
rect 158496 79716 158530 79756
rect 158496 79704 158502 79716
rect 158594 79688 158622 79840
rect 158254 79636 158260 79688
rect 158312 79636 158318 79688
rect 158346 79636 158352 79688
rect 158404 79636 158410 79688
rect 158530 79636 158536 79688
rect 158588 79648 158622 79688
rect 158588 79636 158594 79648
rect 157766 79580 157840 79608
rect 156966 79500 156972 79552
rect 157024 79540 157030 79552
rect 157242 79540 157248 79552
rect 157024 79512 157248 79540
rect 157024 79500 157030 79512
rect 157242 79500 157248 79512
rect 157300 79500 157306 79552
rect 157674 79512 157708 79552
rect 157702 79500 157708 79512
rect 157760 79500 157766 79552
rect 157610 79432 157616 79484
rect 157668 79472 157674 79484
rect 157812 79472 157840 79580
rect 157668 79444 157840 79472
rect 157668 79432 157674 79444
rect 156966 79404 156972 79416
rect 156754 79376 156972 79404
rect 156966 79364 156972 79376
rect 157024 79364 157030 79416
rect 158686 79404 158714 80328
rect 158778 79960 158806 80600
rect 169726 80560 169754 80600
rect 174630 80588 174636 80600
rect 174688 80588 174694 80640
rect 178034 80588 178040 80640
rect 178092 80628 178098 80640
rect 580442 80628 580448 80640
rect 178092 80600 580448 80628
rect 178092 80588 178098 80600
rect 580442 80588 580448 80600
rect 580500 80588 580506 80640
rect 169726 80532 171272 80560
rect 171244 80492 171272 80532
rect 175734 80520 175740 80572
rect 175792 80560 175798 80572
rect 580350 80560 580356 80572
rect 175792 80532 580356 80560
rect 175792 80520 175798 80532
rect 580350 80520 580356 80532
rect 580408 80520 580414 80572
rect 175918 80492 175924 80504
rect 171244 80464 175924 80492
rect 175918 80452 175924 80464
rect 175976 80452 175982 80504
rect 180150 80424 180156 80436
rect 171106 80396 180156 80424
rect 164344 80124 165246 80152
rect 164344 80016 164372 80124
rect 160158 79988 160830 80016
rect 160158 79960 160186 79988
rect 158760 79908 158766 79960
rect 158818 79908 158824 79960
rect 158852 79908 158858 79960
rect 158910 79908 158916 79960
rect 159036 79908 159042 79960
rect 159094 79908 159100 79960
rect 159312 79908 159318 79960
rect 159370 79908 159376 79960
rect 159680 79908 159686 79960
rect 159738 79908 159744 79960
rect 159772 79908 159778 79960
rect 159830 79948 159836 79960
rect 159830 79908 159864 79948
rect 160048 79908 160054 79960
rect 160106 79908 160112 79960
rect 160140 79908 160146 79960
rect 160198 79908 160204 79960
rect 160232 79908 160238 79960
rect 160290 79908 160296 79960
rect 160324 79908 160330 79960
rect 160382 79908 160388 79960
rect 160416 79908 160422 79960
rect 160474 79908 160480 79960
rect 160600 79908 160606 79960
rect 160658 79908 160664 79960
rect 160692 79908 160698 79960
rect 160750 79908 160756 79960
rect 158870 79824 158898 79908
rect 158806 79772 158812 79824
rect 158864 79784 158898 79824
rect 158864 79772 158870 79784
rect 158944 79772 158950 79824
rect 159002 79772 159008 79824
rect 158962 79688 158990 79772
rect 158898 79636 158904 79688
rect 158956 79648 158990 79688
rect 158956 79636 158962 79648
rect 159054 79472 159082 79908
rect 159220 79840 159226 79892
rect 159278 79840 159284 79892
rect 159238 79620 159266 79840
rect 159330 79676 159358 79908
rect 159588 79840 159594 79892
rect 159646 79840 159652 79892
rect 159606 79812 159634 79840
rect 159560 79784 159634 79812
rect 159330 79648 159496 79676
rect 159238 79580 159272 79620
rect 159266 79568 159272 79580
rect 159324 79568 159330 79620
rect 159174 79500 159180 79552
rect 159232 79540 159238 79552
rect 159468 79540 159496 79648
rect 159560 79620 159588 79784
rect 159698 79756 159726 79908
rect 159634 79704 159640 79756
rect 159692 79716 159726 79756
rect 159692 79704 159698 79716
rect 159542 79568 159548 79620
rect 159600 79568 159606 79620
rect 159836 79552 159864 79908
rect 160066 79880 160094 79908
rect 160250 79880 160278 79908
rect 159928 79852 160094 79880
rect 160204 79852 160278 79880
rect 159232 79512 159496 79540
rect 159232 79500 159238 79512
rect 159818 79500 159824 79552
rect 159876 79500 159882 79552
rect 159928 79484 159956 79852
rect 160204 79824 160232 79852
rect 160342 79824 160370 79908
rect 160186 79772 160192 79824
rect 160244 79772 160250 79824
rect 160278 79772 160284 79824
rect 160336 79784 160370 79824
rect 160336 79772 160342 79784
rect 160434 79688 160462 79908
rect 160618 79824 160646 79908
rect 160600 79772 160606 79824
rect 160658 79772 160664 79824
rect 160710 79744 160738 79908
rect 160572 79716 160738 79744
rect 160434 79648 160468 79688
rect 160462 79636 160468 79648
rect 160520 79636 160526 79688
rect 160572 79620 160600 79716
rect 160554 79568 160560 79620
rect 160612 79568 160618 79620
rect 160802 79608 160830 79988
rect 162550 79988 164096 80016
rect 162550 79960 162578 79988
rect 161152 79908 161158 79960
rect 161210 79948 161216 79960
rect 161210 79920 162486 79948
rect 161210 79908 161216 79920
rect 161060 79840 161066 79892
rect 161118 79880 161124 79892
rect 161336 79880 161342 79892
rect 161118 79840 161152 79880
rect 160968 79772 160974 79824
rect 161026 79812 161032 79824
rect 161026 79772 161060 79812
rect 161032 79688 161060 79772
rect 161124 79756 161152 79840
rect 161216 79852 161342 79880
rect 161216 79824 161244 79852
rect 161336 79840 161342 79852
rect 161394 79840 161400 79892
rect 161612 79840 161618 79892
rect 161670 79840 161676 79892
rect 161888 79840 161894 79892
rect 161946 79840 161952 79892
rect 162164 79840 162170 79892
rect 162222 79840 162228 79892
rect 161198 79772 161204 79824
rect 161256 79772 161262 79824
rect 161106 79704 161112 79756
rect 161164 79704 161170 79756
rect 161014 79636 161020 79688
rect 161072 79636 161078 79688
rect 161630 79676 161658 79840
rect 161906 79744 161934 79840
rect 161906 79716 162072 79744
rect 162044 79688 162072 79716
rect 161934 79676 161940 79688
rect 161630 79648 161940 79676
rect 161934 79636 161940 79648
rect 161992 79636 161998 79688
rect 162026 79636 162032 79688
rect 162084 79636 162090 79688
rect 160922 79608 160928 79620
rect 160802 79580 160928 79608
rect 160922 79568 160928 79580
rect 160980 79568 160986 79620
rect 162182 79608 162210 79840
rect 162256 79772 162262 79824
rect 162314 79772 162320 79824
rect 161400 79580 162210 79608
rect 161400 79552 161428 79580
rect 161382 79500 161388 79552
rect 161440 79500 161446 79552
rect 159726 79472 159732 79484
rect 159054 79444 159732 79472
rect 159726 79432 159732 79444
rect 159784 79432 159790 79484
rect 159910 79432 159916 79484
rect 159968 79432 159974 79484
rect 162118 79404 162124 79416
rect 158686 79376 162124 79404
rect 162118 79364 162124 79376
rect 162176 79364 162182 79416
rect 162274 79404 162302 79772
rect 162458 79744 162486 79920
rect 162532 79908 162538 79960
rect 162590 79908 162596 79960
rect 163268 79908 163274 79960
rect 163326 79908 163332 79960
rect 163912 79908 163918 79960
rect 163970 79948 163976 79960
rect 163970 79908 164004 79948
rect 162716 79840 162722 79892
rect 162774 79840 162780 79892
rect 163084 79880 163090 79892
rect 163056 79840 163090 79880
rect 163142 79840 163148 79892
rect 163176 79840 163182 79892
rect 163234 79840 163240 79892
rect 162578 79772 162584 79824
rect 162636 79812 162642 79824
rect 162734 79812 162762 79840
rect 162636 79784 162762 79812
rect 162636 79772 162642 79784
rect 163056 79756 163084 79840
rect 163194 79756 163222 79840
rect 162670 79744 162676 79756
rect 162458 79716 162676 79744
rect 162670 79704 162676 79716
rect 162728 79704 162734 79756
rect 163038 79704 163044 79756
rect 163096 79704 163102 79756
rect 163130 79704 163136 79756
rect 163188 79716 163222 79756
rect 163188 79704 163194 79716
rect 162946 79636 162952 79688
rect 163004 79676 163010 79688
rect 163286 79676 163314 79908
rect 163728 79840 163734 79892
rect 163786 79840 163792 79892
rect 163820 79840 163826 79892
rect 163878 79880 163884 79892
rect 163878 79840 163912 79880
rect 163544 79772 163550 79824
rect 163602 79772 163608 79824
rect 163004 79648 163314 79676
rect 163004 79636 163010 79648
rect 163562 79552 163590 79772
rect 163746 79676 163774 79840
rect 163700 79648 163774 79676
rect 163700 79552 163728 79648
rect 163884 79620 163912 79840
rect 163866 79568 163872 79620
rect 163924 79568 163930 79620
rect 163498 79500 163504 79552
rect 163556 79512 163590 79552
rect 163556 79500 163562 79512
rect 163682 79500 163688 79552
rect 163740 79500 163746 79552
rect 162854 79432 162860 79484
rect 162912 79472 162918 79484
rect 163976 79472 164004 79908
rect 164068 79620 164096 79988
rect 164160 79988 164372 80016
rect 164160 79688 164188 79988
rect 165218 79960 165246 80124
rect 165954 79988 166856 80016
rect 165954 79960 165982 79988
rect 164556 79908 164562 79960
rect 164614 79948 164620 79960
rect 164614 79920 165154 79948
rect 164614 79908 164620 79920
rect 165016 79840 165022 79892
rect 165074 79840 165080 79892
rect 164832 79772 164838 79824
rect 164890 79772 164896 79824
rect 164142 79636 164148 79688
rect 164200 79636 164206 79688
rect 164850 79620 164878 79772
rect 165034 79744 165062 79840
rect 165126 79812 165154 79920
rect 165200 79908 165206 79960
rect 165258 79908 165264 79960
rect 165936 79908 165942 79960
rect 165994 79908 166000 79960
rect 166396 79908 166402 79960
rect 166454 79908 166460 79960
rect 165660 79840 165666 79892
rect 165718 79840 165724 79892
rect 166120 79840 166126 79892
rect 166178 79840 166184 79892
rect 165246 79812 165252 79824
rect 165126 79784 165252 79812
rect 165246 79772 165252 79784
rect 165304 79772 165310 79824
rect 165034 79716 165568 79744
rect 165540 79620 165568 79716
rect 165678 79676 165706 79840
rect 165632 79648 165706 79676
rect 164050 79568 164056 79620
rect 164108 79568 164114 79620
rect 164786 79568 164792 79620
rect 164844 79580 164878 79620
rect 164844 79568 164850 79580
rect 165522 79568 165528 79620
rect 165580 79568 165586 79620
rect 165632 79540 165660 79648
rect 165706 79568 165712 79620
rect 165764 79608 165770 79620
rect 166138 79608 166166 79840
rect 165764 79580 166166 79608
rect 165764 79568 165770 79580
rect 166258 79568 166264 79620
rect 166316 79608 166322 79620
rect 166414 79608 166442 79908
rect 166828 79688 166856 79988
rect 167518 79988 168190 80016
rect 167518 79960 167546 79988
rect 167500 79908 167506 79960
rect 167558 79908 167564 79960
rect 167776 79908 167782 79960
rect 167834 79908 167840 79960
rect 167040 79840 167046 79892
rect 167098 79840 167104 79892
rect 166810 79636 166816 79688
rect 166868 79636 166874 79688
rect 166316 79580 166442 79608
rect 166316 79568 166322 79580
rect 166626 79540 166632 79552
rect 165632 79512 166632 79540
rect 166626 79500 166632 79512
rect 166684 79500 166690 79552
rect 167058 79540 167086 79840
rect 167362 79568 167368 79620
rect 167420 79608 167426 79620
rect 167794 79608 167822 79908
rect 168162 79880 168190 79988
rect 168806 79988 169478 80016
rect 168328 79908 168334 79960
rect 168386 79948 168392 79960
rect 168386 79920 168742 79948
rect 168386 79908 168392 79920
rect 168162 79852 168328 79880
rect 168300 79824 168328 79852
rect 168420 79840 168426 79892
rect 168478 79840 168484 79892
rect 168282 79772 168288 79824
rect 168340 79772 168346 79824
rect 168438 79756 168466 79840
rect 168374 79704 168380 79756
rect 168432 79716 168466 79756
rect 168432 79704 168438 79716
rect 167420 79580 167822 79608
rect 168714 79608 168742 79920
rect 168806 79676 168834 79988
rect 169450 79960 169478 79988
rect 170324 79988 170858 80016
rect 168880 79908 168886 79960
rect 168938 79908 168944 79960
rect 169064 79908 169070 79960
rect 169122 79908 169128 79960
rect 169432 79908 169438 79960
rect 169490 79908 169496 79960
rect 168898 79744 168926 79908
rect 169082 79812 169110 79908
rect 169248 79840 169254 79892
rect 169306 79840 169312 79892
rect 169082 79784 169156 79812
rect 169018 79744 169024 79756
rect 168898 79716 169024 79744
rect 169018 79704 169024 79716
rect 169076 79704 169082 79756
rect 168926 79676 168932 79688
rect 168806 79648 168932 79676
rect 168926 79636 168932 79648
rect 168984 79636 168990 79688
rect 168834 79608 168840 79620
rect 168714 79580 168840 79608
rect 167420 79568 167426 79580
rect 168834 79568 168840 79580
rect 168892 79568 168898 79620
rect 167058 79512 168420 79540
rect 162912 79444 164004 79472
rect 162912 79432 162918 79444
rect 164878 79432 164884 79484
rect 164936 79472 164942 79484
rect 164936 79444 167592 79472
rect 164936 79432 164942 79444
rect 163958 79404 163964 79416
rect 162274 79376 163964 79404
rect 163958 79364 163964 79376
rect 164016 79364 164022 79416
rect 164234 79364 164240 79416
rect 164292 79404 164298 79416
rect 166902 79404 166908 79416
rect 164292 79376 166908 79404
rect 164292 79364 164298 79376
rect 166902 79364 166908 79376
rect 166960 79364 166966 79416
rect 164878 79336 164884 79348
rect 156018 79308 164884 79336
rect 164878 79296 164884 79308
rect 164936 79296 164942 79348
rect 165522 79296 165528 79348
rect 165580 79336 165586 79348
rect 167454 79336 167460 79348
rect 165580 79308 167460 79336
rect 165580 79296 165586 79308
rect 167454 79296 167460 79308
rect 167512 79296 167518 79348
rect 167564 79336 167592 79444
rect 168392 79404 168420 79512
rect 168650 79404 168656 79416
rect 168392 79376 168656 79404
rect 168650 79364 168656 79376
rect 168708 79364 168714 79416
rect 169128 79404 169156 79784
rect 169266 79688 169294 79840
rect 169800 79772 169806 79824
rect 169858 79772 169864 79824
rect 169818 79688 169846 79772
rect 169202 79636 169208 79688
rect 169260 79648 169294 79688
rect 169260 79636 169266 79648
rect 169754 79636 169760 79688
rect 169812 79648 169846 79688
rect 169812 79636 169818 79648
rect 169984 79636 169990 79688
rect 170042 79636 170048 79688
rect 170002 79552 170030 79636
rect 170002 79512 170036 79552
rect 170030 79500 170036 79512
rect 170088 79500 170094 79552
rect 169726 79444 170260 79472
rect 169294 79404 169300 79416
rect 169128 79376 169300 79404
rect 169294 79364 169300 79376
rect 169352 79364 169358 79416
rect 169726 79336 169754 79444
rect 167564 79308 169754 79336
rect 170232 79336 170260 79444
rect 170324 79416 170352 79988
rect 170628 79908 170634 79960
rect 170686 79908 170692 79960
rect 170646 79880 170674 79908
rect 170600 79852 170674 79880
rect 170306 79364 170312 79416
rect 170364 79364 170370 79416
rect 170600 79404 170628 79852
rect 170720 79840 170726 79892
rect 170778 79840 170784 79892
rect 170738 79620 170766 79840
rect 170830 79744 170858 79988
rect 171106 79960 171134 80396
rect 180150 80384 180156 80396
rect 180208 80384 180214 80436
rect 171382 80328 178034 80356
rect 171382 80084 171410 80328
rect 178006 80288 178034 80328
rect 231854 80288 231860 80300
rect 178006 80260 231860 80288
rect 231854 80248 231860 80260
rect 231912 80248 231918 80300
rect 174446 80180 174452 80232
rect 174504 80220 174510 80232
rect 249794 80220 249800 80232
rect 174504 80192 249800 80220
rect 174504 80180 174510 80192
rect 249794 80180 249800 80192
rect 249852 80180 249858 80232
rect 175734 80152 175740 80164
rect 171244 80056 171410 80084
rect 172118 80124 175740 80152
rect 171088 79908 171094 79960
rect 171146 79908 171152 79960
rect 171244 79744 171272 80056
rect 172118 79960 172146 80124
rect 175734 80112 175740 80124
rect 175792 80112 175798 80164
rect 175826 80112 175832 80164
rect 175884 80152 175890 80164
rect 284294 80152 284300 80164
rect 175884 80124 284300 80152
rect 175884 80112 175890 80124
rect 284294 80112 284300 80124
rect 284352 80112 284358 80164
rect 175090 80084 175096 80096
rect 173866 80056 175096 80084
rect 173866 80016 173894 80056
rect 175090 80044 175096 80056
rect 175148 80044 175154 80096
rect 175918 80044 175924 80096
rect 175976 80084 175982 80096
rect 426434 80084 426440 80096
rect 175976 80056 426440 80084
rect 175976 80044 175982 80056
rect 426434 80044 426440 80056
rect 426492 80044 426498 80096
rect 172210 79988 173894 80016
rect 172210 79960 172238 79988
rect 171548 79908 171554 79960
rect 171606 79908 171612 79960
rect 171824 79908 171830 79960
rect 171882 79908 171888 79960
rect 171916 79908 171922 79960
rect 171974 79908 171980 79960
rect 172100 79908 172106 79960
rect 172158 79908 172164 79960
rect 172192 79908 172198 79960
rect 172250 79908 172256 79960
rect 172560 79908 172566 79960
rect 172618 79948 172624 79960
rect 172618 79920 173618 79948
rect 172618 79908 172624 79920
rect 170830 79716 171272 79744
rect 171566 79756 171594 79908
rect 171640 79840 171646 79892
rect 171698 79840 171704 79892
rect 171658 79812 171686 79840
rect 171658 79784 171732 79812
rect 171566 79716 171600 79756
rect 171594 79704 171600 79716
rect 171652 79704 171658 79756
rect 170858 79636 170864 79688
rect 170916 79676 170922 79688
rect 170916 79648 171134 79676
rect 170916 79636 170922 79648
rect 170738 79580 170772 79620
rect 170766 79568 170772 79580
rect 170824 79568 170830 79620
rect 171106 79472 171134 79648
rect 171704 79540 171732 79784
rect 171842 79676 171870 79908
rect 171934 79812 171962 79908
rect 172928 79880 172934 79892
rect 172486 79852 172934 79880
rect 172054 79812 172060 79824
rect 171934 79784 172060 79812
rect 172054 79772 172060 79784
rect 172112 79772 172118 79824
rect 172146 79772 172152 79824
rect 172204 79812 172210 79824
rect 172486 79812 172514 79852
rect 172928 79840 172934 79852
rect 172986 79840 172992 79892
rect 173296 79840 173302 79892
rect 173354 79840 173360 79892
rect 173314 79812 173342 79840
rect 172204 79784 172514 79812
rect 173084 79784 173342 79812
rect 173590 79824 173618 79920
rect 173664 79908 173670 79960
rect 173722 79948 173728 79960
rect 173722 79920 173894 79948
rect 173722 79908 173728 79920
rect 173590 79784 173624 79824
rect 172204 79772 172210 79784
rect 173084 79688 173112 79784
rect 173618 79772 173624 79784
rect 173676 79772 173682 79824
rect 173250 79704 173256 79756
rect 173308 79744 173314 79756
rect 173866 79744 173894 79920
rect 173940 79840 173946 79892
rect 173998 79880 174004 79892
rect 173998 79852 174262 79880
rect 173998 79840 174004 79852
rect 174124 79772 174130 79824
rect 174182 79772 174188 79824
rect 173308 79716 173894 79744
rect 173308 79704 173314 79716
rect 173986 79704 173992 79756
rect 174044 79744 174050 79756
rect 174142 79744 174170 79772
rect 174044 79716 174170 79744
rect 174044 79704 174050 79716
rect 171962 79676 171968 79688
rect 171842 79648 171968 79676
rect 171962 79636 171968 79648
rect 172020 79636 172026 79688
rect 173066 79636 173072 79688
rect 173124 79636 173130 79688
rect 174078 79636 174084 79688
rect 174136 79676 174142 79688
rect 174234 79676 174262 79852
rect 174136 79648 174262 79676
rect 174136 79636 174142 79648
rect 174538 79636 174544 79688
rect 174596 79676 174602 79688
rect 373994 79676 374000 79688
rect 174596 79648 374000 79676
rect 174596 79636 174602 79648
rect 373994 79636 374000 79648
rect 374052 79636 374058 79688
rect 172606 79568 172612 79620
rect 172664 79608 172670 79620
rect 179506 79608 179512 79620
rect 172664 79580 179512 79608
rect 172664 79568 172670 79580
rect 179506 79568 179512 79580
rect 179564 79568 179570 79620
rect 171704 79512 175044 79540
rect 171686 79472 171692 79484
rect 171106 79444 171692 79472
rect 171686 79432 171692 79444
rect 171744 79432 171750 79484
rect 171778 79432 171784 79484
rect 171836 79472 171842 79484
rect 173158 79472 173164 79484
rect 171836 79444 173164 79472
rect 171836 79432 171842 79444
rect 173158 79432 173164 79444
rect 173216 79432 173222 79484
rect 173710 79432 173716 79484
rect 173768 79472 173774 79484
rect 174630 79472 174636 79484
rect 173768 79444 174636 79472
rect 173768 79432 173774 79444
rect 174630 79432 174636 79444
rect 174688 79432 174694 79484
rect 171502 79404 171508 79416
rect 170600 79376 171508 79404
rect 171502 79364 171508 79376
rect 171560 79364 171566 79416
rect 173342 79404 173348 79416
rect 171612 79376 173348 79404
rect 171612 79336 171640 79376
rect 173342 79364 173348 79376
rect 173400 79364 173406 79416
rect 175016 79404 175044 79512
rect 177390 79500 177396 79552
rect 177448 79540 177454 79552
rect 331214 79540 331220 79552
rect 177448 79512 331220 79540
rect 177448 79500 177454 79512
rect 331214 79500 331220 79512
rect 331272 79500 331278 79552
rect 175090 79432 175096 79484
rect 175148 79472 175154 79484
rect 580258 79472 580264 79484
rect 175148 79444 580264 79472
rect 175148 79432 175154 79444
rect 580258 79432 580264 79444
rect 580316 79432 580322 79484
rect 580626 79404 580632 79416
rect 175016 79376 580632 79404
rect 580626 79364 580632 79376
rect 580684 79364 580690 79416
rect 170232 79308 171640 79336
rect 171686 79296 171692 79348
rect 171744 79336 171750 79348
rect 173802 79336 173808 79348
rect 171744 79308 173808 79336
rect 171744 79296 171750 79308
rect 173802 79296 173808 79308
rect 173860 79296 173866 79348
rect 580534 79336 580540 79348
rect 180766 79308 580540 79336
rect 165154 79268 165160 79280
rect 154546 79240 165160 79268
rect 154546 79200 154574 79240
rect 165154 79228 165160 79240
rect 165212 79228 165218 79280
rect 165430 79228 165436 79280
rect 165488 79268 165494 79280
rect 165488 79240 170260 79268
rect 165488 79228 165494 79240
rect 150406 79172 154574 79200
rect 155678 79160 155684 79212
rect 155736 79200 155742 79212
rect 155736 79172 164924 79200
rect 155736 79160 155742 79172
rect 152458 79132 152464 79144
rect 118666 79104 140774 79132
rect 145576 79104 152464 79132
rect 128078 79024 128084 79076
rect 128136 79064 128142 79076
rect 128630 79064 128636 79076
rect 128136 79036 128636 79064
rect 128136 79024 128142 79036
rect 128630 79024 128636 79036
rect 128688 79024 128694 79076
rect 129090 79024 129096 79076
rect 129148 79064 129154 79076
rect 133874 79064 133880 79076
rect 129148 79036 133880 79064
rect 129148 79024 129154 79036
rect 133874 79024 133880 79036
rect 133932 79024 133938 79076
rect 130378 78956 130384 79008
rect 130436 78996 130442 79008
rect 130562 78996 130568 79008
rect 130436 78968 130568 78996
rect 130436 78956 130442 78968
rect 130562 78956 130568 78968
rect 130620 78956 130626 79008
rect 140746 78996 140774 79104
rect 152458 79092 152464 79104
rect 152516 79092 152522 79144
rect 158346 79092 158352 79144
rect 158404 79132 158410 79144
rect 158990 79132 158996 79144
rect 158404 79104 158996 79132
rect 158404 79092 158410 79104
rect 158990 79092 158996 79104
rect 159048 79092 159054 79144
rect 159726 79092 159732 79144
rect 159784 79132 159790 79144
rect 164896 79132 164924 79172
rect 165798 79160 165804 79212
rect 165856 79200 165862 79212
rect 168006 79200 168012 79212
rect 165856 79172 168012 79200
rect 165856 79160 165862 79172
rect 168006 79160 168012 79172
rect 168064 79160 168070 79212
rect 168834 79160 168840 79212
rect 168892 79200 168898 79212
rect 169570 79200 169576 79212
rect 168892 79172 169576 79200
rect 168892 79160 168898 79172
rect 169570 79160 169576 79172
rect 169628 79160 169634 79212
rect 169754 79160 169760 79212
rect 169812 79200 169818 79212
rect 170122 79200 170128 79212
rect 169812 79172 170128 79200
rect 169812 79160 169818 79172
rect 170122 79160 170128 79172
rect 170180 79160 170186 79212
rect 170232 79200 170260 79240
rect 171594 79228 171600 79280
rect 171652 79268 171658 79280
rect 180766 79268 180794 79308
rect 580534 79296 580540 79308
rect 580592 79296 580598 79348
rect 171652 79240 180794 79268
rect 171652 79228 171658 79240
rect 171686 79200 171692 79212
rect 170232 79172 171692 79200
rect 171686 79160 171692 79172
rect 171744 79160 171750 79212
rect 171870 79160 171876 79212
rect 171928 79200 171934 79212
rect 175826 79200 175832 79212
rect 171928 79172 175832 79200
rect 171928 79160 171934 79172
rect 175826 79160 175832 79172
rect 175884 79160 175890 79212
rect 170950 79132 170956 79144
rect 159784 79104 164832 79132
rect 164896 79104 170956 79132
rect 159784 79092 159790 79104
rect 154022 79024 154028 79076
rect 154080 79064 154086 79076
rect 163130 79064 163136 79076
rect 154080 79036 163136 79064
rect 154080 79024 154086 79036
rect 163130 79024 163136 79036
rect 163188 79024 163194 79076
rect 164804 79064 164832 79104
rect 170950 79092 170956 79104
rect 171008 79092 171014 79144
rect 171318 79092 171324 79144
rect 171376 79132 171382 79144
rect 182910 79132 182916 79144
rect 171376 79104 182916 79132
rect 171376 79092 171382 79104
rect 182910 79092 182916 79104
rect 182968 79092 182974 79144
rect 165798 79064 165804 79076
rect 164804 79036 165804 79064
rect 165798 79024 165804 79036
rect 165856 79024 165862 79076
rect 166074 79024 166080 79076
rect 166132 79064 166138 79076
rect 200114 79064 200120 79076
rect 166132 79036 200120 79064
rect 166132 79024 166138 79036
rect 200114 79024 200120 79036
rect 200172 79024 200178 79076
rect 153102 78996 153108 79008
rect 140746 78968 153108 78996
rect 153102 78956 153108 78968
rect 153160 78956 153166 79008
rect 159174 78956 159180 79008
rect 159232 78996 159238 79008
rect 252554 78996 252560 79008
rect 159232 78968 252560 78996
rect 159232 78956 159238 78968
rect 252554 78956 252560 78968
rect 252612 78956 252618 79008
rect 118666 78900 140774 78928
rect 44818 78752 44824 78804
rect 44876 78792 44882 78804
rect 118666 78792 118694 78900
rect 140746 78860 140774 78900
rect 145466 78888 145472 78940
rect 145524 78928 145530 78940
rect 152918 78928 152924 78940
rect 145524 78900 152924 78928
rect 145524 78888 145530 78900
rect 152918 78888 152924 78900
rect 152976 78888 152982 78940
rect 154942 78888 154948 78940
rect 155000 78928 155006 78940
rect 165430 78928 165436 78940
rect 155000 78900 165436 78928
rect 155000 78888 155006 78900
rect 165430 78888 165436 78900
rect 165488 78888 165494 78940
rect 165522 78888 165528 78940
rect 165580 78928 165586 78940
rect 213914 78928 213920 78940
rect 165580 78900 213920 78928
rect 165580 78888 165586 78900
rect 213914 78888 213920 78900
rect 213972 78888 213978 78940
rect 306374 78860 306380 78872
rect 140746 78832 159404 78860
rect 44876 78764 118694 78792
rect 44876 78752 44882 78764
rect 154666 78752 154672 78804
rect 154724 78792 154730 78804
rect 155034 78792 155040 78804
rect 154724 78764 155040 78792
rect 154724 78752 154730 78764
rect 155034 78752 155040 78764
rect 155092 78752 155098 78804
rect 157978 78752 157984 78804
rect 158036 78792 158042 78804
rect 158254 78792 158260 78804
rect 158036 78764 158260 78792
rect 158036 78752 158042 78764
rect 158254 78752 158260 78764
rect 158312 78752 158318 78804
rect 125962 78684 125968 78736
rect 126020 78724 126026 78736
rect 126330 78724 126336 78736
rect 126020 78696 126336 78724
rect 126020 78684 126026 78696
rect 126330 78684 126336 78696
rect 126388 78684 126394 78736
rect 155954 78684 155960 78736
rect 156012 78724 156018 78736
rect 156230 78724 156236 78736
rect 156012 78696 156236 78724
rect 156012 78684 156018 78696
rect 156230 78684 156236 78696
rect 156288 78684 156294 78736
rect 159376 78724 159404 78832
rect 159928 78832 306380 78860
rect 159726 78752 159732 78804
rect 159784 78792 159790 78804
rect 159928 78792 159956 78832
rect 306374 78820 306380 78832
rect 306432 78820 306438 78872
rect 159784 78764 159956 78792
rect 159784 78752 159790 78764
rect 164234 78752 164240 78804
rect 164292 78792 164298 78804
rect 164694 78792 164700 78804
rect 164292 78764 164700 78792
rect 164292 78752 164298 78764
rect 164694 78752 164700 78764
rect 164752 78752 164758 78804
rect 164878 78752 164884 78804
rect 164936 78792 164942 78804
rect 173894 78792 173900 78804
rect 164936 78764 173900 78792
rect 164936 78752 164942 78764
rect 173894 78752 173900 78764
rect 173952 78752 173958 78804
rect 201494 78792 201500 78804
rect 180766 78764 201500 78792
rect 159376 78696 164924 78724
rect 124030 78616 124036 78668
rect 124088 78656 124094 78668
rect 128078 78656 128084 78668
rect 124088 78628 128084 78656
rect 124088 78616 124094 78628
rect 128078 78616 128084 78628
rect 128136 78616 128142 78668
rect 135346 78616 135352 78668
rect 135404 78656 135410 78668
rect 135806 78656 135812 78668
rect 135404 78628 135812 78656
rect 135404 78616 135410 78628
rect 135806 78616 135812 78628
rect 135864 78616 135870 78668
rect 147582 78616 147588 78668
rect 147640 78656 147646 78668
rect 164896 78656 164924 78696
rect 165154 78684 165160 78736
rect 165212 78724 165218 78736
rect 170950 78724 170956 78736
rect 165212 78696 170956 78724
rect 165212 78684 165218 78696
rect 170950 78684 170956 78696
rect 171008 78684 171014 78736
rect 171226 78684 171232 78736
rect 171284 78724 171290 78736
rect 172422 78724 172428 78736
rect 171284 78696 172428 78724
rect 171284 78684 171290 78696
rect 172422 78684 172428 78696
rect 172480 78684 172486 78736
rect 172606 78684 172612 78736
rect 172664 78724 172670 78736
rect 180766 78724 180794 78764
rect 201494 78752 201500 78764
rect 201552 78752 201558 78804
rect 172664 78696 180794 78724
rect 172664 78684 172670 78696
rect 147640 78628 164832 78656
rect 164896 78628 171824 78656
rect 147640 78616 147646 78628
rect 93118 78548 93124 78600
rect 93176 78588 93182 78600
rect 127986 78588 127992 78600
rect 93176 78560 127992 78588
rect 93176 78548 93182 78560
rect 127986 78548 127992 78560
rect 128044 78548 128050 78600
rect 155862 78548 155868 78600
rect 155920 78588 155926 78600
rect 157978 78588 157984 78600
rect 155920 78560 157984 78588
rect 155920 78548 155926 78560
rect 157978 78548 157984 78560
rect 158036 78548 158042 78600
rect 164694 78588 164700 78600
rect 159376 78560 164700 78588
rect 126146 78480 126152 78532
rect 126204 78520 126210 78532
rect 126330 78520 126336 78532
rect 126204 78492 126336 78520
rect 126204 78480 126210 78492
rect 126330 78480 126336 78492
rect 126388 78480 126394 78532
rect 130010 78480 130016 78532
rect 130068 78520 130074 78532
rect 130746 78520 130752 78532
rect 130068 78492 130752 78520
rect 130068 78480 130074 78492
rect 130746 78480 130752 78492
rect 130804 78480 130810 78532
rect 141234 78480 141240 78532
rect 141292 78520 141298 78532
rect 159376 78520 159404 78560
rect 164694 78548 164700 78560
rect 164752 78548 164758 78600
rect 141292 78492 159404 78520
rect 164804 78520 164832 78628
rect 166902 78548 166908 78600
rect 166960 78588 166966 78600
rect 171686 78588 171692 78600
rect 166960 78560 171692 78588
rect 166960 78548 166966 78560
rect 171686 78548 171692 78560
rect 171744 78548 171750 78600
rect 171796 78588 171824 78628
rect 171962 78616 171968 78668
rect 172020 78656 172026 78668
rect 182266 78656 182272 78668
rect 172020 78628 182272 78656
rect 172020 78616 172026 78628
rect 182266 78616 182272 78628
rect 182324 78616 182330 78668
rect 173526 78588 173532 78600
rect 171796 78560 173532 78588
rect 173526 78548 173532 78560
rect 173584 78548 173590 78600
rect 170858 78520 170864 78532
rect 164804 78492 170864 78520
rect 141292 78480 141298 78492
rect 170858 78480 170864 78492
rect 170916 78480 170922 78532
rect 170950 78480 170956 78532
rect 171008 78520 171014 78532
rect 171134 78520 171140 78532
rect 171008 78492 171140 78520
rect 171008 78480 171014 78492
rect 171134 78480 171140 78492
rect 171192 78480 171198 78532
rect 172882 78480 172888 78532
rect 172940 78520 172946 78532
rect 180794 78520 180800 78532
rect 172940 78492 180800 78520
rect 172940 78480 172946 78492
rect 180794 78480 180800 78492
rect 180852 78480 180858 78532
rect 123662 78412 123668 78464
rect 123720 78452 123726 78464
rect 134886 78452 134892 78464
rect 123720 78424 134892 78452
rect 123720 78412 123726 78424
rect 134886 78412 134892 78424
rect 134944 78412 134950 78464
rect 153194 78412 153200 78464
rect 153252 78452 153258 78464
rect 156230 78452 156236 78464
rect 153252 78424 156236 78452
rect 153252 78412 153258 78424
rect 156230 78412 156236 78424
rect 156288 78412 156294 78464
rect 157702 78412 157708 78464
rect 157760 78452 157766 78464
rect 158070 78452 158076 78464
rect 157760 78424 158076 78452
rect 157760 78412 157766 78424
rect 158070 78412 158076 78424
rect 158128 78412 158134 78464
rect 161658 78412 161664 78464
rect 161716 78452 161722 78464
rect 161716 78424 167040 78452
rect 161716 78412 161722 78424
rect 127066 78344 127072 78396
rect 127124 78384 127130 78396
rect 135254 78384 135260 78396
rect 127124 78356 135260 78384
rect 127124 78344 127130 78356
rect 135254 78344 135260 78356
rect 135312 78344 135318 78396
rect 149514 78344 149520 78396
rect 149572 78384 149578 78396
rect 159726 78384 159732 78396
rect 149572 78356 159732 78384
rect 149572 78344 149578 78356
rect 159726 78344 159732 78356
rect 159784 78344 159790 78396
rect 162118 78344 162124 78396
rect 162176 78384 162182 78396
rect 165154 78384 165160 78396
rect 162176 78356 165160 78384
rect 162176 78344 162182 78356
rect 165154 78344 165160 78356
rect 165212 78344 165218 78396
rect 167012 78384 167040 78424
rect 167638 78412 167644 78464
rect 167696 78452 167702 78464
rect 242158 78452 242164 78464
rect 167696 78424 242164 78452
rect 167696 78412 167702 78424
rect 242158 78412 242164 78424
rect 242216 78412 242222 78464
rect 315298 78384 315304 78396
rect 167012 78356 315304 78384
rect 315298 78344 315304 78356
rect 315356 78344 315362 78396
rect 125870 78316 125876 78328
rect 118666 78288 125876 78316
rect 113818 78208 113824 78260
rect 113876 78248 113882 78260
rect 118666 78248 118694 78288
rect 125870 78276 125876 78288
rect 125928 78276 125934 78328
rect 142246 78276 142252 78328
rect 142304 78316 142310 78328
rect 165522 78316 165528 78328
rect 142304 78288 165528 78316
rect 142304 78276 142310 78288
rect 165522 78276 165528 78288
rect 165580 78276 165586 78328
rect 165798 78276 165804 78328
rect 165856 78316 165862 78328
rect 430574 78316 430580 78328
rect 165856 78288 430580 78316
rect 165856 78276 165862 78288
rect 430574 78276 430580 78288
rect 430632 78276 430638 78328
rect 129642 78248 129648 78260
rect 113876 78220 118694 78248
rect 123496 78220 129648 78248
rect 113876 78208 113882 78220
rect 110414 78140 110420 78192
rect 110472 78180 110478 78192
rect 123496 78180 123524 78220
rect 129642 78208 129648 78220
rect 129700 78208 129706 78260
rect 144914 78248 144920 78260
rect 144840 78220 144920 78248
rect 110472 78152 123524 78180
rect 110472 78140 110478 78152
rect 132494 78112 132500 78124
rect 124186 78084 132500 78112
rect 89714 78004 89720 78056
rect 89772 78044 89778 78056
rect 124186 78044 124214 78084
rect 132494 78072 132500 78084
rect 132552 78072 132558 78124
rect 89772 78016 124214 78044
rect 144840 78044 144868 78220
rect 144914 78208 144920 78220
rect 144972 78208 144978 78260
rect 154758 78208 154764 78260
rect 154816 78248 154822 78260
rect 161290 78248 161296 78260
rect 154816 78220 161296 78248
rect 154816 78208 154822 78220
rect 161290 78208 161296 78220
rect 161348 78208 161354 78260
rect 162762 78208 162768 78260
rect 162820 78248 162826 78260
rect 436738 78248 436744 78260
rect 162820 78220 436744 78248
rect 162820 78208 162826 78220
rect 436738 78208 436744 78220
rect 436796 78208 436802 78260
rect 145282 78140 145288 78192
rect 145340 78180 145346 78192
rect 145340 78152 150434 78180
rect 145340 78140 145346 78152
rect 150406 78112 150434 78152
rect 150802 78140 150808 78192
rect 150860 78180 150866 78192
rect 151170 78180 151176 78192
rect 150860 78152 151176 78180
rect 150860 78140 150866 78152
rect 151170 78140 151176 78152
rect 151228 78140 151234 78192
rect 155310 78140 155316 78192
rect 155368 78180 155374 78192
rect 159726 78180 159732 78192
rect 155368 78152 159732 78180
rect 155368 78140 155374 78152
rect 159726 78140 159732 78152
rect 159784 78140 159790 78192
rect 164694 78140 164700 78192
rect 164752 78180 164758 78192
rect 164752 78152 165108 78180
rect 164752 78140 164758 78152
rect 159174 78112 159180 78124
rect 150406 78084 159180 78112
rect 159174 78072 159180 78084
rect 159232 78072 159238 78124
rect 164418 78072 164424 78124
rect 164476 78112 164482 78124
rect 164970 78112 164976 78124
rect 164476 78084 164976 78112
rect 164476 78072 164482 78084
rect 164970 78072 164976 78084
rect 165028 78072 165034 78124
rect 165080 78112 165108 78152
rect 165430 78140 165436 78192
rect 165488 78180 165494 78192
rect 480254 78180 480260 78192
rect 165488 78152 480260 78180
rect 165488 78140 165494 78152
rect 480254 78140 480260 78152
rect 480312 78140 480318 78192
rect 171502 78112 171508 78124
rect 165080 78084 171508 78112
rect 171502 78072 171508 78084
rect 171560 78072 171566 78124
rect 171686 78072 171692 78124
rect 171744 78112 171750 78124
rect 498194 78112 498200 78124
rect 171744 78084 498200 78112
rect 171744 78072 171750 78084
rect 498194 78072 498200 78084
rect 498252 78072 498258 78124
rect 145282 78044 145288 78056
rect 144840 78016 145288 78044
rect 89772 78004 89778 78016
rect 145282 78004 145288 78016
rect 145340 78004 145346 78056
rect 150710 78004 150716 78056
rect 150768 78044 150774 78056
rect 157242 78044 157248 78056
rect 150768 78016 157248 78044
rect 150768 78004 150774 78016
rect 157242 78004 157248 78016
rect 157300 78004 157306 78056
rect 168374 78004 168380 78056
rect 168432 78044 168438 78056
rect 170766 78044 170772 78056
rect 168432 78016 170772 78044
rect 168432 78004 168438 78016
rect 170766 78004 170772 78016
rect 170824 78004 170830 78056
rect 170858 78004 170864 78056
rect 170916 78044 170922 78056
rect 170916 78016 174400 78044
rect 170916 78004 170922 78016
rect 53834 77936 53840 77988
rect 53892 77976 53898 77988
rect 129734 77976 129740 77988
rect 53892 77948 129740 77976
rect 53892 77936 53898 77948
rect 129734 77936 129740 77948
rect 129792 77936 129798 77988
rect 137830 77936 137836 77988
rect 137888 77976 137894 77988
rect 138014 77976 138020 77988
rect 137888 77948 138020 77976
rect 137888 77936 137894 77948
rect 138014 77936 138020 77948
rect 138072 77936 138078 77988
rect 139486 77936 139492 77988
rect 139544 77976 139550 77988
rect 145834 77976 145840 77988
rect 139544 77948 145840 77976
rect 139544 77936 139550 77948
rect 145834 77936 145840 77948
rect 145892 77936 145898 77988
rect 154206 77936 154212 77988
rect 154264 77976 154270 77988
rect 162762 77976 162768 77988
rect 154264 77948 162768 77976
rect 154264 77936 154270 77948
rect 162762 77936 162768 77948
rect 162820 77936 162826 77988
rect 166810 77936 166816 77988
rect 166868 77976 166874 77988
rect 171870 77976 171876 77988
rect 166868 77948 171876 77976
rect 166868 77936 166874 77948
rect 171870 77936 171876 77948
rect 171928 77936 171934 77988
rect 171962 77936 171968 77988
rect 172020 77976 172026 77988
rect 174078 77976 174084 77988
rect 172020 77948 174084 77976
rect 172020 77936 172026 77948
rect 174078 77936 174084 77948
rect 174136 77936 174142 77988
rect 174372 77976 174400 78016
rect 174538 78004 174544 78056
rect 174596 78044 174602 78056
rect 574738 78044 574744 78056
rect 174596 78016 574744 78044
rect 174596 78004 174602 78016
rect 574738 78004 574744 78016
rect 574796 78004 574802 78056
rect 581086 77976 581092 77988
rect 174372 77948 581092 77976
rect 581086 77936 581092 77948
rect 581144 77936 581150 77988
rect 125318 77868 125324 77920
rect 125376 77908 125382 77920
rect 133046 77908 133052 77920
rect 125376 77880 133052 77908
rect 125376 77868 125382 77880
rect 133046 77868 133052 77880
rect 133104 77868 133110 77920
rect 141142 77868 141148 77920
rect 141200 77908 141206 77920
rect 152826 77908 152832 77920
rect 141200 77880 152832 77908
rect 141200 77868 141206 77880
rect 152826 77868 152832 77880
rect 152884 77868 152890 77920
rect 154758 77868 154764 77920
rect 154816 77908 154822 77920
rect 155586 77908 155592 77920
rect 154816 77880 155592 77908
rect 154816 77868 154822 77880
rect 155586 77868 155592 77880
rect 155644 77868 155650 77920
rect 157058 77868 157064 77920
rect 157116 77908 157122 77920
rect 171318 77908 171324 77920
rect 157116 77880 171324 77908
rect 157116 77868 157122 77880
rect 171318 77868 171324 77880
rect 171376 77868 171382 77920
rect 116578 77800 116584 77852
rect 116636 77840 116642 77852
rect 129182 77840 129188 77852
rect 116636 77812 129188 77840
rect 116636 77800 116642 77812
rect 129182 77800 129188 77812
rect 129240 77800 129246 77852
rect 129918 77800 129924 77852
rect 129976 77840 129982 77852
rect 131666 77840 131672 77852
rect 129976 77812 131672 77840
rect 129976 77800 129982 77812
rect 131666 77800 131672 77812
rect 131724 77800 131730 77852
rect 151998 77800 152004 77852
rect 152056 77840 152062 77852
rect 152550 77840 152556 77852
rect 152056 77812 152556 77840
rect 152056 77800 152062 77812
rect 152550 77800 152556 77812
rect 152608 77800 152614 77852
rect 157426 77800 157432 77852
rect 157484 77840 157490 77852
rect 171778 77840 171784 77852
rect 157484 77812 171784 77840
rect 157484 77800 157490 77812
rect 171778 77800 171784 77812
rect 171836 77800 171842 77852
rect 143534 77732 143540 77784
rect 143592 77772 143598 77784
rect 143592 77744 152504 77772
rect 143592 77732 143598 77744
rect 125410 77664 125416 77716
rect 125468 77704 125474 77716
rect 133690 77704 133696 77716
rect 125468 77676 133696 77704
rect 125468 77664 125474 77676
rect 133690 77664 133696 77676
rect 133748 77664 133754 77716
rect 152476 77704 152504 77744
rect 154574 77732 154580 77784
rect 154632 77772 154638 77784
rect 158622 77772 158628 77784
rect 154632 77744 158628 77772
rect 154632 77732 154638 77744
rect 158622 77732 158628 77744
rect 158680 77732 158686 77784
rect 159266 77732 159272 77784
rect 159324 77772 159330 77784
rect 159324 77744 160094 77772
rect 159324 77732 159330 77744
rect 159174 77704 159180 77716
rect 152476 77676 159180 77704
rect 159174 77664 159180 77676
rect 159232 77664 159238 77716
rect 160066 77704 160094 77744
rect 164878 77732 164884 77784
rect 164936 77772 164942 77784
rect 172146 77772 172152 77784
rect 164936 77744 172152 77772
rect 164936 77732 164942 77744
rect 172146 77732 172152 77744
rect 172204 77732 172210 77784
rect 171686 77704 171692 77716
rect 160066 77676 171692 77704
rect 171686 77664 171692 77676
rect 171744 77664 171750 77716
rect 122374 77596 122380 77648
rect 122432 77636 122438 77648
rect 125226 77636 125232 77648
rect 122432 77608 125232 77636
rect 122432 77596 122438 77608
rect 125226 77596 125232 77608
rect 125284 77596 125290 77648
rect 145006 77596 145012 77648
rect 145064 77636 145070 77648
rect 159266 77636 159272 77648
rect 145064 77608 159272 77636
rect 145064 77596 145070 77608
rect 159266 77596 159272 77608
rect 159324 77596 159330 77648
rect 166074 77636 166080 77648
rect 160066 77608 166080 77636
rect 120810 77528 120816 77580
rect 120868 77568 120874 77580
rect 128262 77568 128268 77580
rect 120868 77540 128268 77568
rect 120868 77528 120874 77540
rect 128262 77528 128268 77540
rect 128320 77528 128326 77580
rect 141878 77528 141884 77580
rect 141936 77568 141942 77580
rect 160066 77568 160094 77608
rect 166074 77596 166080 77608
rect 166132 77596 166138 77648
rect 169294 77596 169300 77648
rect 169352 77636 169358 77648
rect 170306 77636 170312 77648
rect 169352 77608 170312 77636
rect 169352 77596 169358 77608
rect 170306 77596 170312 77608
rect 170364 77596 170370 77648
rect 179138 77596 179144 77648
rect 179196 77636 179202 77648
rect 580074 77636 580080 77648
rect 179196 77608 580080 77636
rect 179196 77596 179202 77608
rect 580074 77596 580080 77608
rect 580132 77596 580138 77648
rect 141936 77540 160094 77568
rect 141936 77528 141942 77540
rect 164878 77528 164884 77580
rect 164936 77568 164942 77580
rect 174446 77568 174452 77580
rect 164936 77540 174452 77568
rect 164936 77528 164942 77540
rect 174446 77528 174452 77540
rect 174504 77528 174510 77580
rect 3510 77460 3516 77512
rect 3568 77500 3574 77512
rect 173986 77500 173992 77512
rect 3568 77472 173992 77500
rect 3568 77460 3574 77472
rect 173986 77460 173992 77472
rect 174044 77460 174050 77512
rect 125686 77392 125692 77444
rect 125744 77432 125750 77444
rect 135438 77432 135444 77444
rect 125744 77404 135444 77432
rect 125744 77392 125750 77404
rect 135438 77392 135444 77404
rect 135496 77392 135502 77444
rect 151446 77392 151452 77444
rect 151504 77432 151510 77444
rect 153838 77432 153844 77444
rect 151504 77404 153844 77432
rect 151504 77392 151510 77404
rect 153838 77392 153844 77404
rect 153896 77392 153902 77444
rect 159174 77392 159180 77444
rect 159232 77432 159238 77444
rect 168834 77432 168840 77444
rect 159232 77404 168840 77432
rect 159232 77392 159238 77404
rect 168834 77392 168840 77404
rect 168892 77392 168898 77444
rect 171594 77392 171600 77444
rect 171652 77432 171658 77444
rect 171778 77432 171784 77444
rect 171652 77404 171784 77432
rect 171652 77392 171658 77404
rect 171778 77392 171784 77404
rect 171836 77392 171842 77444
rect 125226 77324 125232 77376
rect 125284 77364 125290 77376
rect 132402 77364 132408 77376
rect 125284 77336 132408 77364
rect 125284 77324 125290 77336
rect 132402 77324 132408 77336
rect 132460 77324 132466 77376
rect 158346 77324 158352 77376
rect 158404 77364 158410 77376
rect 166810 77364 166816 77376
rect 158404 77336 166816 77364
rect 158404 77324 158410 77336
rect 166810 77324 166816 77336
rect 166868 77324 166874 77376
rect 126238 77256 126244 77308
rect 126296 77296 126302 77308
rect 130562 77296 130568 77308
rect 126296 77268 130568 77296
rect 126296 77256 126302 77268
rect 130562 77256 130568 77268
rect 130620 77256 130626 77308
rect 151814 77256 151820 77308
rect 151872 77296 151878 77308
rect 152734 77296 152740 77308
rect 151872 77268 152740 77296
rect 151872 77256 151878 77268
rect 152734 77256 152740 77268
rect 152792 77256 152798 77308
rect 158806 77256 158812 77308
rect 158864 77296 158870 77308
rect 158990 77296 158996 77308
rect 158864 77268 158996 77296
rect 158864 77256 158870 77268
rect 158990 77256 158996 77268
rect 159048 77256 159054 77308
rect 159266 77256 159272 77308
rect 159324 77296 159330 77308
rect 164878 77296 164884 77308
rect 159324 77268 164884 77296
rect 159324 77256 159330 77268
rect 164878 77256 164884 77268
rect 164936 77256 164942 77308
rect 166626 77256 166632 77308
rect 166684 77296 166690 77308
rect 170490 77296 170496 77308
rect 166684 77268 170496 77296
rect 166684 77256 166690 77268
rect 170490 77256 170496 77268
rect 170548 77256 170554 77308
rect 125870 77188 125876 77240
rect 125928 77228 125934 77240
rect 126790 77228 126796 77240
rect 125928 77200 126796 77228
rect 125928 77188 125934 77200
rect 126790 77188 126796 77200
rect 126848 77188 126854 77240
rect 127158 77188 127164 77240
rect 127216 77228 127222 77240
rect 127434 77228 127440 77240
rect 127216 77200 127440 77228
rect 127216 77188 127222 77200
rect 127434 77188 127440 77200
rect 127492 77188 127498 77240
rect 127526 77188 127532 77240
rect 127584 77228 127590 77240
rect 127802 77228 127808 77240
rect 127584 77200 127808 77228
rect 127584 77188 127590 77200
rect 127802 77188 127808 77200
rect 127860 77188 127866 77240
rect 128078 77188 128084 77240
rect 128136 77228 128142 77240
rect 128354 77228 128360 77240
rect 128136 77200 128360 77228
rect 128136 77188 128142 77200
rect 128354 77188 128360 77200
rect 128412 77188 128418 77240
rect 151998 77188 152004 77240
rect 152056 77228 152062 77240
rect 152458 77228 152464 77240
rect 152056 77200 152464 77228
rect 152056 77188 152062 77200
rect 152458 77188 152464 77200
rect 152516 77188 152522 77240
rect 154298 77188 154304 77240
rect 154356 77228 154362 77240
rect 155770 77228 155776 77240
rect 154356 77200 155776 77228
rect 154356 77188 154362 77200
rect 155770 77188 155776 77200
rect 155828 77188 155834 77240
rect 160278 77188 160284 77240
rect 160336 77228 160342 77240
rect 160830 77228 160836 77240
rect 160336 77200 160836 77228
rect 160336 77188 160342 77200
rect 160830 77188 160836 77200
rect 160888 77188 160894 77240
rect 163038 77188 163044 77240
rect 163096 77228 163102 77240
rect 163590 77228 163596 77240
rect 163096 77200 163596 77228
rect 163096 77188 163102 77200
rect 163590 77188 163596 77200
rect 163648 77188 163654 77240
rect 163958 77188 163964 77240
rect 164016 77228 164022 77240
rect 169294 77228 169300 77240
rect 164016 77200 169300 77228
rect 164016 77188 164022 77200
rect 169294 77188 169300 77200
rect 169352 77188 169358 77240
rect 172330 77188 172336 77240
rect 172388 77228 172394 77240
rect 527174 77228 527180 77240
rect 172388 77200 527180 77228
rect 172388 77188 172394 77200
rect 527174 77188 527180 77200
rect 527232 77188 527238 77240
rect 143626 77120 143632 77172
rect 143684 77160 143690 77172
rect 143902 77160 143908 77172
rect 143684 77132 143908 77160
rect 143684 77120 143690 77132
rect 143902 77120 143908 77132
rect 143960 77120 143966 77172
rect 152734 77120 152740 77172
rect 152792 77160 152798 77172
rect 226334 77160 226340 77172
rect 152792 77132 226340 77160
rect 152792 77120 152798 77132
rect 226334 77120 226340 77132
rect 226392 77120 226398 77172
rect 149238 77052 149244 77104
rect 149296 77092 149302 77104
rect 149514 77092 149520 77104
rect 149296 77064 149520 77092
rect 149296 77052 149302 77064
rect 149514 77052 149520 77064
rect 149572 77052 149578 77104
rect 152458 77052 152464 77104
rect 152516 77092 152522 77104
rect 240134 77092 240140 77104
rect 152516 77064 240140 77092
rect 152516 77052 152522 77064
rect 240134 77052 240140 77064
rect 240192 77052 240198 77104
rect 129090 76984 129096 77036
rect 129148 77024 129154 77036
rect 130194 77024 130200 77036
rect 129148 76996 130200 77024
rect 129148 76984 129154 76996
rect 130194 76984 130200 76996
rect 130252 76984 130258 77036
rect 145926 76984 145932 77036
rect 145984 77024 145990 77036
rect 260834 77024 260840 77036
rect 145984 76996 260840 77024
rect 145984 76984 145990 76996
rect 260834 76984 260840 76996
rect 260892 76984 260898 77036
rect 146110 76916 146116 76968
rect 146168 76956 146174 76968
rect 267734 76956 267740 76968
rect 146168 76928 267740 76956
rect 146168 76916 146174 76928
rect 267734 76916 267740 76928
rect 267792 76916 267798 76968
rect 133046 76848 133052 76900
rect 133104 76888 133110 76900
rect 135530 76888 135536 76900
rect 133104 76860 135536 76888
rect 133104 76848 133110 76860
rect 135530 76848 135536 76860
rect 135588 76848 135594 76900
rect 143994 76848 144000 76900
rect 144052 76888 144058 76900
rect 144178 76888 144184 76900
rect 144052 76860 144184 76888
rect 144052 76848 144058 76860
rect 144178 76848 144184 76860
rect 144236 76848 144242 76900
rect 146570 76848 146576 76900
rect 146628 76888 146634 76900
rect 147030 76888 147036 76900
rect 146628 76860 147036 76888
rect 146628 76848 146634 76860
rect 147030 76848 147036 76860
rect 147088 76848 147094 76900
rect 148042 76848 148048 76900
rect 148100 76888 148106 76900
rect 288434 76888 288440 76900
rect 148100 76860 288440 76888
rect 148100 76848 148106 76860
rect 288434 76848 288440 76860
rect 288492 76848 288498 76900
rect 122834 76780 122840 76832
rect 122892 76820 122898 76832
rect 133322 76820 133328 76832
rect 122892 76792 133328 76820
rect 122892 76780 122898 76792
rect 133322 76780 133328 76792
rect 133380 76780 133386 76832
rect 143902 76780 143908 76832
rect 143960 76820 143966 76832
rect 144086 76820 144092 76832
rect 143960 76792 144092 76820
rect 143960 76780 143966 76792
rect 144086 76780 144092 76792
rect 144144 76780 144150 76832
rect 148594 76780 148600 76832
rect 148652 76820 148658 76832
rect 296714 76820 296720 76832
rect 148652 76792 296720 76820
rect 148652 76780 148658 76792
rect 296714 76780 296720 76792
rect 296772 76780 296778 76832
rect 118694 76712 118700 76764
rect 118752 76752 118758 76764
rect 133782 76752 133788 76764
rect 118752 76724 133788 76752
rect 118752 76712 118758 76724
rect 133782 76712 133788 76724
rect 133840 76712 133846 76764
rect 136910 76712 136916 76764
rect 136968 76752 136974 76764
rect 137094 76752 137100 76764
rect 136968 76724 137100 76752
rect 136968 76712 136974 76724
rect 137094 76712 137100 76724
rect 137152 76712 137158 76764
rect 138842 76712 138848 76764
rect 138900 76752 138906 76764
rect 139302 76752 139308 76764
rect 138900 76724 139308 76752
rect 138900 76712 138906 76724
rect 139302 76712 139308 76724
rect 139360 76712 139366 76764
rect 139486 76712 139492 76764
rect 139544 76752 139550 76764
rect 140038 76752 140044 76764
rect 139544 76724 140044 76752
rect 139544 76712 139550 76724
rect 140038 76712 140044 76724
rect 140096 76712 140102 76764
rect 143810 76712 143816 76764
rect 143868 76752 143874 76764
rect 143994 76752 144000 76764
rect 143868 76724 144000 76752
rect 143868 76712 143874 76724
rect 143994 76712 144000 76724
rect 144052 76712 144058 76764
rect 146202 76712 146208 76764
rect 146260 76752 146266 76764
rect 146662 76752 146668 76764
rect 146260 76724 146668 76752
rect 146260 76712 146266 76724
rect 146662 76712 146668 76724
rect 146720 76712 146726 76764
rect 149146 76712 149152 76764
rect 149204 76752 149210 76764
rect 302234 76752 302240 76764
rect 149204 76724 302240 76752
rect 149204 76712 149210 76724
rect 302234 76712 302240 76724
rect 302292 76712 302298 76764
rect 93854 76644 93860 76696
rect 93912 76684 93918 76696
rect 130930 76684 130936 76696
rect 93912 76656 130936 76684
rect 93912 76644 93918 76656
rect 130930 76644 130936 76656
rect 130988 76644 130994 76696
rect 132402 76644 132408 76696
rect 132460 76684 132466 76696
rect 140498 76684 140504 76696
rect 132460 76656 140504 76684
rect 132460 76644 132466 76656
rect 140498 76644 140504 76656
rect 140556 76644 140562 76696
rect 142890 76644 142896 76696
rect 142948 76684 142954 76696
rect 142948 76656 148456 76684
rect 142948 76644 142954 76656
rect 70394 76576 70400 76628
rect 70452 76616 70458 76628
rect 131022 76616 131028 76628
rect 70452 76588 131028 76616
rect 70452 76576 70458 76588
rect 131022 76576 131028 76588
rect 131080 76576 131086 76628
rect 131758 76576 131764 76628
rect 131816 76616 131822 76628
rect 132034 76616 132040 76628
rect 131816 76588 132040 76616
rect 131816 76576 131822 76588
rect 132034 76576 132040 76588
rect 132092 76576 132098 76628
rect 132678 76576 132684 76628
rect 132736 76616 132742 76628
rect 133230 76616 133236 76628
rect 132736 76588 133236 76616
rect 132736 76576 132742 76588
rect 133230 76576 133236 76588
rect 133288 76576 133294 76628
rect 133414 76576 133420 76628
rect 133472 76616 133478 76628
rect 133690 76616 133696 76628
rect 133472 76588 133696 76616
rect 133472 76576 133478 76588
rect 133690 76576 133696 76588
rect 133748 76576 133754 76628
rect 135806 76576 135812 76628
rect 135864 76616 135870 76628
rect 136450 76616 136456 76628
rect 135864 76588 136456 76616
rect 135864 76576 135870 76588
rect 136450 76576 136456 76588
rect 136508 76576 136514 76628
rect 138290 76576 138296 76628
rect 138348 76616 138354 76628
rect 138842 76616 138848 76628
rect 138348 76588 138848 76616
rect 138348 76576 138354 76588
rect 138842 76576 138848 76588
rect 138900 76576 138906 76628
rect 140774 76576 140780 76628
rect 140832 76616 140838 76628
rect 141694 76616 141700 76628
rect 140832 76588 141700 76616
rect 140832 76576 140838 76588
rect 141694 76576 141700 76588
rect 141752 76576 141758 76628
rect 143810 76576 143816 76628
rect 143868 76616 143874 76628
rect 144454 76616 144460 76628
rect 143868 76588 144460 76616
rect 143868 76576 143874 76588
rect 144454 76576 144460 76588
rect 144512 76576 144518 76628
rect 145006 76576 145012 76628
rect 145064 76616 145070 76628
rect 145374 76616 145380 76628
rect 145064 76588 145380 76616
rect 145064 76576 145070 76588
rect 145374 76576 145380 76588
rect 145432 76576 145438 76628
rect 146386 76576 146392 76628
rect 146444 76616 146450 76628
rect 146662 76616 146668 76628
rect 146444 76588 146668 76616
rect 146444 76576 146450 76588
rect 146662 76576 146668 76588
rect 146720 76576 146726 76628
rect 148042 76576 148048 76628
rect 148100 76616 148106 76628
rect 148318 76616 148324 76628
rect 148100 76588 148324 76616
rect 148100 76576 148106 76588
rect 148318 76576 148324 76588
rect 148376 76576 148382 76628
rect 148428 76616 148456 76656
rect 149330 76644 149336 76696
rect 149388 76684 149394 76696
rect 149882 76684 149888 76696
rect 149388 76656 149888 76684
rect 149388 76644 149394 76656
rect 149882 76644 149888 76656
rect 149940 76644 149946 76696
rect 150250 76644 150256 76696
rect 150308 76684 150314 76696
rect 152458 76684 152464 76696
rect 150308 76656 152464 76684
rect 150308 76644 150314 76656
rect 152458 76644 152464 76656
rect 152516 76644 152522 76696
rect 154390 76644 154396 76696
rect 154448 76684 154454 76696
rect 356054 76684 356060 76696
rect 154448 76656 356060 76684
rect 154448 76644 154454 76656
rect 356054 76644 356060 76656
rect 356112 76644 356118 76696
rect 152734 76616 152740 76628
rect 148428 76588 152740 76616
rect 152734 76576 152740 76588
rect 152792 76576 152798 76628
rect 159266 76576 159272 76628
rect 159324 76616 159330 76628
rect 159542 76616 159548 76628
rect 159324 76588 159548 76616
rect 159324 76576 159330 76588
rect 159542 76576 159548 76588
rect 159600 76576 159606 76628
rect 160186 76576 160192 76628
rect 160244 76616 160250 76628
rect 160370 76616 160376 76628
rect 160244 76588 160376 76616
rect 160244 76576 160250 76588
rect 160370 76576 160376 76588
rect 160428 76576 160434 76628
rect 160462 76576 160468 76628
rect 160520 76616 160526 76628
rect 160646 76616 160652 76628
rect 160520 76588 160652 76616
rect 160520 76576 160526 76588
rect 160646 76576 160652 76588
rect 160704 76576 160710 76628
rect 161566 76576 161572 76628
rect 161624 76616 161630 76628
rect 162210 76616 162216 76628
rect 161624 76588 162216 76616
rect 161624 76576 161630 76588
rect 162210 76576 162216 76588
rect 162268 76576 162274 76628
rect 163038 76576 163044 76628
rect 163096 76616 163102 76628
rect 163498 76616 163504 76628
rect 163096 76588 163504 76616
rect 163096 76576 163102 76588
rect 163498 76576 163504 76588
rect 163556 76576 163562 76628
rect 165798 76576 165804 76628
rect 165856 76616 165862 76628
rect 166350 76616 166356 76628
rect 165856 76588 166356 76616
rect 165856 76576 165862 76588
rect 166350 76576 166356 76588
rect 166408 76576 166414 76628
rect 166442 76576 166448 76628
rect 166500 76616 166506 76628
rect 166626 76616 166632 76628
rect 166500 76588 166632 76616
rect 166500 76576 166506 76588
rect 166626 76576 166632 76588
rect 166684 76576 166690 76628
rect 167638 76576 167644 76628
rect 167696 76616 167702 76628
rect 167822 76616 167828 76628
rect 167696 76588 167828 76616
rect 167696 76576 167702 76588
rect 167822 76576 167828 76588
rect 167880 76576 167886 76628
rect 168650 76576 168656 76628
rect 168708 76616 168714 76628
rect 169386 76616 169392 76628
rect 168708 76588 169392 76616
rect 168708 76576 168714 76588
rect 169386 76576 169392 76588
rect 169444 76576 169450 76628
rect 171778 76616 171784 76628
rect 169726 76588 171784 76616
rect 69014 76508 69020 76560
rect 69072 76548 69078 76560
rect 131114 76548 131120 76560
rect 69072 76520 131120 76548
rect 69072 76508 69078 76520
rect 131114 76508 131120 76520
rect 131172 76508 131178 76560
rect 139578 76508 139584 76560
rect 139636 76548 139642 76560
rect 139946 76548 139952 76560
rect 139636 76520 139952 76548
rect 139636 76508 139642 76520
rect 139946 76508 139952 76520
rect 140004 76508 140010 76560
rect 141234 76508 141240 76560
rect 141292 76548 141298 76560
rect 141510 76548 141516 76560
rect 141292 76520 141516 76548
rect 141292 76508 141298 76520
rect 141510 76508 141516 76520
rect 141568 76508 141574 76560
rect 142246 76508 142252 76560
rect 142304 76548 142310 76560
rect 142798 76548 142804 76560
rect 142304 76520 142804 76548
rect 142304 76508 142310 76520
rect 142798 76508 142804 76520
rect 142856 76508 142862 76560
rect 146846 76508 146852 76560
rect 146904 76548 146910 76560
rect 147122 76548 147128 76560
rect 146904 76520 147128 76548
rect 146904 76508 146910 76520
rect 147122 76508 147128 76520
rect 147180 76508 147186 76560
rect 149238 76508 149244 76560
rect 149296 76548 149302 76560
rect 149698 76548 149704 76560
rect 149296 76520 149704 76548
rect 149296 76508 149302 76520
rect 149698 76508 149704 76520
rect 149756 76508 149762 76560
rect 152458 76508 152464 76560
rect 152516 76548 152522 76560
rect 152918 76548 152924 76560
rect 152516 76520 152924 76548
rect 152516 76508 152522 76520
rect 152918 76508 152924 76520
rect 152976 76508 152982 76560
rect 161658 76508 161664 76560
rect 161716 76548 161722 76560
rect 162302 76548 162308 76560
rect 161716 76520 162308 76548
rect 161716 76508 161722 76520
rect 162302 76508 162308 76520
rect 162360 76508 162366 76560
rect 164326 76508 164332 76560
rect 164384 76548 164390 76560
rect 164786 76548 164792 76560
rect 164384 76520 164792 76548
rect 164384 76508 164390 76520
rect 164786 76508 164792 76520
rect 164844 76508 164850 76560
rect 168374 76508 168380 76560
rect 168432 76548 168438 76560
rect 169110 76548 169116 76560
rect 168432 76520 169116 76548
rect 168432 76508 168438 76520
rect 169110 76508 169116 76520
rect 169168 76508 169174 76560
rect 169294 76508 169300 76560
rect 169352 76548 169358 76560
rect 169726 76548 169754 76588
rect 171778 76576 171784 76588
rect 171836 76576 171842 76628
rect 172146 76576 172152 76628
rect 172204 76616 172210 76628
rect 557534 76616 557540 76628
rect 172204 76588 557540 76616
rect 172204 76576 172210 76588
rect 557534 76576 557540 76588
rect 557592 76576 557598 76628
rect 169352 76520 169754 76548
rect 169352 76508 169358 76520
rect 170306 76508 170312 76560
rect 170364 76548 170370 76560
rect 558914 76548 558920 76560
rect 170364 76520 558920 76548
rect 170364 76508 170370 76520
rect 558914 76508 558920 76520
rect 558972 76508 558978 76560
rect 131022 76440 131028 76492
rect 131080 76480 131086 76492
rect 132586 76480 132592 76492
rect 131080 76452 132592 76480
rect 131080 76440 131086 76452
rect 132586 76440 132592 76452
rect 132644 76440 132650 76492
rect 137922 76440 137928 76492
rect 137980 76480 137986 76492
rect 138658 76480 138664 76492
rect 137980 76452 138664 76480
rect 137980 76440 137986 76452
rect 138658 76440 138664 76452
rect 138716 76440 138722 76492
rect 139762 76440 139768 76492
rect 139820 76480 139826 76492
rect 182174 76480 182180 76492
rect 139820 76452 182180 76480
rect 139820 76440 139826 76452
rect 182174 76440 182180 76452
rect 182232 76440 182238 76492
rect 124858 76372 124864 76424
rect 124916 76412 124922 76424
rect 131574 76412 131580 76424
rect 124916 76384 131580 76412
rect 124916 76372 124922 76384
rect 131574 76372 131580 76384
rect 131632 76372 131638 76424
rect 145374 76372 145380 76424
rect 145432 76412 145438 76424
rect 145650 76412 145656 76424
rect 145432 76384 145656 76412
rect 145432 76372 145438 76384
rect 145650 76372 145656 76384
rect 145708 76372 145714 76424
rect 145834 76372 145840 76424
rect 145892 76412 145898 76424
rect 178034 76412 178040 76424
rect 145892 76384 178040 76412
rect 145892 76372 145898 76384
rect 178034 76372 178040 76384
rect 178092 76372 178098 76424
rect 139762 76304 139768 76356
rect 139820 76344 139826 76356
rect 140222 76344 140228 76356
rect 139820 76316 140228 76344
rect 139820 76304 139826 76316
rect 140222 76304 140228 76316
rect 140280 76304 140286 76356
rect 147766 76304 147772 76356
rect 147824 76344 147830 76356
rect 148318 76344 148324 76356
rect 147824 76316 148324 76344
rect 147824 76304 147830 76316
rect 148318 76304 148324 76316
rect 148376 76304 148382 76356
rect 150894 76304 150900 76356
rect 150952 76344 150958 76356
rect 151446 76344 151452 76356
rect 150952 76316 151452 76344
rect 150952 76304 150958 76316
rect 151446 76304 151452 76316
rect 151504 76304 151510 76356
rect 160370 76304 160376 76356
rect 160428 76344 160434 76356
rect 160738 76344 160744 76356
rect 160428 76316 160744 76344
rect 160428 76304 160434 76316
rect 160738 76304 160744 76316
rect 160796 76304 160802 76356
rect 161474 76304 161480 76356
rect 161532 76344 161538 76356
rect 167822 76344 167828 76356
rect 161532 76316 167828 76344
rect 161532 76304 161538 76316
rect 167822 76304 167828 76316
rect 167880 76304 167886 76356
rect 168466 76304 168472 76356
rect 168524 76344 168530 76356
rect 168834 76344 168840 76356
rect 168524 76316 168840 76344
rect 168524 76304 168530 76316
rect 168834 76304 168840 76316
rect 168892 76304 168898 76356
rect 171502 76304 171508 76356
rect 171560 76344 171566 76356
rect 195974 76344 195980 76356
rect 171560 76316 195980 76344
rect 171560 76304 171566 76316
rect 195974 76304 195980 76316
rect 196032 76304 196038 76356
rect 125134 76236 125140 76288
rect 125192 76276 125198 76288
rect 126698 76276 126704 76288
rect 125192 76248 126704 76276
rect 125192 76236 125198 76248
rect 126698 76236 126704 76248
rect 126756 76236 126762 76288
rect 131574 76236 131580 76288
rect 131632 76276 131638 76288
rect 131942 76276 131948 76288
rect 131632 76248 131948 76276
rect 131632 76236 131638 76248
rect 131942 76236 131948 76248
rect 132000 76236 132006 76288
rect 135622 76236 135628 76288
rect 135680 76276 135686 76288
rect 136634 76276 136640 76288
rect 135680 76248 136640 76276
rect 135680 76236 135686 76248
rect 136634 76236 136640 76248
rect 136692 76236 136698 76288
rect 164142 76236 164148 76288
rect 164200 76276 164206 76288
rect 164418 76276 164424 76288
rect 164200 76248 164424 76276
rect 164200 76236 164206 76248
rect 164418 76236 164424 76248
rect 164476 76236 164482 76288
rect 166994 76236 167000 76288
rect 167052 76276 167058 76288
rect 167914 76276 167920 76288
rect 167052 76248 167920 76276
rect 167052 76236 167058 76248
rect 167914 76236 167920 76248
rect 167972 76236 167978 76288
rect 160462 76168 160468 76220
rect 160520 76208 160526 76220
rect 161014 76208 161020 76220
rect 160520 76180 161020 76208
rect 160520 76168 160526 76180
rect 161014 76168 161020 76180
rect 161072 76168 161078 76220
rect 168466 76168 168472 76220
rect 168524 76208 168530 76220
rect 169018 76208 169024 76220
rect 168524 76180 169024 76208
rect 168524 76168 168530 76180
rect 169018 76168 169024 76180
rect 169076 76168 169082 76220
rect 128722 76100 128728 76152
rect 128780 76140 128786 76152
rect 129458 76140 129464 76152
rect 128780 76112 129464 76140
rect 128780 76100 128786 76112
rect 129458 76100 129464 76112
rect 129516 76100 129522 76152
rect 136634 76100 136640 76152
rect 136692 76140 136698 76152
rect 137738 76140 137744 76152
rect 136692 76112 137744 76140
rect 136692 76100 136698 76112
rect 137738 76100 137744 76112
rect 137796 76100 137802 76152
rect 144914 76100 144920 76152
rect 144972 76140 144978 76152
rect 146018 76140 146024 76152
rect 144972 76112 146024 76140
rect 144972 76100 144978 76112
rect 146018 76100 146024 76112
rect 146076 76100 146082 76152
rect 159450 76100 159456 76152
rect 159508 76140 159514 76152
rect 159818 76140 159824 76152
rect 159508 76112 159824 76140
rect 159508 76100 159514 76112
rect 159818 76100 159824 76112
rect 159876 76100 159882 76152
rect 160738 76100 160744 76152
rect 160796 76140 160802 76152
rect 160922 76140 160928 76152
rect 160796 76112 160928 76140
rect 160796 76100 160802 76112
rect 160922 76100 160928 76112
rect 160980 76100 160986 76152
rect 165706 76100 165712 76152
rect 165764 76140 165770 76152
rect 166258 76140 166264 76152
rect 165764 76112 166264 76140
rect 165764 76100 165770 76112
rect 166258 76100 166264 76112
rect 166316 76100 166322 76152
rect 125042 76032 125048 76084
rect 125100 76072 125106 76084
rect 126974 76072 126980 76084
rect 125100 76044 126980 76072
rect 125100 76032 125106 76044
rect 126974 76032 126980 76044
rect 127032 76032 127038 76084
rect 129734 76032 129740 76084
rect 129792 76072 129798 76084
rect 135898 76072 135904 76084
rect 129792 76044 135904 76072
rect 129792 76032 129798 76044
rect 135898 76032 135904 76044
rect 135956 76032 135962 76084
rect 131482 75964 131488 76016
rect 131540 76004 131546 76016
rect 132126 76004 132132 76016
rect 131540 75976 132132 76004
rect 131540 75964 131546 75976
rect 132126 75964 132132 75976
rect 132184 75964 132190 76016
rect 163130 75964 163136 76016
rect 163188 76004 163194 76016
rect 163866 76004 163872 76016
rect 163188 75976 163872 76004
rect 163188 75964 163194 75976
rect 163866 75964 163872 75976
rect 163924 75964 163930 76016
rect 137370 75896 137376 75948
rect 137428 75936 137434 75948
rect 144454 75936 144460 75948
rect 137428 75908 144460 75936
rect 137428 75896 137434 75908
rect 144454 75896 144460 75908
rect 144512 75896 144518 75948
rect 153378 75896 153384 75948
rect 153436 75936 153442 75948
rect 153562 75936 153568 75948
rect 153436 75908 153568 75936
rect 153436 75896 153442 75908
rect 153562 75896 153568 75908
rect 153620 75896 153626 75948
rect 170950 75896 170956 75948
rect 171008 75936 171014 75948
rect 173342 75936 173348 75948
rect 171008 75908 173348 75936
rect 171008 75896 171014 75908
rect 173342 75896 173348 75908
rect 173400 75896 173406 75948
rect 134058 75828 134064 75880
rect 134116 75868 134122 75880
rect 134702 75868 134708 75880
rect 134116 75840 134708 75868
rect 134116 75828 134122 75840
rect 134702 75828 134708 75840
rect 134760 75828 134766 75880
rect 130378 75760 130384 75812
rect 130436 75800 130442 75812
rect 133046 75800 133052 75812
rect 130436 75772 133052 75800
rect 130436 75760 130442 75772
rect 133046 75760 133052 75772
rect 133104 75760 133110 75812
rect 129182 75692 129188 75744
rect 129240 75732 129246 75744
rect 129550 75732 129556 75744
rect 129240 75704 129556 75732
rect 129240 75692 129246 75704
rect 129550 75692 129556 75704
rect 129608 75692 129614 75744
rect 159634 75692 159640 75744
rect 159692 75732 159698 75744
rect 164878 75732 164884 75744
rect 159692 75704 164884 75732
rect 159692 75692 159698 75704
rect 164878 75692 164884 75704
rect 164936 75692 164942 75744
rect 155034 75624 155040 75676
rect 155092 75664 155098 75676
rect 155310 75664 155316 75676
rect 155092 75636 155316 75664
rect 155092 75624 155098 75636
rect 155310 75624 155316 75636
rect 155368 75624 155374 75676
rect 157334 75624 157340 75676
rect 157392 75664 157398 75676
rect 157886 75664 157892 75676
rect 157392 75636 157892 75664
rect 157392 75624 157398 75636
rect 157886 75624 157892 75636
rect 157944 75624 157950 75676
rect 160066 75636 173894 75664
rect 125778 75488 125784 75540
rect 125836 75528 125842 75540
rect 126606 75528 126612 75540
rect 125836 75500 126612 75528
rect 125836 75488 125842 75500
rect 126606 75488 126612 75500
rect 126664 75488 126670 75540
rect 128538 75488 128544 75540
rect 128596 75528 128602 75540
rect 129918 75528 129924 75540
rect 128596 75500 129924 75528
rect 128596 75488 128602 75500
rect 129918 75488 129924 75500
rect 129976 75488 129982 75540
rect 135530 75488 135536 75540
rect 135588 75528 135594 75540
rect 136266 75528 136272 75540
rect 135588 75500 136272 75528
rect 135588 75488 135594 75500
rect 136266 75488 136272 75500
rect 136324 75488 136330 75540
rect 142522 75488 142528 75540
rect 142580 75528 142586 75540
rect 142706 75528 142712 75540
rect 142580 75500 142712 75528
rect 142580 75488 142586 75500
rect 142706 75488 142712 75500
rect 142764 75488 142770 75540
rect 152826 75488 152832 75540
rect 152884 75528 152890 75540
rect 160066 75528 160094 75636
rect 167454 75556 167460 75608
rect 167512 75596 167518 75608
rect 167822 75596 167828 75608
rect 167512 75568 167828 75596
rect 167512 75556 167518 75568
rect 167822 75556 167828 75568
rect 167880 75556 167886 75608
rect 152884 75500 160094 75528
rect 173866 75528 173894 75636
rect 197354 75528 197360 75540
rect 173866 75500 197360 75528
rect 152884 75488 152890 75500
rect 197354 75488 197360 75500
rect 197412 75488 197418 75540
rect 123570 75420 123576 75472
rect 123628 75460 123634 75472
rect 130102 75460 130108 75472
rect 123628 75432 130108 75460
rect 123628 75420 123634 75432
rect 130102 75420 130108 75432
rect 130160 75420 130166 75472
rect 153654 75420 153660 75472
rect 153712 75460 153718 75472
rect 155586 75460 155592 75472
rect 153712 75432 155592 75460
rect 153712 75420 153718 75432
rect 155586 75420 155592 75432
rect 155644 75420 155650 75472
rect 167086 75420 167092 75472
rect 167144 75460 167150 75472
rect 167454 75460 167460 75472
rect 167144 75432 167460 75460
rect 167144 75420 167150 75432
rect 167454 75420 167460 75432
rect 167512 75420 167518 75472
rect 171134 75420 171140 75472
rect 171192 75460 171198 75472
rect 358814 75460 358820 75472
rect 171192 75432 358820 75460
rect 171192 75420 171198 75432
rect 358814 75420 358820 75432
rect 358872 75420 358878 75472
rect 107654 75352 107660 75404
rect 107712 75392 107718 75404
rect 132218 75392 132224 75404
rect 107712 75364 132224 75392
rect 107712 75352 107718 75364
rect 132218 75352 132224 75364
rect 132276 75352 132282 75404
rect 142522 75352 142528 75404
rect 142580 75392 142586 75404
rect 143074 75392 143080 75404
rect 142580 75364 143080 75392
rect 142580 75352 142586 75364
rect 143074 75352 143080 75364
rect 143132 75352 143138 75404
rect 157334 75352 157340 75404
rect 157392 75392 157398 75404
rect 157702 75392 157708 75404
rect 157392 75364 157708 75392
rect 157392 75352 157398 75364
rect 157702 75352 157708 75364
rect 157760 75352 157766 75404
rect 164878 75352 164884 75404
rect 164936 75392 164942 75404
rect 438854 75392 438860 75404
rect 164936 75364 438860 75392
rect 164936 75352 164942 75364
rect 438854 75352 438860 75364
rect 438912 75352 438918 75404
rect 51074 75284 51080 75336
rect 51132 75324 51138 75336
rect 125502 75324 125508 75336
rect 51132 75296 125508 75324
rect 51132 75284 51138 75296
rect 125502 75284 125508 75296
rect 125560 75284 125566 75336
rect 129274 75324 129280 75336
rect 125796 75296 129280 75324
rect 49694 75216 49700 75268
rect 49752 75256 49758 75268
rect 125796 75256 125824 75296
rect 129274 75284 129280 75296
rect 129332 75284 129338 75336
rect 134334 75284 134340 75336
rect 134392 75324 134398 75336
rect 134610 75324 134616 75336
rect 134392 75296 134616 75324
rect 134392 75284 134398 75296
rect 134610 75284 134616 75296
rect 134668 75284 134674 75336
rect 150710 75284 150716 75336
rect 150768 75324 150774 75336
rect 151078 75324 151084 75336
rect 150768 75296 151084 75324
rect 150768 75284 150774 75296
rect 151078 75284 151084 75296
rect 151136 75284 151142 75336
rect 154574 75284 154580 75336
rect 154632 75324 154638 75336
rect 155494 75324 155500 75336
rect 154632 75296 155500 75324
rect 154632 75284 154638 75296
rect 155494 75284 155500 75296
rect 155552 75284 155558 75336
rect 156046 75284 156052 75336
rect 156104 75324 156110 75336
rect 156598 75324 156604 75336
rect 156104 75296 156604 75324
rect 156104 75284 156110 75296
rect 156598 75284 156604 75296
rect 156656 75284 156662 75336
rect 163774 75284 163780 75336
rect 163832 75324 163838 75336
rect 489914 75324 489920 75336
rect 163832 75296 489920 75324
rect 163832 75284 163838 75296
rect 489914 75284 489920 75296
rect 489972 75284 489978 75336
rect 49752 75228 125824 75256
rect 49752 75216 49758 75228
rect 150802 75216 150808 75268
rect 150860 75256 150866 75268
rect 151262 75256 151268 75268
rect 150860 75228 151268 75256
rect 150860 75216 150866 75228
rect 151262 75216 151268 75228
rect 151320 75216 151326 75268
rect 154942 75216 154948 75268
rect 155000 75256 155006 75268
rect 155218 75256 155224 75268
rect 155000 75228 155224 75256
rect 155000 75216 155006 75228
rect 155218 75216 155224 75228
rect 155276 75216 155282 75268
rect 156322 75216 156328 75268
rect 156380 75256 156386 75268
rect 156506 75256 156512 75268
rect 156380 75228 156512 75256
rect 156380 75216 156386 75228
rect 156506 75216 156512 75228
rect 156564 75216 156570 75268
rect 157702 75216 157708 75268
rect 157760 75256 157766 75268
rect 158162 75256 158168 75268
rect 157760 75228 158168 75256
rect 157760 75216 157766 75228
rect 158162 75216 158168 75228
rect 158220 75216 158226 75268
rect 167822 75216 167828 75268
rect 167880 75256 167886 75268
rect 506474 75256 506480 75268
rect 167880 75228 506480 75256
rect 167880 75216 167886 75228
rect 506474 75216 506480 75228
rect 506532 75216 506538 75268
rect 46934 75148 46940 75200
rect 46992 75188 46998 75200
rect 46992 75160 118694 75188
rect 46992 75148 46998 75160
rect 118666 75052 118694 75160
rect 134150 75148 134156 75200
rect 134208 75188 134214 75200
rect 135162 75188 135168 75200
rect 134208 75160 135168 75188
rect 134208 75148 134214 75160
rect 135162 75148 135168 75160
rect 135220 75148 135226 75200
rect 150894 75148 150900 75200
rect 150952 75188 150958 75200
rect 151354 75188 151360 75200
rect 150952 75160 151360 75188
rect 150952 75148 150958 75160
rect 151354 75148 151360 75160
rect 151412 75148 151418 75200
rect 155034 75148 155040 75200
rect 155092 75188 155098 75200
rect 155402 75188 155408 75200
rect 155092 75160 155408 75188
rect 155092 75148 155098 75160
rect 155402 75148 155408 75160
rect 155460 75148 155466 75200
rect 156046 75148 156052 75200
rect 156104 75188 156110 75200
rect 156966 75188 156972 75200
rect 156104 75160 156972 75188
rect 156104 75148 156110 75160
rect 156966 75148 156972 75160
rect 157024 75148 157030 75200
rect 157518 75148 157524 75200
rect 157576 75188 157582 75200
rect 158254 75188 158260 75200
rect 157576 75160 158260 75188
rect 157576 75148 157582 75160
rect 158254 75148 158260 75160
rect 158312 75148 158318 75200
rect 168006 75148 168012 75200
rect 168064 75188 168070 75200
rect 517514 75188 517520 75200
rect 168064 75160 517520 75188
rect 168064 75148 168070 75160
rect 517514 75148 517520 75160
rect 517572 75148 517578 75200
rect 147766 75080 147772 75132
rect 147824 75120 147830 75132
rect 148410 75120 148416 75132
rect 147824 75092 148416 75120
rect 147824 75080 147830 75092
rect 148410 75080 148416 75092
rect 148468 75080 148474 75132
rect 152182 75080 152188 75132
rect 152240 75120 152246 75132
rect 152642 75120 152648 75132
rect 152240 75092 152648 75120
rect 152240 75080 152246 75092
rect 152642 75080 152648 75092
rect 152700 75080 152706 75132
rect 153562 75080 153568 75132
rect 153620 75120 153626 75132
rect 154114 75120 154120 75132
rect 153620 75092 154120 75120
rect 153620 75080 153626 75092
rect 154114 75080 154120 75092
rect 154172 75080 154178 75132
rect 169938 75080 169944 75132
rect 169996 75120 170002 75132
rect 170214 75120 170220 75132
rect 169996 75092 170220 75120
rect 169996 75080 170002 75092
rect 170214 75080 170220 75092
rect 170272 75080 170278 75132
rect 124030 75052 124036 75064
rect 118666 75024 124036 75052
rect 124030 75012 124036 75024
rect 124088 75012 124094 75064
rect 135438 75012 135444 75064
rect 135496 75052 135502 75064
rect 136174 75052 136180 75064
rect 135496 75024 136180 75052
rect 135496 75012 135502 75024
rect 136174 75012 136180 75024
rect 136232 75012 136238 75064
rect 156230 75012 156236 75064
rect 156288 75052 156294 75064
rect 156782 75052 156788 75064
rect 156288 75024 156788 75052
rect 156288 75012 156294 75024
rect 156782 75012 156788 75024
rect 156840 75012 156846 75064
rect 163222 75012 163228 75064
rect 163280 75052 163286 75064
rect 163682 75052 163688 75064
rect 163280 75024 163688 75052
rect 163280 75012 163286 75024
rect 163682 75012 163688 75024
rect 163740 75012 163746 75064
rect 156138 74944 156144 74996
rect 156196 74984 156202 74996
rect 156874 74984 156880 74996
rect 156196 74956 156880 74984
rect 156196 74944 156202 74956
rect 156874 74944 156880 74956
rect 156932 74944 156938 74996
rect 136726 74604 136732 74656
rect 136784 74644 136790 74656
rect 137002 74644 137008 74656
rect 136784 74616 137008 74644
rect 136784 74604 136790 74616
rect 137002 74604 137008 74616
rect 137060 74604 137066 74656
rect 139486 74604 139492 74656
rect 139544 74644 139550 74656
rect 140314 74644 140320 74656
rect 139544 74616 140320 74644
rect 139544 74604 139550 74616
rect 140314 74604 140320 74616
rect 140372 74604 140378 74656
rect 138474 74536 138480 74588
rect 138532 74576 138538 74588
rect 138750 74576 138756 74588
rect 138532 74548 138756 74576
rect 138532 74536 138538 74548
rect 138750 74536 138756 74548
rect 138808 74536 138814 74588
rect 144086 74536 144092 74588
rect 144144 74576 144150 74588
rect 144362 74576 144368 74588
rect 144144 74548 144368 74576
rect 144144 74536 144150 74548
rect 144362 74536 144368 74548
rect 144420 74536 144426 74588
rect 171226 74468 171232 74520
rect 171284 74508 171290 74520
rect 171686 74508 171692 74520
rect 171284 74480 171692 74508
rect 171284 74468 171290 74480
rect 171686 74468 171692 74480
rect 171744 74468 171750 74520
rect 149146 74400 149152 74452
rect 149204 74440 149210 74452
rect 150066 74440 150072 74452
rect 149204 74412 150072 74440
rect 149204 74400 149210 74412
rect 150066 74400 150072 74412
rect 150124 74400 150130 74452
rect 145466 74264 145472 74316
rect 145524 74304 145530 74316
rect 145742 74304 145748 74316
rect 145524 74276 145748 74304
rect 145524 74264 145530 74276
rect 145742 74264 145748 74276
rect 145800 74264 145806 74316
rect 141786 74128 141792 74180
rect 141844 74168 141850 74180
rect 209774 74168 209780 74180
rect 141844 74140 209780 74168
rect 141844 74128 141850 74140
rect 209774 74128 209780 74140
rect 209832 74128 209838 74180
rect 146294 74060 146300 74112
rect 146352 74100 146358 74112
rect 216674 74100 216680 74112
rect 146352 74072 216680 74100
rect 146352 74060 146358 74072
rect 216674 74060 216680 74072
rect 216732 74060 216738 74112
rect 119338 73992 119344 74044
rect 119396 74032 119402 74044
rect 130470 74032 130476 74044
rect 119396 74004 130476 74032
rect 119396 73992 119402 74004
rect 130470 73992 130476 74004
rect 130528 73992 130534 74044
rect 131114 73992 131120 74044
rect 131172 74032 131178 74044
rect 134978 74032 134984 74044
rect 131172 74004 134984 74032
rect 131172 73992 131178 74004
rect 134978 73992 134984 74004
rect 135036 73992 135042 74044
rect 143350 73992 143356 74044
rect 143408 74032 143414 74044
rect 223574 74032 223580 74044
rect 143408 74004 223580 74032
rect 143408 73992 143414 74004
rect 223574 73992 223580 74004
rect 223632 73992 223638 74044
rect 93946 73924 93952 73976
rect 94004 73964 94010 73976
rect 131022 73964 131028 73976
rect 94004 73936 131028 73964
rect 94004 73924 94010 73936
rect 131022 73924 131028 73936
rect 131080 73924 131086 73976
rect 147214 73924 147220 73976
rect 147272 73964 147278 73976
rect 251174 73964 251180 73976
rect 147272 73936 251180 73964
rect 147272 73924 147278 73936
rect 251174 73924 251180 73936
rect 251232 73924 251238 73976
rect 69106 73856 69112 73908
rect 69164 73896 69170 73908
rect 130838 73896 130844 73908
rect 69164 73868 130844 73896
rect 69164 73856 69170 73868
rect 130838 73856 130844 73868
rect 130896 73856 130902 73908
rect 137462 73856 137468 73908
rect 137520 73896 137526 73908
rect 139210 73896 139216 73908
rect 137520 73868 139216 73896
rect 137520 73856 137526 73868
rect 139210 73856 139216 73868
rect 139268 73856 139274 73908
rect 153286 73856 153292 73908
rect 153344 73896 153350 73908
rect 347774 73896 347780 73908
rect 153344 73868 347780 73896
rect 153344 73856 153350 73868
rect 347774 73856 347780 73868
rect 347832 73856 347838 73908
rect 30374 73788 30380 73840
rect 30432 73828 30438 73840
rect 127894 73828 127900 73840
rect 30432 73800 127900 73828
rect 30432 73788 30438 73800
rect 127894 73788 127900 73800
rect 127952 73788 127958 73840
rect 141326 73788 141332 73840
rect 141384 73828 141390 73840
rect 141602 73828 141608 73840
rect 141384 73800 141608 73828
rect 141384 73788 141390 73800
rect 141602 73788 141608 73800
rect 141660 73788 141666 73840
rect 157978 73788 157984 73840
rect 158036 73828 158042 73840
rect 390554 73828 390560 73840
rect 158036 73800 390560 73828
rect 158036 73788 158042 73800
rect 390554 73788 390560 73800
rect 390612 73788 390618 73840
rect 136726 73720 136732 73772
rect 136784 73760 136790 73772
rect 137554 73760 137560 73772
rect 136784 73732 137560 73760
rect 136784 73720 136790 73732
rect 137554 73720 137560 73732
rect 137612 73720 137618 73772
rect 138014 73244 138020 73296
rect 138072 73284 138078 73296
rect 142982 73284 142988 73296
rect 138072 73256 142988 73284
rect 138072 73244 138078 73256
rect 142982 73244 142988 73256
rect 143040 73244 143046 73296
rect 171042 73108 171048 73160
rect 171100 73148 171106 73160
rect 580166 73148 580172 73160
rect 171100 73120 580172 73148
rect 171100 73108 171106 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 150066 72768 150072 72820
rect 150124 72808 150130 72820
rect 307754 72808 307760 72820
rect 150124 72780 307760 72808
rect 150124 72768 150130 72780
rect 307754 72768 307760 72780
rect 307812 72768 307818 72820
rect 122282 72700 122288 72752
rect 122340 72740 122346 72752
rect 130562 72740 130568 72752
rect 122340 72712 130568 72740
rect 122340 72700 122346 72712
rect 130562 72700 130568 72712
rect 130620 72700 130626 72752
rect 149698 72700 149704 72752
rect 149756 72740 149762 72752
rect 311894 72740 311900 72752
rect 149756 72712 311900 72740
rect 149756 72700 149762 72712
rect 311894 72700 311900 72712
rect 311952 72700 311958 72752
rect 114554 72632 114560 72684
rect 114612 72672 114618 72684
rect 134518 72672 134524 72684
rect 114612 72644 134524 72672
rect 114612 72632 114618 72644
rect 134518 72632 134524 72644
rect 134576 72632 134582 72684
rect 151446 72632 151452 72684
rect 151504 72672 151510 72684
rect 325694 72672 325700 72684
rect 151504 72644 325700 72672
rect 151504 72632 151510 72644
rect 325694 72632 325700 72644
rect 325752 72632 325758 72684
rect 96614 72564 96620 72616
rect 96672 72604 96678 72616
rect 133138 72604 133144 72616
rect 96672 72576 133144 72604
rect 96672 72564 96678 72576
rect 133138 72564 133144 72576
rect 133196 72564 133202 72616
rect 151722 72564 151728 72616
rect 151780 72604 151786 72616
rect 332594 72604 332600 72616
rect 151780 72576 332600 72604
rect 151780 72564 151786 72576
rect 332594 72564 332600 72576
rect 332652 72564 332658 72616
rect 85574 72496 85580 72548
rect 85632 72536 85638 72548
rect 132310 72536 132316 72548
rect 85632 72508 132316 72536
rect 85632 72496 85638 72508
rect 132310 72496 132316 72508
rect 132368 72496 132374 72548
rect 154482 72496 154488 72548
rect 154540 72536 154546 72548
rect 340874 72536 340880 72548
rect 154540 72508 340880 72536
rect 154540 72496 154546 72508
rect 340874 72496 340880 72508
rect 340932 72496 340938 72548
rect 26234 72428 26240 72480
rect 26292 72468 26298 72480
rect 127802 72468 127808 72480
rect 26292 72440 127808 72468
rect 26292 72428 26298 72440
rect 127802 72428 127808 72440
rect 127860 72428 127866 72480
rect 152458 72428 152464 72480
rect 152516 72468 152522 72480
rect 343634 72468 343640 72480
rect 152516 72440 343640 72468
rect 152516 72428 152522 72440
rect 343634 72428 343640 72440
rect 343692 72428 343698 72480
rect 166626 72360 166632 72412
rect 166684 72400 166690 72412
rect 173250 72400 173256 72412
rect 166684 72372 173256 72400
rect 166684 72360 166690 72372
rect 173250 72360 173256 72372
rect 173308 72360 173314 72412
rect 132586 71680 132592 71732
rect 132644 71720 132650 71732
rect 135346 71720 135352 71732
rect 132644 71692 135352 71720
rect 132644 71680 132650 71692
rect 135346 71680 135352 71692
rect 135404 71680 135410 71732
rect 3418 71612 3424 71664
rect 3476 71652 3482 71664
rect 9030 71652 9036 71664
rect 3476 71624 9036 71652
rect 3476 71612 3482 71624
rect 9030 71612 9036 71624
rect 9088 71612 9094 71664
rect 121454 71408 121460 71460
rect 121512 71448 121518 71460
rect 134886 71448 134892 71460
rect 121512 71420 134892 71448
rect 121512 71408 121518 71420
rect 134886 71408 134892 71420
rect 134944 71408 134950 71460
rect 100754 71340 100760 71392
rect 100812 71380 100818 71392
rect 133690 71380 133696 71392
rect 100812 71352 133696 71380
rect 100812 71340 100818 71352
rect 133690 71340 133696 71352
rect 133748 71340 133754 71392
rect 82814 71272 82820 71324
rect 82872 71312 82878 71324
rect 131298 71312 131304 71324
rect 82872 71284 131304 71312
rect 82872 71272 82878 71284
rect 131298 71272 131304 71284
rect 131356 71272 131362 71324
rect 155310 71272 155316 71324
rect 155368 71312 155374 71324
rect 382274 71312 382280 71324
rect 155368 71284 382280 71312
rect 155368 71272 155374 71284
rect 382274 71272 382280 71284
rect 382332 71272 382338 71324
rect 48314 71204 48320 71256
rect 48372 71244 48378 71256
rect 129366 71244 129372 71256
rect 48372 71216 129372 71244
rect 48372 71204 48378 71216
rect 129366 71204 129372 71216
rect 129424 71204 129430 71256
rect 157886 71204 157892 71256
rect 157944 71244 157950 71256
rect 408494 71244 408500 71256
rect 157944 71216 408500 71244
rect 157944 71204 157950 71216
rect 408494 71204 408500 71216
rect 408552 71204 408558 71256
rect 28994 71136 29000 71188
rect 29052 71176 29058 71188
rect 128078 71176 128084 71188
rect 29052 71148 128084 71176
rect 29052 71136 29058 71148
rect 128078 71136 128084 71148
rect 128136 71136 128142 71188
rect 165246 71136 165252 71188
rect 165304 71176 165310 71188
rect 500954 71176 500960 71188
rect 165304 71148 500960 71176
rect 165304 71136 165310 71148
rect 500954 71136 500960 71148
rect 501012 71136 501018 71188
rect 16574 71068 16580 71120
rect 16632 71108 16638 71120
rect 126606 71108 126612 71120
rect 16632 71080 126612 71108
rect 16632 71068 16638 71080
rect 126606 71068 126612 71080
rect 126664 71068 126670 71120
rect 164878 71068 164884 71120
rect 164936 71108 164942 71120
rect 507854 71108 507860 71120
rect 164936 71080 507860 71108
rect 164936 71068 164942 71080
rect 507854 71068 507860 71080
rect 507912 71068 507918 71120
rect 11054 71000 11060 71052
rect 11112 71040 11118 71052
rect 126514 71040 126520 71052
rect 11112 71012 126520 71040
rect 11112 71000 11118 71012
rect 126514 71000 126520 71012
rect 126572 71000 126578 71052
rect 139302 71000 139308 71052
rect 139360 71040 139366 71052
rect 165062 71040 165068 71052
rect 139360 71012 165068 71040
rect 139360 71000 139366 71012
rect 165062 71000 165068 71012
rect 165120 71000 165126 71052
rect 166166 71000 166172 71052
rect 166224 71040 166230 71052
rect 523034 71040 523040 71052
rect 166224 71012 523040 71040
rect 166224 71000 166230 71012
rect 523034 71000 523040 71012
rect 523092 71000 523098 71052
rect 141510 69980 141516 70032
rect 141568 70020 141574 70032
rect 209866 70020 209872 70032
rect 141568 69992 209872 70020
rect 141568 69980 141574 69992
rect 209866 69980 209872 69992
rect 209924 69980 209930 70032
rect 159358 69912 159364 69964
rect 159416 69952 159422 69964
rect 431954 69952 431960 69964
rect 159416 69924 431960 69952
rect 159416 69912 159422 69924
rect 431954 69912 431960 69924
rect 432012 69912 432018 69964
rect 103514 69844 103520 69896
rect 103572 69884 103578 69896
rect 133046 69884 133052 69896
rect 103572 69856 133052 69884
rect 103572 69844 103578 69856
rect 133046 69844 133052 69856
rect 133104 69844 133110 69896
rect 159266 69844 159272 69896
rect 159324 69884 159330 69896
rect 437474 69884 437480 69896
rect 159324 69856 437480 69884
rect 159324 69844 159330 69856
rect 437474 69844 437480 69856
rect 437532 69844 437538 69896
rect 78674 69776 78680 69828
rect 78732 69816 78738 69828
rect 131850 69816 131856 69828
rect 78732 69788 131856 69816
rect 78732 69776 78738 69788
rect 131850 69776 131856 69788
rect 131908 69776 131914 69828
rect 160830 69776 160836 69828
rect 160888 69816 160894 69828
rect 447134 69816 447140 69828
rect 160888 69788 447140 69816
rect 160888 69776 160894 69788
rect 447134 69776 447140 69788
rect 447192 69776 447198 69828
rect 60734 69708 60740 69760
rect 60792 69748 60798 69760
rect 129090 69748 129096 69760
rect 60792 69720 129096 69748
rect 60792 69708 60798 69720
rect 129090 69708 129096 69720
rect 129148 69708 129154 69760
rect 167914 69708 167920 69760
rect 167972 69748 167978 69760
rect 536834 69748 536840 69760
rect 167972 69720 536840 69748
rect 167972 69708 167978 69720
rect 536834 69708 536840 69720
rect 536892 69708 536898 69760
rect 44174 69640 44180 69692
rect 44232 69680 44238 69692
rect 128906 69680 128912 69692
rect 44232 69652 128912 69680
rect 44232 69640 44238 69652
rect 128906 69640 128912 69652
rect 128964 69640 128970 69692
rect 169478 69640 169484 69692
rect 169536 69680 169542 69692
rect 564434 69680 564440 69692
rect 169536 69652 564440 69680
rect 169536 69640 169542 69652
rect 564434 69640 564440 69652
rect 564492 69640 564498 69692
rect 137278 68960 137284 69012
rect 137336 69000 137342 69012
rect 138750 69000 138756 69012
rect 137336 68972 138756 69000
rect 137336 68960 137342 68972
rect 138750 68960 138756 68972
rect 138808 68960 138814 69012
rect 138658 68892 138664 68944
rect 138716 68932 138722 68944
rect 140130 68932 140136 68944
rect 138716 68904 140136 68932
rect 138716 68892 138722 68904
rect 140130 68892 140136 68904
rect 140188 68892 140194 68944
rect 141418 68552 141424 68604
rect 141476 68592 141482 68604
rect 202874 68592 202880 68604
rect 141476 68564 202880 68592
rect 141476 68552 141482 68564
rect 202874 68552 202880 68564
rect 202932 68552 202938 68604
rect 144270 68484 144276 68536
rect 144328 68524 144334 68536
rect 238754 68524 238760 68536
rect 144328 68496 238760 68524
rect 144328 68484 144334 68496
rect 238754 68484 238760 68496
rect 238812 68484 238818 68536
rect 157150 68416 157156 68468
rect 157208 68456 157214 68468
rect 320174 68456 320180 68468
rect 157208 68428 320180 68456
rect 157208 68416 157214 68428
rect 320174 68416 320180 68428
rect 320232 68416 320238 68468
rect 162118 68348 162124 68400
rect 162176 68388 162182 68400
rect 467834 68388 467840 68400
rect 162176 68360 467840 68388
rect 162176 68348 162182 68360
rect 467834 68348 467840 68360
rect 467892 68348 467898 68400
rect 115934 68280 115940 68332
rect 115992 68320 115998 68332
rect 134242 68320 134248 68332
rect 115992 68292 134248 68320
rect 115992 68280 115998 68292
rect 134242 68280 134248 68292
rect 134300 68280 134306 68332
rect 169018 68280 169024 68332
rect 169076 68320 169082 68332
rect 561674 68320 561680 68332
rect 169076 68292 561680 68320
rect 169076 68280 169082 68292
rect 561674 68280 561680 68292
rect 561732 68280 561738 68332
rect 145558 67056 145564 67108
rect 145616 67096 145622 67108
rect 256694 67096 256700 67108
rect 145616 67068 256700 67096
rect 145616 67056 145622 67068
rect 256694 67056 256700 67068
rect 256752 67056 256758 67108
rect 156690 66988 156696 67040
rect 156748 67028 156754 67040
rect 396074 67028 396080 67040
rect 156748 67000 396080 67028
rect 156748 66988 156754 67000
rect 396074 66988 396080 67000
rect 396132 66988 396138 67040
rect 167730 66920 167736 66972
rect 167788 66960 167794 66972
rect 539594 66960 539600 66972
rect 167788 66932 539600 66960
rect 167788 66920 167794 66932
rect 539594 66920 539600 66932
rect 539652 66920 539658 66972
rect 33134 66852 33140 66904
rect 33192 66892 33198 66904
rect 127526 66892 127532 66904
rect 33192 66864 127532 66892
rect 33192 66852 33198 66864
rect 127526 66852 127532 66864
rect 127584 66852 127590 66904
rect 167638 66852 167644 66904
rect 167696 66892 167702 66904
rect 543734 66892 543740 66904
rect 167696 66864 543740 66892
rect 167696 66852 167702 66864
rect 543734 66852 543740 66864
rect 543792 66852 543798 66904
rect 138566 66172 138572 66224
rect 138624 66212 138630 66224
rect 140222 66212 140228 66224
rect 138624 66184 140228 66212
rect 138624 66172 138630 66184
rect 140222 66172 140228 66184
rect 140280 66172 140286 66224
rect 142706 65628 142712 65680
rect 142764 65668 142770 65680
rect 218054 65668 218060 65680
rect 142764 65640 218060 65668
rect 142764 65628 142770 65640
rect 218054 65628 218060 65640
rect 218112 65628 218118 65680
rect 144178 65560 144184 65612
rect 144236 65600 144242 65612
rect 234614 65600 234620 65612
rect 144236 65572 234620 65600
rect 144236 65560 144242 65572
rect 234614 65560 234620 65572
rect 234672 65560 234678 65612
rect 155770 65492 155776 65544
rect 155828 65532 155834 65544
rect 367094 65532 367100 65544
rect 155828 65504 367100 65532
rect 155828 65492 155834 65504
rect 367094 65492 367100 65504
rect 367152 65492 367158 65544
rect 141326 64404 141332 64456
rect 141384 64444 141390 64456
rect 207014 64444 207020 64456
rect 141384 64416 207020 64444
rect 141384 64404 141390 64416
rect 207014 64404 207020 64416
rect 207072 64404 207078 64456
rect 142614 64336 142620 64388
rect 142672 64376 142678 64388
rect 220814 64376 220820 64388
rect 142672 64348 220820 64376
rect 142672 64336 142678 64348
rect 220814 64336 220820 64348
rect 220872 64336 220878 64388
rect 153654 64268 153660 64320
rect 153712 64308 153718 64320
rect 362954 64308 362960 64320
rect 153712 64280 362960 64308
rect 153712 64268 153718 64280
rect 362954 64268 362960 64280
rect 363012 64268 363018 64320
rect 158346 64200 158352 64252
rect 158404 64240 158410 64252
rect 374086 64240 374092 64252
rect 158404 64212 374092 64240
rect 158404 64200 158410 64212
rect 374086 64200 374092 64212
rect 374144 64200 374150 64252
rect 155126 64132 155132 64184
rect 155184 64172 155190 64184
rect 376754 64172 376760 64184
rect 155184 64144 376760 64172
rect 155184 64132 155190 64144
rect 376754 64132 376760 64144
rect 376812 64132 376818 64184
rect 144086 62908 144092 62960
rect 144144 62948 144150 62960
rect 242894 62948 242900 62960
rect 144144 62920 242900 62948
rect 144144 62908 144150 62920
rect 242894 62908 242900 62920
rect 242952 62908 242958 62960
rect 151078 62840 151084 62892
rect 151136 62880 151142 62892
rect 324314 62880 324320 62892
rect 151136 62852 324320 62880
rect 151136 62840 151142 62852
rect 324314 62840 324320 62852
rect 324372 62840 324378 62892
rect 137186 62772 137192 62824
rect 137244 62812 137250 62824
rect 144178 62812 144184 62824
rect 137244 62784 144184 62812
rect 137244 62772 137250 62784
rect 144178 62772 144184 62784
rect 144236 62772 144242 62824
rect 163590 62772 163596 62824
rect 163648 62812 163654 62824
rect 481634 62812 481640 62824
rect 163648 62784 481640 62812
rect 163648 62772 163654 62784
rect 481634 62772 481640 62784
rect 481692 62772 481698 62824
rect 142522 61616 142528 61668
rect 142580 61656 142586 61668
rect 224954 61656 224960 61668
rect 142580 61628 224960 61656
rect 142580 61616 142586 61628
rect 224954 61616 224960 61628
rect 225012 61616 225018 61668
rect 162302 61548 162308 61600
rect 162360 61588 162366 61600
rect 368474 61588 368480 61600
rect 162360 61560 368480 61588
rect 162360 61548 162366 61560
rect 368474 61548 368480 61560
rect 368532 61548 368538 61600
rect 156598 61480 156604 61532
rect 156656 61520 156662 61532
rect 390646 61520 390652 61532
rect 156656 61492 390652 61520
rect 156656 61480 156662 61492
rect 390646 61480 390652 61492
rect 390704 61480 390710 61532
rect 157886 61412 157892 61464
rect 157944 61452 157950 61464
rect 412634 61452 412640 61464
rect 157944 61424 412640 61452
rect 157944 61412 157950 61424
rect 412634 61412 412640 61424
rect 412692 61412 412698 61464
rect 102134 61344 102140 61396
rect 102192 61384 102198 61396
rect 125410 61384 125416 61396
rect 102192 61356 125416 61384
rect 102192 61344 102198 61356
rect 125410 61344 125416 61356
rect 125468 61344 125474 61396
rect 159174 61344 159180 61396
rect 159232 61384 159238 61396
rect 440234 61384 440240 61396
rect 159232 61356 440240 61384
rect 159232 61344 159238 61356
rect 440234 61344 440240 61356
rect 440292 61344 440298 61396
rect 137094 60664 137100 60716
rect 137152 60704 137158 60716
rect 142798 60704 142804 60716
rect 137152 60676 142804 60704
rect 137152 60664 137158 60676
rect 142798 60664 142804 60676
rect 142856 60664 142862 60716
rect 183002 60664 183008 60716
rect 183060 60704 183066 60716
rect 580166 60704 580172 60716
rect 183060 60676 580172 60704
rect 183060 60664 183066 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 140038 60324 140044 60376
rect 140096 60364 140102 60376
rect 180794 60364 180800 60376
rect 140096 60336 180800 60364
rect 140096 60324 140102 60336
rect 180794 60324 180800 60336
rect 180852 60324 180858 60376
rect 120074 60256 120080 60308
rect 120132 60296 120138 60308
rect 123662 60296 123668 60308
rect 120132 60268 123668 60296
rect 120132 60256 120138 60268
rect 123662 60256 123668 60268
rect 123720 60256 123726 60308
rect 145466 60256 145472 60308
rect 145524 60296 145530 60308
rect 259454 60296 259460 60308
rect 145524 60268 259460 60296
rect 145524 60256 145530 60268
rect 259454 60256 259460 60268
rect 259512 60256 259518 60308
rect 150986 60188 150992 60240
rect 151044 60228 151050 60240
rect 327074 60228 327080 60240
rect 151044 60200 327080 60228
rect 151044 60188 151050 60200
rect 327074 60188 327080 60200
rect 327132 60188 327138 60240
rect 160738 60120 160744 60172
rect 160796 60160 160802 60172
rect 444374 60160 444380 60172
rect 160796 60132 444380 60160
rect 160796 60120 160802 60132
rect 444374 60120 444380 60132
rect 444432 60120 444438 60172
rect 163498 60052 163504 60104
rect 163556 60092 163562 60104
rect 481726 60092 481732 60104
rect 163556 60064 481732 60092
rect 163556 60052 163562 60064
rect 481726 60052 481732 60064
rect 481784 60052 481790 60104
rect 164786 59984 164792 60036
rect 164844 60024 164850 60036
rect 498286 60024 498292 60036
rect 164844 59996 498292 60024
rect 164844 59984 164850 59996
rect 498286 59984 498292 59996
rect 498344 59984 498350 60036
rect 3050 59304 3056 59356
rect 3108 59344 3114 59356
rect 181530 59344 181536 59356
rect 3108 59316 181536 59344
rect 3108 59304 3114 59316
rect 181530 59304 181536 59316
rect 181588 59304 181594 59356
rect 149606 58760 149612 58812
rect 149664 58800 149670 58812
rect 309134 58800 309140 58812
rect 149664 58772 309140 58800
rect 149664 58760 149670 58772
rect 309134 58760 309140 58772
rect 309192 58760 309198 58812
rect 152458 58692 152464 58744
rect 152516 58732 152522 58744
rect 340966 58732 340972 58744
rect 152516 58704 340972 58732
rect 152516 58692 152522 58704
rect 340966 58692 340972 58704
rect 341024 58692 341030 58744
rect 155034 58624 155040 58676
rect 155092 58664 155098 58676
rect 383654 58664 383660 58676
rect 155092 58636 383660 58664
rect 155092 58624 155098 58636
rect 383654 58624 383660 58636
rect 383712 58624 383718 58676
rect 137002 57876 137008 57928
rect 137060 57916 137066 57928
rect 140038 57916 140044 57928
rect 137060 57888 140044 57916
rect 137060 57876 137066 57888
rect 140038 57876 140044 57888
rect 140096 57876 140102 57928
rect 139946 57536 139952 57588
rect 140004 57576 140010 57588
rect 179414 57576 179420 57588
rect 140004 57548 179420 57576
rect 140004 57536 140010 57548
rect 179414 57536 179420 57548
rect 179472 57536 179478 57588
rect 152366 57468 152372 57520
rect 152424 57508 152430 57520
rect 345014 57508 345020 57520
rect 152424 57480 345020 57508
rect 152424 57468 152430 57480
rect 345014 57468 345020 57480
rect 345072 57468 345078 57520
rect 156506 57400 156512 57452
rect 156564 57440 156570 57452
rect 394694 57440 394700 57452
rect 156564 57412 394700 57440
rect 156564 57400 156570 57412
rect 394694 57400 394700 57412
rect 394752 57400 394758 57452
rect 159082 57332 159088 57384
rect 159140 57372 159146 57384
rect 433334 57372 433340 57384
rect 159140 57344 433340 57372
rect 159140 57332 159146 57344
rect 433334 57332 433340 57344
rect 433392 57332 433398 57384
rect 164694 57264 164700 57316
rect 164752 57304 164758 57316
rect 505094 57304 505100 57316
rect 164752 57276 505100 57304
rect 164752 57264 164758 57276
rect 505094 57264 505100 57276
rect 505152 57264 505158 57316
rect 95234 57196 95240 57248
rect 95292 57236 95298 57248
rect 125318 57236 125324 57248
rect 95292 57208 125324 57236
rect 95292 57196 95298 57208
rect 125318 57196 125324 57208
rect 125376 57196 125382 57248
rect 168926 57196 168932 57248
rect 168984 57236 168990 57248
rect 564526 57236 564532 57248
rect 168984 57208 564532 57236
rect 168984 57196 168990 57208
rect 564526 57196 564532 57208
rect 564584 57196 564590 57248
rect 153562 55904 153568 55956
rect 153620 55944 153626 55956
rect 365714 55944 365720 55956
rect 153620 55916 365720 55944
rect 153620 55904 153626 55916
rect 365714 55904 365720 55916
rect 365772 55904 365778 55956
rect 88334 55836 88340 55888
rect 88392 55876 88398 55888
rect 125226 55876 125232 55888
rect 88392 55848 125232 55876
rect 88392 55836 88398 55848
rect 125226 55836 125232 55848
rect 125284 55836 125290 55888
rect 157794 55836 157800 55888
rect 157852 55876 157858 55888
rect 415394 55876 415400 55888
rect 157852 55848 415400 55876
rect 157852 55836 157858 55848
rect 415394 55836 415400 55848
rect 415452 55836 415458 55888
rect 150894 54748 150900 54800
rect 150952 54788 150958 54800
rect 331214 54788 331220 54800
rect 150952 54760 331220 54788
rect 150952 54748 150958 54760
rect 331214 54748 331220 54760
rect 331272 54748 331278 54800
rect 154942 54680 154948 54732
rect 155000 54720 155006 54732
rect 380894 54720 380900 54732
rect 155000 54692 380900 54720
rect 155000 54680 155006 54692
rect 380894 54680 380900 54692
rect 380952 54680 380958 54732
rect 156414 54612 156420 54664
rect 156472 54652 156478 54664
rect 398834 54652 398840 54664
rect 156472 54624 398840 54652
rect 156472 54612 156478 54624
rect 398834 54612 398840 54624
rect 398892 54612 398898 54664
rect 160646 54544 160652 54596
rect 160704 54584 160710 54596
rect 448514 54584 448520 54596
rect 160704 54556 448520 54584
rect 160704 54544 160710 54556
rect 448514 54544 448520 54556
rect 448572 54544 448578 54596
rect 163406 54476 163412 54528
rect 163464 54516 163470 54528
rect 487154 54516 487160 54528
rect 163464 54488 487160 54516
rect 163464 54476 163470 54488
rect 487154 54476 487160 54488
rect 487212 54476 487218 54528
rect 157702 53320 157708 53372
rect 157760 53360 157766 53372
rect 419534 53360 419540 53372
rect 157760 53332 419540 53360
rect 157760 53320 157766 53332
rect 419534 53320 419540 53332
rect 419592 53320 419598 53372
rect 160554 53252 160560 53304
rect 160612 53292 160618 53304
rect 451274 53292 451280 53304
rect 160612 53264 451280 53292
rect 160612 53252 160618 53264
rect 451274 53252 451280 53264
rect 451332 53252 451338 53304
rect 167546 53184 167552 53236
rect 167604 53224 167610 53236
rect 538214 53224 538220 53236
rect 167604 53196 538220 53224
rect 167604 53184 167610 53196
rect 538214 53184 538220 53196
rect 538272 53184 538278 53236
rect 168834 53116 168840 53168
rect 168892 53156 168898 53168
rect 552014 53156 552020 53168
rect 168892 53128 552020 53156
rect 168892 53116 168898 53128
rect 552014 53116 552020 53128
rect 552072 53116 552078 53168
rect 170122 53048 170128 53100
rect 170180 53088 170186 53100
rect 571334 53088 571340 53100
rect 170180 53060 571340 53088
rect 170180 53048 170186 53060
rect 571334 53048 571340 53060
rect 571392 53048 571398 53100
rect 141234 51824 141240 51876
rect 141292 51864 141298 51876
rect 204254 51864 204260 51876
rect 141292 51836 204260 51864
rect 141292 51824 141298 51836
rect 204254 51824 204260 51836
rect 204312 51824 204318 51876
rect 166074 51756 166080 51808
rect 166132 51796 166138 51808
rect 527174 51796 527180 51808
rect 166132 51768 527180 51796
rect 166132 51756 166138 51768
rect 527174 51756 527180 51768
rect 527232 51756 527238 51808
rect 13814 51688 13820 51740
rect 13872 51728 13878 51740
rect 125134 51728 125140 51740
rect 13872 51700 125140 51728
rect 13872 51688 13878 51700
rect 125134 51688 125140 51700
rect 125192 51688 125198 51740
rect 138474 51688 138480 51740
rect 138532 51728 138538 51740
rect 166258 51728 166264 51740
rect 138532 51700 166264 51728
rect 138532 51688 138538 51700
rect 166258 51688 166264 51700
rect 166316 51688 166322 51740
rect 167454 51688 167460 51740
rect 167512 51728 167518 51740
rect 534074 51728 534080 51740
rect 167512 51700 534080 51728
rect 167512 51688 167518 51700
rect 534074 51688 534080 51700
rect 534132 51688 534138 51740
rect 143994 50600 144000 50652
rect 144052 50640 144058 50652
rect 233234 50640 233240 50652
rect 144052 50612 233240 50640
rect 144052 50600 144058 50612
rect 233234 50600 233240 50612
rect 233292 50600 233298 50652
rect 165982 50532 165988 50584
rect 166040 50572 166046 50584
rect 520274 50572 520280 50584
rect 166040 50544 520280 50572
rect 166040 50532 166046 50544
rect 520274 50532 520280 50544
rect 520332 50532 520338 50584
rect 165798 50464 165804 50516
rect 165856 50504 165862 50516
rect 523126 50504 523132 50516
rect 165856 50476 523132 50504
rect 165856 50464 165862 50476
rect 523126 50464 523132 50476
rect 523184 50464 523190 50516
rect 170766 50396 170772 50448
rect 170824 50436 170830 50448
rect 550634 50436 550640 50448
rect 170824 50408 550640 50436
rect 170824 50396 170830 50408
rect 550634 50396 550640 50408
rect 550692 50396 550698 50448
rect 170030 50328 170036 50380
rect 170088 50368 170094 50380
rect 569954 50368 569960 50380
rect 170088 50340 569960 50368
rect 170088 50328 170094 50340
rect 569954 50328 569960 50340
rect 570012 50328 570018 50380
rect 139854 49240 139860 49292
rect 139912 49280 139918 49292
rect 183554 49280 183560 49292
rect 139912 49252 183560 49280
rect 139912 49240 139918 49252
rect 183554 49240 183560 49252
rect 183612 49240 183618 49292
rect 153470 49172 153476 49224
rect 153528 49212 153534 49224
rect 357434 49212 357440 49224
rect 153528 49184 357440 49212
rect 153528 49172 153534 49184
rect 357434 49172 357440 49184
rect 357492 49172 357498 49224
rect 159726 49104 159732 49156
rect 159784 49144 159790 49156
rect 382366 49144 382372 49156
rect 159784 49116 382372 49144
rect 159784 49104 159790 49116
rect 382366 49104 382372 49116
rect 382424 49104 382430 49156
rect 171594 49036 171600 49088
rect 171652 49076 171658 49088
rect 432046 49076 432052 49088
rect 171652 49048 432052 49076
rect 171652 49036 171658 49048
rect 432046 49036 432052 49048
rect 432104 49036 432110 49088
rect 138382 48968 138388 49020
rect 138440 49008 138446 49020
rect 165798 49008 165804 49020
rect 138440 48980 165804 49008
rect 138440 48968 138446 48980
rect 165798 48968 165804 48980
rect 165856 48968 165862 49020
rect 165890 48968 165896 49020
rect 165948 49008 165954 49020
rect 516134 49008 516140 49020
rect 165948 48980 516140 49008
rect 165948 48968 165954 48980
rect 516134 48968 516140 48980
rect 516192 48968 516198 49020
rect 142430 47676 142436 47728
rect 142488 47716 142494 47728
rect 215294 47716 215300 47728
rect 142488 47688 215300 47716
rect 142488 47676 142494 47688
rect 215294 47676 215300 47688
rect 215352 47676 215358 47728
rect 164602 47608 164608 47660
rect 164660 47648 164666 47660
rect 502334 47648 502340 47660
rect 164660 47620 502340 47648
rect 164660 47608 164666 47620
rect 502334 47608 502340 47620
rect 502392 47608 502398 47660
rect 168650 47540 168656 47592
rect 168708 47580 168714 47592
rect 563054 47580 563060 47592
rect 168708 47552 563060 47580
rect 168708 47540 168714 47552
rect 563054 47540 563060 47552
rect 563112 47540 563118 47592
rect 118510 46860 118516 46912
rect 118568 46900 118574 46912
rect 580166 46900 580172 46912
rect 118568 46872 580172 46900
rect 118568 46860 118574 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 139762 46316 139768 46368
rect 139820 46356 139826 46368
rect 187694 46356 187700 46368
rect 139820 46328 187700 46356
rect 139820 46316 139826 46328
rect 187694 46316 187700 46328
rect 187752 46316 187758 46368
rect 143902 46248 143908 46300
rect 143960 46288 143966 46300
rect 235994 46288 236000 46300
rect 143960 46260 236000 46288
rect 143960 46248 143966 46260
rect 235994 46248 236000 46260
rect 236052 46248 236058 46300
rect 158990 46180 158996 46232
rect 159048 46220 159054 46232
rect 427814 46220 427820 46232
rect 159048 46192 427820 46220
rect 159048 46180 159054 46192
rect 427814 46180 427820 46192
rect 427872 46180 427878 46232
rect 3418 45500 3424 45552
rect 3476 45540 3482 45552
rect 173986 45540 173992 45552
rect 3476 45512 173992 45540
rect 3476 45500 3482 45512
rect 173986 45500 173992 45512
rect 174044 45500 174050 45552
rect 141142 45024 141148 45076
rect 141200 45064 141206 45076
rect 208394 45064 208400 45076
rect 141200 45036 208400 45064
rect 141200 45024 141206 45036
rect 208394 45024 208400 45036
rect 208452 45024 208458 45076
rect 152274 44956 152280 45008
rect 152332 44996 152338 45008
rect 339494 44996 339500 45008
rect 152332 44968 339500 44996
rect 152332 44956 152338 44968
rect 339494 44956 339500 44968
rect 339552 44956 339558 45008
rect 138290 44888 138296 44940
rect 138348 44928 138354 44940
rect 168650 44928 168656 44940
rect 138348 44900 168656 44928
rect 138348 44888 138354 44900
rect 168650 44888 168656 44900
rect 168708 44888 168714 44940
rect 171686 44888 171692 44940
rect 171744 44928 171750 44940
rect 425054 44928 425060 44940
rect 171744 44900 425060 44928
rect 171744 44888 171750 44900
rect 425054 44888 425060 44900
rect 425112 44888 425118 44940
rect 81434 44820 81440 44872
rect 81492 44860 81498 44872
rect 131574 44860 131580 44872
rect 81492 44832 131580 44860
rect 81492 44820 81498 44832
rect 131574 44820 131580 44832
rect 131632 44820 131638 44872
rect 163314 44820 163320 44872
rect 163372 44860 163378 44872
rect 485774 44860 485780 44872
rect 163372 44832 485780 44860
rect 163372 44820 163378 44832
rect 485774 44820 485780 44832
rect 485832 44820 485838 44872
rect 139670 43528 139676 43580
rect 139728 43568 139734 43580
rect 185026 43568 185032 43580
rect 139728 43540 185032 43568
rect 139728 43528 139734 43540
rect 185026 43528 185032 43540
rect 185084 43528 185090 43580
rect 152182 43460 152188 43512
rect 152240 43500 152246 43512
rect 349154 43500 349160 43512
rect 152240 43472 349160 43500
rect 152240 43460 152246 43472
rect 349154 43460 349160 43472
rect 349212 43460 349218 43512
rect 168742 43392 168748 43444
rect 168800 43432 168806 43444
rect 556154 43432 556160 43444
rect 168800 43404 556160 43432
rect 168800 43392 168806 43404
rect 556154 43392 556160 43404
rect 556212 43392 556218 43444
rect 142338 42168 142344 42220
rect 142396 42208 142402 42220
rect 218146 42208 218152 42220
rect 142396 42180 218152 42208
rect 142396 42168 142402 42180
rect 218146 42168 218152 42180
rect 218204 42168 218210 42220
rect 148318 42100 148324 42152
rect 148376 42140 148382 42152
rect 285674 42140 285680 42152
rect 148376 42112 285680 42140
rect 148376 42100 148382 42112
rect 285674 42100 285680 42112
rect 285732 42100 285738 42152
rect 150802 42032 150808 42084
rect 150860 42072 150866 42084
rect 328454 42072 328460 42084
rect 150860 42044 328460 42072
rect 150860 42032 150866 42044
rect 328454 42032 328460 42044
rect 328512 42032 328518 42084
rect 145374 37952 145380 38004
rect 145432 37992 145438 38004
rect 258074 37992 258080 38004
rect 145432 37964 258080 37992
rect 145432 37952 145438 37964
rect 258074 37952 258080 37964
rect 258132 37952 258138 38004
rect 45554 37884 45560 37936
rect 45612 37924 45618 37936
rect 116578 37924 116584 37936
rect 45612 37896 116584 37924
rect 45612 37884 45618 37896
rect 116578 37884 116584 37896
rect 116636 37884 116642 37936
rect 152090 37884 152096 37936
rect 152148 37924 152154 37936
rect 338114 37924 338120 37936
rect 152148 37896 338120 37924
rect 152148 37884 152154 37896
rect 338114 37884 338120 37896
rect 338172 37884 338178 37936
rect 7558 36524 7564 36576
rect 7616 36564 7622 36576
rect 124214 36564 124220 36576
rect 7616 36536 124220 36564
rect 7616 36524 7622 36536
rect 124214 36524 124220 36536
rect 124272 36524 124278 36576
rect 166626 36524 166632 36576
rect 166684 36564 166690 36576
rect 418154 36564 418160 36576
rect 166684 36536 418160 36564
rect 166684 36524 166690 36536
rect 418154 36524 418160 36536
rect 418212 36524 418218 36576
rect 148226 35368 148232 35420
rect 148284 35408 148290 35420
rect 291194 35408 291200 35420
rect 148284 35380 291200 35408
rect 148284 35368 148290 35380
rect 291194 35368 291200 35380
rect 291252 35368 291258 35420
rect 149514 35300 149520 35352
rect 149572 35340 149578 35352
rect 304994 35340 305000 35352
rect 149572 35312 305000 35340
rect 149572 35300 149578 35312
rect 304994 35300 305000 35312
rect 305052 35300 305058 35352
rect 160922 35232 160928 35284
rect 160980 35272 160986 35284
rect 375374 35272 375380 35284
rect 160980 35244 375380 35272
rect 160980 35232 160986 35244
rect 375374 35232 375380 35244
rect 375432 35232 375438 35284
rect 38654 35164 38660 35216
rect 38712 35204 38718 35216
rect 122374 35204 122380 35216
rect 38712 35176 122380 35204
rect 38712 35164 38718 35176
rect 122374 35164 122380 35176
rect 122432 35164 122438 35216
rect 163222 35164 163228 35216
rect 163280 35204 163286 35216
rect 490006 35204 490012 35216
rect 163280 35176 490012 35204
rect 163280 35164 163286 35176
rect 490006 35164 490012 35176
rect 490064 35164 490070 35216
rect 145282 33940 145288 33992
rect 145340 33980 145346 33992
rect 259546 33980 259552 33992
rect 145340 33952 259552 33980
rect 145340 33940 145346 33952
rect 259546 33940 259552 33952
rect 259604 33940 259610 33992
rect 148134 33872 148140 33924
rect 148192 33912 148198 33924
rect 287054 33912 287060 33924
rect 148192 33884 287060 33912
rect 148192 33872 148198 33884
rect 287054 33872 287060 33884
rect 287112 33872 287118 33924
rect 158898 33804 158904 33856
rect 158956 33844 158962 33856
rect 429194 33844 429200 33856
rect 158956 33816 429200 33844
rect 158956 33804 158962 33816
rect 429194 33804 429200 33816
rect 429252 33804 429258 33856
rect 169938 33736 169944 33788
rect 169996 33776 170002 33788
rect 572714 33776 572720 33788
rect 169996 33748 572720 33776
rect 169996 33736 170002 33748
rect 572714 33736 572720 33748
rect 572772 33736 572778 33788
rect 3142 33056 3148 33108
rect 3200 33096 3206 33108
rect 7650 33096 7656 33108
rect 3200 33068 7656 33096
rect 3200 33056 3206 33068
rect 7650 33056 7656 33068
rect 7708 33056 7714 33108
rect 173342 33056 173348 33108
rect 173400 33096 173406 33108
rect 580166 33096 580172 33108
rect 173400 33068 580172 33096
rect 173400 33056 173406 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 31754 32376 31760 32428
rect 31812 32416 31818 32428
rect 120810 32416 120816 32428
rect 31812 32388 120816 32416
rect 31812 32376 31818 32388
rect 120810 32376 120816 32388
rect 120868 32376 120874 32428
rect 142246 32376 142252 32428
rect 142304 32416 142310 32428
rect 219434 32416 219440 32428
rect 142304 32388 219440 32416
rect 142304 32376 142310 32388
rect 219434 32376 219440 32388
rect 219492 32376 219498 32428
rect 154114 31152 154120 31204
rect 154172 31192 154178 31204
rect 332686 31192 332692 31204
rect 154172 31164 332692 31192
rect 154172 31152 154178 31164
rect 332686 31152 332692 31164
rect 332744 31152 332750 31204
rect 150710 31084 150716 31136
rect 150768 31124 150774 31136
rect 329834 31124 329840 31136
rect 150768 31096 329840 31124
rect 150768 31084 150774 31096
rect 329834 31084 329840 31096
rect 329892 31084 329898 31136
rect 167362 31016 167368 31068
rect 167420 31056 167426 31068
rect 542354 31056 542360 31068
rect 167420 31028 542360 31056
rect 167420 31016 167426 31028
rect 542354 31016 542360 31028
rect 542412 31016 542418 31068
rect 145098 29928 145104 29980
rect 145156 29968 145162 29980
rect 251266 29968 251272 29980
rect 145156 29940 251272 29968
rect 145156 29928 145162 29940
rect 251266 29928 251272 29940
rect 251324 29928 251330 29980
rect 145190 29860 145196 29912
rect 145248 29900 145254 29912
rect 253934 29900 253940 29912
rect 145248 29872 253940 29900
rect 145248 29860 145254 29872
rect 253934 29860 253940 29872
rect 253992 29860 253998 29912
rect 150618 29792 150624 29844
rect 150676 29832 150682 29844
rect 324406 29832 324412 29844
rect 150676 29804 324412 29832
rect 150676 29792 150682 29804
rect 324406 29792 324412 29804
rect 324464 29792 324470 29844
rect 156322 29724 156328 29776
rect 156380 29764 156386 29776
rect 391934 29764 391940 29776
rect 156380 29736 391940 29764
rect 156380 29724 156386 29736
rect 391934 29724 391940 29736
rect 391992 29724 391998 29776
rect 160002 29656 160008 29708
rect 160060 29696 160066 29708
rect 434714 29696 434720 29708
rect 160060 29668 434720 29696
rect 160060 29656 160066 29668
rect 434714 29656 434720 29668
rect 434772 29656 434778 29708
rect 167270 29588 167276 29640
rect 167328 29628 167334 29640
rect 535454 29628 535460 29640
rect 167328 29600 535460 29628
rect 167328 29588 167334 29600
rect 535454 29588 535460 29600
rect 535512 29588 535518 29640
rect 141050 28500 141056 28552
rect 141108 28540 141114 28552
rect 201494 28540 201500 28552
rect 141108 28512 201500 28540
rect 141108 28500 141114 28512
rect 201494 28500 201500 28512
rect 201552 28500 201558 28552
rect 143810 28432 143816 28484
rect 143868 28472 143874 28484
rect 242986 28472 242992 28484
rect 143868 28444 242992 28472
rect 143868 28432 143874 28444
rect 242986 28432 242992 28444
rect 243044 28432 243050 28484
rect 151998 28364 152004 28416
rect 152056 28404 152062 28416
rect 346394 28404 346400 28416
rect 152056 28376 346400 28404
rect 152056 28364 152062 28376
rect 346394 28364 346400 28376
rect 346452 28364 346458 28416
rect 154850 28296 154856 28348
rect 154908 28336 154914 28348
rect 378134 28336 378140 28348
rect 154908 28308 378140 28336
rect 154908 28296 154914 28308
rect 378134 28296 378140 28308
rect 378192 28296 378198 28348
rect 171410 28228 171416 28280
rect 171468 28268 171474 28280
rect 397454 28268 397460 28280
rect 171468 28240 397460 28268
rect 171468 28228 171474 28240
rect 397454 28228 397460 28240
rect 397512 28228 397518 28280
rect 139578 27072 139584 27124
rect 139636 27112 139642 27124
rect 186314 27112 186320 27124
rect 139636 27084 186320 27112
rect 139636 27072 139642 27084
rect 186314 27072 186320 27084
rect 186372 27072 186378 27124
rect 171502 27004 171508 27056
rect 171560 27044 171566 27056
rect 411254 27044 411260 27056
rect 171560 27016 411260 27044
rect 171560 27004 171566 27016
rect 411254 27004 411260 27016
rect 411312 27004 411318 27056
rect 156230 26936 156236 26988
rect 156288 26976 156294 26988
rect 398926 26976 398932 26988
rect 156288 26948 398932 26976
rect 156288 26936 156294 26948
rect 398926 26936 398932 26948
rect 398984 26936 398990 26988
rect 165706 26868 165712 26920
rect 165764 26908 165770 26920
rect 524414 26908 524420 26920
rect 165764 26880 524420 26908
rect 165764 26868 165770 26880
rect 524414 26868 524420 26880
rect 524472 26868 524478 26920
rect 140958 25848 140964 25900
rect 141016 25888 141022 25900
rect 201586 25888 201592 25900
rect 141016 25860 201592 25888
rect 141016 25848 141022 25860
rect 201586 25848 201592 25860
rect 201644 25848 201650 25900
rect 149422 25780 149428 25832
rect 149480 25820 149486 25832
rect 303614 25820 303620 25832
rect 149480 25792 303620 25820
rect 149480 25780 149486 25792
rect 303614 25780 303620 25792
rect 303672 25780 303678 25832
rect 156138 25712 156144 25764
rect 156196 25752 156202 25764
rect 401594 25752 401600 25764
rect 156196 25724 401600 25752
rect 156196 25712 156202 25724
rect 401594 25712 401600 25724
rect 401652 25712 401658 25764
rect 157610 25644 157616 25696
rect 157668 25684 157674 25696
rect 414014 25684 414020 25696
rect 157668 25656 414020 25684
rect 157668 25644 157674 25656
rect 414014 25644 414020 25656
rect 414072 25644 414078 25696
rect 167178 25576 167184 25628
rect 167236 25616 167242 25628
rect 540974 25616 540980 25628
rect 167236 25588 540980 25616
rect 167236 25576 167242 25588
rect 540974 25576 540980 25588
rect 541032 25576 541038 25628
rect 167086 25508 167092 25560
rect 167144 25548 167150 25560
rect 545114 25548 545120 25560
rect 167144 25520 545120 25548
rect 167144 25508 167150 25520
rect 545114 25508 545120 25520
rect 545172 25508 545178 25560
rect 135806 24964 135812 25016
rect 135864 25004 135870 25016
rect 140958 25004 140964 25016
rect 135864 24976 140964 25004
rect 135864 24964 135870 24976
rect 140958 24964 140964 24976
rect 141016 24964 141022 25016
rect 140866 24352 140872 24404
rect 140924 24392 140930 24404
rect 198734 24392 198740 24404
rect 140924 24364 198740 24392
rect 140924 24352 140930 24364
rect 198734 24352 198740 24364
rect 198792 24352 198798 24404
rect 148042 24284 148048 24336
rect 148100 24324 148106 24336
rect 292666 24324 292672 24336
rect 148100 24296 292672 24324
rect 148100 24284 148106 24296
rect 292666 24284 292672 24296
rect 292724 24284 292730 24336
rect 97994 24216 98000 24268
rect 98052 24256 98058 24268
rect 132862 24256 132868 24268
rect 98052 24228 132868 24256
rect 98052 24216 98058 24228
rect 132862 24216 132868 24228
rect 132920 24216 132926 24268
rect 149330 24216 149336 24268
rect 149388 24256 149394 24268
rect 313274 24256 313280 24268
rect 149388 24228 313280 24256
rect 149388 24216 149394 24228
rect 313274 24216 313280 24228
rect 313332 24216 313338 24268
rect 27614 24148 27620 24200
rect 27672 24188 27678 24200
rect 127434 24188 127440 24200
rect 27672 24160 127440 24188
rect 27672 24148 27678 24160
rect 127434 24148 127440 24160
rect 127492 24148 127498 24200
rect 157518 24148 157524 24200
rect 157576 24188 157582 24200
rect 416774 24188 416780 24200
rect 157576 24160 416780 24188
rect 157576 24148 157582 24160
rect 416774 24148 416780 24160
rect 416832 24148 416838 24200
rect 3326 24080 3332 24132
rect 3384 24120 3390 24132
rect 179874 24120 179880 24132
rect 3384 24092 179880 24120
rect 3384 24080 3390 24092
rect 179874 24080 179880 24092
rect 179932 24080 179938 24132
rect 182818 24080 182824 24132
rect 182876 24120 182882 24132
rect 579614 24120 579620 24132
rect 182876 24092 579620 24120
rect 182876 24080 182882 24092
rect 579614 24080 579620 24092
rect 579672 24080 579678 24132
rect 135714 23876 135720 23928
rect 135772 23916 135778 23928
rect 139578 23916 139584 23928
rect 135772 23888 139584 23916
rect 135772 23876 135778 23888
rect 139578 23876 139584 23888
rect 139636 23876 139642 23928
rect 3418 23060 3424 23112
rect 3476 23100 3482 23112
rect 174078 23100 174084 23112
rect 3476 23072 174084 23100
rect 3476 23060 3482 23072
rect 174078 23060 174084 23072
rect 174136 23060 174142 23112
rect 172054 22992 172060 23044
rect 172112 23032 172118 23044
rect 404354 23032 404360 23044
rect 172112 23004 404360 23032
rect 172112 22992 172118 23004
rect 404354 22992 404360 23004
rect 404412 22992 404418 23044
rect 42794 22924 42800 22976
rect 42852 22964 42858 22976
rect 128630 22964 128636 22976
rect 42852 22936 128636 22964
rect 42852 22924 42858 22936
rect 128630 22924 128636 22936
rect 128688 22924 128694 22976
rect 157426 22924 157432 22976
rect 157484 22964 157490 22976
rect 409874 22964 409880 22976
rect 157484 22936 409880 22964
rect 157484 22924 157490 22936
rect 409874 22924 409880 22936
rect 409932 22924 409938 22976
rect 11146 22856 11152 22908
rect 11204 22896 11210 22908
rect 125962 22896 125968 22908
rect 11204 22868 125968 22896
rect 11204 22856 11210 22868
rect 125962 22856 125968 22868
rect 126020 22856 126026 22908
rect 160462 22856 160468 22908
rect 160520 22896 160526 22908
rect 455414 22896 455420 22908
rect 160520 22868 455420 22896
rect 160520 22856 160526 22868
rect 455414 22856 455420 22868
rect 455472 22856 455478 22908
rect 9674 22788 9680 22840
rect 9732 22828 9738 22840
rect 126054 22828 126060 22840
rect 9732 22800 126060 22828
rect 9732 22788 9738 22800
rect 126054 22788 126060 22800
rect 126112 22788 126118 22840
rect 136910 22788 136916 22840
rect 136968 22828 136974 22840
rect 148042 22828 148048 22840
rect 136968 22800 148048 22828
rect 136968 22788 136974 22800
rect 148042 22788 148048 22800
rect 148100 22788 148106 22840
rect 164510 22788 164516 22840
rect 164568 22828 164574 22840
rect 499574 22828 499580 22840
rect 164568 22800 499580 22828
rect 164568 22788 164574 22800
rect 499574 22788 499580 22800
rect 499632 22788 499638 22840
rect 118326 22720 118332 22772
rect 118384 22760 118390 22772
rect 580258 22760 580264 22772
rect 118384 22732 580264 22760
rect 118384 22720 118390 22732
rect 580258 22720 580264 22732
rect 580316 22720 580322 22772
rect 138842 22040 138848 22092
rect 138900 22080 138906 22092
rect 143810 22080 143816 22092
rect 138900 22052 143816 22080
rect 138900 22040 138906 22052
rect 143810 22040 143816 22052
rect 143868 22040 143874 22092
rect 160370 21428 160376 21480
rect 160428 21468 160434 21480
rect 454034 21468 454040 21480
rect 160428 21440 454040 21468
rect 160428 21428 160434 21440
rect 454034 21428 454040 21440
rect 454092 21428 454098 21480
rect 170490 21360 170496 21412
rect 170548 21400 170554 21412
rect 514846 21400 514852 21412
rect 170548 21372 514852 21400
rect 170548 21360 170554 21372
rect 514846 21360 514852 21372
rect 514904 21360 514910 21412
rect 144914 20136 144920 20188
rect 144972 20176 144978 20188
rect 262214 20176 262220 20188
rect 144972 20148 262220 20176
rect 144972 20136 144978 20148
rect 262214 20136 262220 20148
rect 262272 20136 262278 20188
rect 145006 20068 145012 20120
rect 145064 20108 145070 20120
rect 255314 20108 255320 20120
rect 145064 20080 255320 20108
rect 145064 20068 145070 20080
rect 255314 20068 255320 20080
rect 255372 20068 255378 20120
rect 255958 20068 255964 20120
rect 256016 20108 256022 20120
rect 456886 20108 456892 20120
rect 256016 20080 456892 20108
rect 256016 20068 256022 20080
rect 456886 20068 456892 20080
rect 456944 20068 456950 20120
rect 124214 20000 124220 20052
rect 124272 20040 124278 20052
rect 134150 20040 134156 20052
rect 124272 20012 134156 20040
rect 124272 20000 124278 20012
rect 134150 20000 134156 20012
rect 134208 20000 134214 20052
rect 143718 20000 143724 20052
rect 143776 20040 143782 20052
rect 241514 20040 241520 20052
rect 143776 20012 241520 20040
rect 143776 20000 143782 20012
rect 241514 20000 241520 20012
rect 241572 20000 241578 20052
rect 242158 20000 242164 20052
rect 242216 20040 242222 20052
rect 449894 20040 449900 20052
rect 242216 20012 449900 20040
rect 242216 20000 242222 20012
rect 449894 20000 449900 20012
rect 449952 20000 449958 20052
rect 67634 19932 67640 19984
rect 67692 19972 67698 19984
rect 130010 19972 130016 19984
rect 67692 19944 130016 19972
rect 67692 19932 67698 19944
rect 130010 19932 130016 19944
rect 130068 19932 130074 19984
rect 157334 19932 157340 19984
rect 157392 19972 157398 19984
rect 415486 19972 415492 19984
rect 157392 19944 415492 19972
rect 157392 19932 157398 19944
rect 415486 19932 415492 19944
rect 415544 19932 415550 19984
rect 143626 18844 143632 18896
rect 143684 18884 143690 18896
rect 234706 18884 234712 18896
rect 143684 18856 234712 18884
rect 143684 18844 143690 18856
rect 234706 18844 234712 18856
rect 234764 18844 234770 18896
rect 164418 18776 164424 18828
rect 164476 18816 164482 18828
rect 509234 18816 509240 18828
rect 164476 18788 509240 18816
rect 164476 18776 164482 18788
rect 509234 18776 509240 18788
rect 509292 18776 509298 18828
rect 168558 18708 168564 18760
rect 168616 18748 168622 18760
rect 553394 18748 553400 18760
rect 168616 18720 553400 18748
rect 168616 18708 168622 18720
rect 553394 18708 553400 18720
rect 553452 18708 553458 18760
rect 168466 18640 168472 18692
rect 168524 18680 168530 18692
rect 556246 18680 556252 18692
rect 168524 18652 556252 18680
rect 168524 18640 168530 18652
rect 556246 18640 556252 18652
rect 556304 18640 556310 18692
rect 168374 18572 168380 18624
rect 168432 18612 168438 18624
rect 560294 18612 560300 18624
rect 168432 18584 560300 18612
rect 168432 18572 168438 18584
rect 560294 18572 560300 18584
rect 560352 18572 560358 18624
rect 160278 17348 160284 17400
rect 160336 17388 160342 17400
rect 445754 17388 445760 17400
rect 160336 17360 445760 17388
rect 160336 17348 160342 17360
rect 445754 17348 445760 17360
rect 445812 17348 445818 17400
rect 160186 17280 160192 17332
rect 160244 17320 160250 17332
rect 448606 17320 448612 17332
rect 160244 17292 448612 17320
rect 160244 17280 160250 17292
rect 448606 17280 448612 17292
rect 448664 17280 448670 17332
rect 164326 17212 164332 17264
rect 164384 17252 164390 17264
rect 506566 17252 506572 17264
rect 164384 17224 506572 17252
rect 164384 17212 164390 17224
rect 506566 17212 506572 17224
rect 506624 17212 506630 17264
rect 144546 16056 144552 16108
rect 144604 16096 144610 16108
rect 237650 16096 237656 16108
rect 144604 16068 237656 16096
rect 144604 16056 144610 16068
rect 237650 16056 237656 16068
rect 237708 16056 237714 16108
rect 151906 15988 151912 16040
rect 151964 16028 151970 16040
rect 342898 16028 342904 16040
rect 151964 16000 342904 16028
rect 151964 15988 151970 16000
rect 342898 15988 342904 16000
rect 342956 15988 342962 16040
rect 153378 15920 153384 15972
rect 153436 15960 153442 15972
rect 361114 15960 361120 15972
rect 153436 15932 361120 15960
rect 153436 15920 153442 15932
rect 361114 15920 361120 15932
rect 361172 15920 361178 15972
rect 163130 15852 163136 15904
rect 163188 15892 163194 15904
rect 492306 15892 492312 15904
rect 163188 15864 492312 15892
rect 163188 15852 163194 15864
rect 492306 15852 492312 15864
rect 492364 15852 492370 15904
rect 147950 14696 147956 14748
rect 148008 14736 148014 14748
rect 289814 14736 289820 14748
rect 148008 14708 289820 14736
rect 148008 14696 148014 14708
rect 289814 14696 289820 14708
rect 289872 14696 289878 14748
rect 149238 14628 149244 14680
rect 149296 14668 149302 14680
rect 311434 14668 311440 14680
rect 149296 14640 311440 14668
rect 149296 14628 149302 14640
rect 311434 14628 311440 14640
rect 311492 14628 311498 14680
rect 154758 14560 154764 14612
rect 154816 14600 154822 14612
rect 386690 14600 386696 14612
rect 154816 14572 386696 14600
rect 154816 14560 154822 14572
rect 386690 14560 386696 14572
rect 386748 14560 386754 14612
rect 160094 14492 160100 14544
rect 160152 14532 160158 14544
rect 453298 14532 453304 14544
rect 160152 14504 453304 14532
rect 160152 14492 160158 14504
rect 453298 14492 453304 14504
rect 453356 14492 453362 14544
rect 163038 14424 163044 14476
rect 163096 14464 163102 14476
rect 488810 14464 488816 14476
rect 163096 14436 488816 14464
rect 163096 14424 163102 14436
rect 488810 14424 488816 14436
rect 488868 14424 488874 14476
rect 151814 13200 151820 13252
rect 151872 13240 151878 13252
rect 349246 13240 349252 13252
rect 151872 13212 349252 13240
rect 151872 13200 151878 13212
rect 349246 13200 349252 13212
rect 349304 13200 349310 13252
rect 155678 13132 155684 13184
rect 155736 13172 155742 13184
rect 361850 13172 361856 13184
rect 155736 13144 361856 13172
rect 155736 13132 155742 13144
rect 361850 13132 361856 13144
rect 361908 13132 361914 13184
rect 162946 13064 162952 13116
rect 163004 13104 163010 13116
rect 484762 13104 484768 13116
rect 163004 13076 484768 13104
rect 163004 13064 163010 13076
rect 484762 13064 484768 13076
rect 484820 13064 484826 13116
rect 106458 11772 106464 11824
rect 106516 11812 106522 11824
rect 132770 11812 132776 11824
rect 106516 11784 132776 11812
rect 106516 11772 106522 11784
rect 132770 11772 132776 11784
rect 132828 11772 132834 11824
rect 136818 11772 136824 11824
rect 136876 11812 136882 11824
rect 145466 11812 145472 11824
rect 136876 11784 145472 11812
rect 136876 11772 136882 11784
rect 145466 11772 145472 11784
rect 145524 11772 145530 11824
rect 156046 11772 156052 11824
rect 156104 11812 156110 11824
rect 400858 11812 400864 11824
rect 156104 11784 400864 11812
rect 156104 11772 156110 11784
rect 400858 11772 400864 11784
rect 400916 11772 400922 11824
rect 63218 11704 63224 11756
rect 63276 11744 63282 11756
rect 129918 11744 129924 11756
rect 63276 11716 129924 11744
rect 63276 11704 63282 11716
rect 129918 11704 129924 11716
rect 129976 11704 129982 11756
rect 138198 11704 138204 11756
rect 138256 11744 138262 11756
rect 167178 11744 167184 11756
rect 138256 11716 167184 11744
rect 138256 11704 138262 11716
rect 167178 11704 167184 11716
rect 167236 11704 167242 11756
rect 169846 11704 169852 11756
rect 169904 11744 169910 11756
rect 574646 11744 574652 11756
rect 169904 11716 574652 11744
rect 169904 11704 169910 11716
rect 574646 11704 574652 11716
rect 574704 11704 574710 11756
rect 234614 11636 234620 11688
rect 234672 11676 234678 11688
rect 235810 11676 235816 11688
rect 234672 11648 235816 11676
rect 234672 11636 234678 11648
rect 235810 11636 235816 11648
rect 235868 11636 235874 11688
rect 259454 11636 259460 11688
rect 259512 11676 259518 11688
rect 260650 11676 260656 11688
rect 259512 11648 260656 11676
rect 259512 11636 259518 11648
rect 260650 11636 260656 11648
rect 260708 11636 260714 11688
rect 150526 10412 150532 10464
rect 150584 10452 150590 10464
rect 322106 10452 322112 10464
rect 150584 10424 322112 10452
rect 150584 10412 150590 10424
rect 322106 10412 322112 10424
rect 322164 10412 322170 10464
rect 117314 10344 117320 10396
rect 117372 10384 117378 10396
rect 134058 10384 134064 10396
rect 117372 10356 134064 10384
rect 117372 10344 117378 10356
rect 134058 10344 134064 10356
rect 134116 10344 134122 10396
rect 154666 10344 154672 10396
rect 154724 10384 154730 10396
rect 379514 10384 379520 10396
rect 154724 10356 379520 10384
rect 154724 10344 154730 10356
rect 379514 10344 379520 10356
rect 379572 10344 379578 10396
rect 25314 10276 25320 10328
rect 25372 10316 25378 10328
rect 93118 10316 93124 10328
rect 25372 10288 93124 10316
rect 25372 10276 25378 10288
rect 93118 10276 93124 10288
rect 93176 10276 93182 10328
rect 99834 10276 99840 10328
rect 99892 10316 99898 10328
rect 132678 10316 132684 10328
rect 99892 10288 132684 10316
rect 99892 10276 99898 10288
rect 132678 10276 132684 10288
rect 132736 10276 132742 10328
rect 168190 10276 168196 10328
rect 168248 10316 168254 10328
rect 539686 10316 539692 10328
rect 168248 10288 539692 10316
rect 168248 10276 168254 10288
rect 539686 10276 539692 10288
rect 539744 10276 539750 10328
rect 147030 9392 147036 9444
rect 147088 9432 147094 9444
rect 270034 9432 270040 9444
rect 147088 9404 270040 9432
rect 147088 9392 147094 9404
rect 270034 9392 270040 9404
rect 270092 9392 270098 9444
rect 146846 9324 146852 9376
rect 146904 9364 146910 9376
rect 277118 9364 277124 9376
rect 146904 9336 277124 9364
rect 146904 9324 146910 9336
rect 277118 9324 277124 9336
rect 277176 9324 277182 9376
rect 146938 9256 146944 9308
rect 146996 9296 147002 9308
rect 276014 9296 276020 9308
rect 146996 9268 276020 9296
rect 146996 9256 147002 9268
rect 276014 9256 276020 9268
rect 276072 9256 276078 9308
rect 149146 9188 149152 9240
rect 149204 9228 149210 9240
rect 315022 9228 315028 9240
rect 149204 9200 315028 9228
rect 149204 9188 149210 9200
rect 315022 9188 315028 9200
rect 315080 9188 315086 9240
rect 315298 9188 315304 9240
rect 315356 9228 315362 9240
rect 465166 9228 465172 9240
rect 315356 9200 465172 9228
rect 315356 9188 315362 9200
rect 465166 9188 465172 9200
rect 465224 9188 465230 9240
rect 153286 9120 153292 9172
rect 153344 9160 153350 9172
rect 358722 9160 358728 9172
rect 153344 9132 358728 9160
rect 153344 9120 153350 9132
rect 358722 9120 358728 9132
rect 358780 9120 358786 9172
rect 85666 9052 85672 9104
rect 85724 9092 85730 9104
rect 131482 9092 131488 9104
rect 85724 9064 131488 9092
rect 85724 9052 85730 9064
rect 131482 9052 131488 9064
rect 131540 9052 131546 9104
rect 161934 9052 161940 9104
rect 161992 9092 161998 9104
rect 463970 9092 463976 9104
rect 161992 9064 463976 9092
rect 161992 9052 161998 9064
rect 463970 9052 463976 9064
rect 464028 9052 464034 9104
rect 78582 8984 78588 9036
rect 78640 9024 78646 9036
rect 128354 9024 128360 9036
rect 78640 8996 128360 9024
rect 78640 8984 78646 8996
rect 128354 8984 128360 8996
rect 128412 8984 128418 9036
rect 162026 8984 162032 9036
rect 162084 9024 162090 9036
rect 467466 9024 467472 9036
rect 162084 8996 467472 9024
rect 162084 8984 162090 8996
rect 467466 8984 467472 8996
rect 467524 8984 467530 9036
rect 64322 8916 64328 8968
rect 64380 8956 64386 8968
rect 126238 8956 126244 8968
rect 64380 8928 126244 8956
rect 64380 8916 64386 8928
rect 126238 8916 126244 8928
rect 126296 8916 126302 8968
rect 165614 8916 165620 8968
rect 165672 8956 165678 8968
rect 521838 8956 521844 8968
rect 165672 8928 521844 8956
rect 165672 8916 165678 8928
rect 521838 8916 521844 8928
rect 521896 8916 521902 8968
rect 142154 7896 142160 7948
rect 142212 7936 142218 7948
rect 222746 7936 222752 7948
rect 142212 7908 222752 7936
rect 142212 7896 142218 7908
rect 222746 7896 222752 7908
rect 222804 7896 222810 7948
rect 53742 7828 53748 7880
rect 53800 7868 53806 7880
rect 129182 7868 129188 7880
rect 53800 7840 129188 7868
rect 53800 7828 53806 7840
rect 129182 7828 129188 7840
rect 129240 7828 129246 7880
rect 149054 7828 149060 7880
rect 149112 7868 149118 7880
rect 307938 7868 307944 7880
rect 149112 7840 307944 7868
rect 149112 7828 149118 7840
rect 307938 7828 307944 7840
rect 307996 7828 308002 7880
rect 45462 7760 45468 7812
rect 45520 7800 45526 7812
rect 128814 7800 128820 7812
rect 45520 7772 128820 7800
rect 45520 7760 45526 7772
rect 128814 7760 128820 7772
rect 128872 7760 128878 7812
rect 150434 7760 150440 7812
rect 150492 7800 150498 7812
rect 323302 7800 323308 7812
rect 150492 7772 323308 7800
rect 150492 7760 150498 7772
rect 323302 7760 323308 7772
rect 323360 7760 323366 7812
rect 35986 7692 35992 7744
rect 36044 7732 36050 7744
rect 127250 7732 127256 7744
rect 36044 7704 127256 7732
rect 36044 7692 36050 7704
rect 127250 7692 127256 7704
rect 127308 7692 127314 7744
rect 154574 7692 154580 7744
rect 154632 7732 154638 7744
rect 385954 7732 385960 7744
rect 154632 7704 385960 7732
rect 154632 7692 154638 7704
rect 385954 7692 385960 7704
rect 386012 7692 386018 7744
rect 34790 7624 34796 7676
rect 34848 7664 34854 7676
rect 127802 7664 127808 7676
rect 34848 7636 127808 7664
rect 34848 7624 34854 7636
rect 127802 7624 127808 7636
rect 127860 7624 127866 7676
rect 172238 7624 172244 7676
rect 172296 7664 172302 7676
rect 440326 7664 440332 7676
rect 172296 7636 440332 7664
rect 172296 7624 172302 7636
rect 440326 7624 440332 7636
rect 440384 7624 440390 7676
rect 24210 7556 24216 7608
rect 24268 7596 24274 7608
rect 122190 7596 122196 7608
rect 24268 7568 122196 7596
rect 24268 7556 24274 7568
rect 122190 7556 122196 7568
rect 122248 7556 122254 7608
rect 164234 7556 164240 7608
rect 164292 7596 164298 7608
rect 504174 7596 504180 7608
rect 164292 7568 504180 7596
rect 164292 7556 164298 7568
rect 504174 7556 504180 7568
rect 504232 7556 504238 7608
rect 102134 7488 102140 7540
rect 102192 7528 102198 7540
rect 103330 7528 103336 7540
rect 102192 7500 103336 7528
rect 102192 7488 102198 7500
rect 103330 7488 103336 7500
rect 103388 7488 103394 7540
rect 146662 6808 146668 6860
rect 146720 6848 146726 6860
rect 268838 6848 268844 6860
rect 146720 6820 268844 6848
rect 146720 6808 146726 6820
rect 268838 6808 268844 6820
rect 268896 6808 268902 6860
rect 146570 6740 146576 6792
rect 146628 6780 146634 6792
rect 272426 6780 272432 6792
rect 146628 6752 272432 6780
rect 146628 6740 146634 6752
rect 272426 6740 272432 6752
rect 272484 6740 272490 6792
rect 146754 6672 146760 6724
rect 146812 6712 146818 6724
rect 273622 6712 273628 6724
rect 146812 6684 273628 6712
rect 146812 6672 146818 6684
rect 273622 6672 273628 6684
rect 273680 6672 273686 6724
rect 147858 6604 147864 6656
rect 147916 6644 147922 6656
rect 296070 6644 296076 6656
rect 147916 6616 296076 6644
rect 147916 6604 147922 6616
rect 296070 6604 296076 6616
rect 296128 6604 296134 6656
rect 105722 6536 105728 6588
rect 105780 6576 105786 6588
rect 133046 6576 133052 6588
rect 105780 6548 133052 6576
rect 105780 6536 105786 6548
rect 133046 6536 133052 6548
rect 133104 6536 133110 6588
rect 155954 6536 155960 6588
rect 156012 6576 156018 6588
rect 394234 6576 394240 6588
rect 156012 6548 394240 6576
rect 156012 6536 156018 6548
rect 394234 6536 394240 6548
rect 394292 6536 394298 6588
rect 84470 6468 84476 6520
rect 84528 6508 84534 6520
rect 131758 6508 131764 6520
rect 84528 6480 131764 6508
rect 84528 6468 84534 6480
rect 131758 6468 131764 6480
rect 131816 6468 131822 6520
rect 161750 6468 161756 6520
rect 161808 6508 161814 6520
rect 462774 6508 462780 6520
rect 161808 6480 462780 6508
rect 161808 6468 161814 6480
rect 462774 6468 462780 6480
rect 462832 6468 462838 6520
rect 80882 6400 80888 6452
rect 80940 6440 80946 6452
rect 131666 6440 131672 6452
rect 80940 6412 131672 6440
rect 80940 6400 80946 6412
rect 131666 6400 131672 6412
rect 131724 6400 131730 6452
rect 161842 6400 161848 6452
rect 161900 6440 161906 6452
rect 466270 6440 466276 6452
rect 161900 6412 466276 6440
rect 161900 6400 161906 6412
rect 466270 6400 466276 6412
rect 466328 6400 466334 6452
rect 77386 6332 77392 6384
rect 77444 6372 77450 6384
rect 131390 6372 131396 6384
rect 77444 6344 131396 6372
rect 77444 6332 77450 6344
rect 131390 6332 131396 6344
rect 131448 6332 131454 6384
rect 161566 6332 161572 6384
rect 161624 6372 161630 6384
rect 469858 6372 469864 6384
rect 161624 6344 469864 6372
rect 161624 6332 161630 6344
rect 469858 6332 469864 6344
rect 469916 6332 469922 6384
rect 52546 6264 52552 6316
rect 52604 6304 52610 6316
rect 128722 6304 128728 6316
rect 52604 6276 128728 6304
rect 52604 6264 52610 6276
rect 128722 6264 128728 6276
rect 128780 6264 128786 6316
rect 161474 6264 161480 6316
rect 161532 6304 161538 6316
rect 471054 6304 471060 6316
rect 161532 6276 471060 6304
rect 161532 6264 161538 6276
rect 471054 6264 471060 6276
rect 471112 6264 471118 6316
rect 19426 6196 19432 6248
rect 19484 6236 19490 6248
rect 125042 6236 125048 6248
rect 19484 6208 125048 6236
rect 19484 6196 19490 6208
rect 125042 6196 125048 6208
rect 125100 6196 125106 6248
rect 161658 6196 161664 6248
rect 161716 6236 161722 6248
rect 473446 6236 473452 6248
rect 161716 6208 473452 6236
rect 161716 6196 161722 6208
rect 473446 6196 473452 6208
rect 473504 6196 473510 6248
rect 18230 6128 18236 6180
rect 18288 6168 18294 6180
rect 125870 6168 125876 6180
rect 18288 6140 125876 6168
rect 18288 6128 18294 6140
rect 125870 6128 125876 6140
rect 125928 6128 125934 6180
rect 169754 6128 169760 6180
rect 169812 6168 169818 6180
rect 572714 6168 572720 6180
rect 169812 6140 572720 6168
rect 169812 6128 169818 6140
rect 572714 6128 572720 6140
rect 572772 6128 572778 6180
rect 132402 6060 132408 6112
rect 132460 6100 132466 6112
rect 190822 6100 190828 6112
rect 132460 6072 190828 6100
rect 132460 6060 132466 6072
rect 190822 6060 190828 6072
rect 190880 6060 190886 6112
rect 136726 5176 136732 5228
rect 136784 5216 136790 5228
rect 154206 5216 154212 5228
rect 136784 5188 154212 5216
rect 136784 5176 136790 5188
rect 154206 5176 154212 5188
rect 154264 5176 154270 5228
rect 101398 5108 101404 5160
rect 101456 5148 101462 5160
rect 113818 5148 113824 5160
rect 101456 5120 113824 5148
rect 101456 5108 101462 5120
rect 113818 5108 113824 5120
rect 113876 5108 113882 5160
rect 114002 5108 114008 5160
rect 114060 5148 114066 5160
rect 134426 5148 134432 5160
rect 114060 5120 134432 5148
rect 114060 5108 114066 5120
rect 134426 5108 134432 5120
rect 134484 5108 134490 5160
rect 138014 5108 138020 5160
rect 138072 5148 138078 5160
rect 169570 5148 169576 5160
rect 138072 5120 169576 5148
rect 138072 5108 138078 5120
rect 169570 5108 169576 5120
rect 169628 5108 169634 5160
rect 66714 5040 66720 5092
rect 66772 5080 66778 5092
rect 103514 5080 103520 5092
rect 66772 5052 103520 5080
rect 66772 5040 66778 5052
rect 103514 5040 103520 5052
rect 103572 5040 103578 5092
rect 103698 5040 103704 5092
rect 103756 5080 103762 5092
rect 130286 5080 130292 5092
rect 103756 5052 130292 5080
rect 103756 5040 103762 5052
rect 130286 5040 130292 5052
rect 130344 5040 130350 5092
rect 140774 5040 140780 5092
rect 140832 5080 140838 5092
rect 206186 5080 206192 5092
rect 140832 5052 206192 5080
rect 140832 5040 140838 5052
rect 206186 5040 206192 5052
rect 206244 5040 206250 5092
rect 15930 4972 15936 5024
rect 15988 5012 15994 5024
rect 101398 5012 101404 5024
rect 15988 4984 101404 5012
rect 15988 4972 15994 4984
rect 101398 4972 101404 4984
rect 101456 4972 101462 5024
rect 147766 4972 147772 5024
rect 147824 5012 147830 5024
rect 294874 5012 294880 5024
rect 147824 4984 294880 5012
rect 147824 4972 147830 4984
rect 294874 4972 294880 4984
rect 294932 4972 294938 5024
rect 436738 4972 436744 5024
rect 436796 5012 436802 5024
rect 436796 4984 451274 5012
rect 436796 4972 436802 4984
rect 28902 4904 28908 4956
rect 28960 4944 28966 4956
rect 127710 4944 127716 4956
rect 28960 4916 127716 4944
rect 28960 4904 28966 4916
rect 127710 4904 127716 4916
rect 127768 4904 127774 4956
rect 154390 4904 154396 4956
rect 154448 4944 154454 4956
rect 364610 4944 364616 4956
rect 154448 4916 364616 4944
rect 154448 4904 154454 4916
rect 364610 4904 364616 4916
rect 364668 4904 364674 4956
rect 6454 4836 6460 4888
rect 6512 4876 6518 4888
rect 10318 4876 10324 4888
rect 6512 4848 10324 4876
rect 6512 4836 6518 4848
rect 10318 4836 10324 4848
rect 10376 4836 10382 4888
rect 13538 4836 13544 4888
rect 13596 4876 13602 4888
rect 125778 4876 125784 4888
rect 13596 4848 125784 4876
rect 13596 4836 13602 4848
rect 125778 4836 125784 4848
rect 125836 4836 125842 4888
rect 136634 4836 136640 4888
rect 136692 4876 136698 4888
rect 157794 4876 157800 4888
rect 136692 4848 157800 4876
rect 136692 4836 136698 4848
rect 157794 4836 157800 4848
rect 157852 4836 157858 4888
rect 159818 4836 159824 4888
rect 159876 4876 159882 4888
rect 436738 4876 436744 4888
rect 159876 4848 436744 4876
rect 159876 4836 159882 4848
rect 436738 4836 436744 4848
rect 436796 4836 436802 4888
rect 451246 4876 451274 4984
rect 479334 4876 479340 4888
rect 451246 4848 479340 4876
rect 479334 4836 479340 4848
rect 479392 4836 479398 4888
rect 8754 4768 8760 4820
rect 8812 4808 8818 4820
rect 126422 4808 126428 4820
rect 8812 4780 126428 4808
rect 8812 4768 8818 4780
rect 126422 4768 126428 4780
rect 126480 4768 126486 4820
rect 138106 4768 138112 4820
rect 138164 4808 138170 4820
rect 162486 4808 162492 4820
rect 138164 4780 162492 4808
rect 138164 4768 138170 4780
rect 162486 4768 162492 4780
rect 162544 4768 162550 4820
rect 162854 4768 162860 4820
rect 162912 4808 162918 4820
rect 493502 4808 493508 4820
rect 162912 4780 493508 4808
rect 162912 4768 162918 4780
rect 493502 4768 493508 4780
rect 493560 4768 493566 4820
rect 566 4088 572 4140
rect 624 4128 630 4140
rect 7558 4128 7564 4140
rect 624 4100 7564 4128
rect 624 4088 630 4100
rect 7558 4088 7564 4100
rect 7616 4088 7622 4140
rect 135622 4088 135628 4140
rect 135680 4128 135686 4140
rect 136542 4128 136548 4140
rect 135680 4100 136548 4128
rect 135680 4088 135686 4100
rect 136542 4088 136548 4100
rect 136600 4088 136606 4140
rect 140314 4088 140320 4140
rect 140372 4128 140378 4140
rect 186130 4128 186136 4140
rect 140372 4100 186136 4128
rect 140372 4088 140378 4100
rect 186130 4088 186136 4100
rect 186188 4088 186194 4140
rect 139486 4020 139492 4072
rect 139544 4060 139550 4072
rect 189718 4060 189724 4072
rect 139544 4032 189724 4060
rect 139544 4020 139550 4032
rect 189718 4020 189724 4032
rect 189776 4020 189782 4072
rect 251174 4020 251180 4072
rect 251232 4060 251238 4072
rect 252370 4060 252376 4072
rect 251232 4032 252376 4060
rect 251232 4020 251238 4032
rect 252370 4020 252376 4032
rect 252428 4020 252434 4072
rect 146386 3952 146392 4004
rect 146444 3992 146450 4004
rect 271230 3992 271236 4004
rect 146444 3964 271236 3992
rect 146444 3952 146450 3964
rect 271230 3952 271236 3964
rect 271288 3952 271294 4004
rect 146478 3884 146484 3936
rect 146536 3924 146542 3936
rect 274818 3924 274824 3936
rect 146536 3896 274824 3924
rect 146536 3884 146542 3896
rect 274818 3884 274824 3896
rect 274876 3884 274882 3936
rect 102226 3816 102232 3868
rect 102284 3856 102290 3868
rect 124858 3856 124864 3868
rect 102284 3828 124864 3856
rect 102284 3816 102290 3828
rect 124858 3816 124864 3828
rect 124916 3816 124922 3868
rect 146294 3816 146300 3868
rect 146352 3856 146358 3868
rect 278314 3856 278320 3868
rect 146352 3828 278320 3856
rect 146352 3816 146358 3828
rect 278314 3816 278320 3828
rect 278372 3816 278378 3868
rect 284294 3816 284300 3868
rect 284352 3856 284358 3868
rect 285030 3856 285036 3868
rect 284352 3828 285036 3856
rect 284352 3816 284358 3828
rect 285030 3816 285036 3828
rect 285088 3816 285094 3868
rect 87966 3748 87972 3800
rect 88024 3788 88030 3800
rect 123478 3788 123484 3800
rect 88024 3760 123484 3788
rect 88024 3748 88030 3760
rect 123478 3748 123484 3760
rect 123536 3748 123542 3800
rect 147674 3748 147680 3800
rect 147732 3788 147738 3800
rect 292574 3788 292580 3800
rect 147732 3760 292580 3788
rect 147732 3748 147738 3760
rect 292574 3748 292580 3760
rect 292632 3748 292638 3800
rect 461578 3788 461584 3800
rect 451246 3760 461584 3788
rect 65518 3680 65524 3732
rect 65576 3720 65582 3732
rect 122374 3720 122380 3732
rect 65576 3692 122380 3720
rect 65576 3680 65582 3692
rect 122374 3680 122380 3692
rect 122432 3680 122438 3732
rect 173158 3680 173164 3732
rect 173216 3720 173222 3732
rect 451246 3720 451274 3760
rect 461578 3748 461584 3760
rect 461636 3748 461642 3800
rect 173216 3692 451274 3720
rect 173216 3680 173222 3692
rect 462222 3680 462228 3732
rect 462280 3720 462286 3732
rect 577406 3720 577412 3732
rect 462280 3692 577412 3720
rect 462280 3680 462286 3692
rect 577406 3680 577412 3692
rect 577464 3680 577470 3732
rect 2866 3612 2872 3664
rect 2924 3652 2930 3664
rect 120718 3652 120724 3664
rect 2924 3624 120724 3652
rect 2924 3612 2930 3624
rect 120718 3612 120724 3624
rect 120776 3612 120782 3664
rect 135530 3612 135536 3664
rect 135588 3652 135594 3664
rect 138842 3652 138848 3664
rect 135588 3624 138848 3652
rect 135588 3612 135594 3624
rect 138842 3612 138848 3624
rect 138900 3612 138906 3664
rect 142982 3612 142988 3664
rect 143040 3652 143046 3664
rect 155402 3652 155408 3664
rect 143040 3624 155408 3652
rect 143040 3612 143046 3624
rect 155402 3612 155408 3624
rect 155460 3612 155466 3664
rect 171778 3612 171784 3664
rect 171836 3652 171842 3664
rect 472250 3652 472256 3664
rect 171836 3624 472256 3652
rect 171836 3612 171842 3624
rect 472250 3612 472256 3624
rect 472308 3612 472314 3664
rect 5258 3544 5264 3596
rect 5316 3584 5322 3596
rect 122098 3584 122104 3596
rect 5316 3556 122104 3584
rect 5316 3544 5322 3556
rect 122098 3544 122104 3556
rect 122156 3544 122162 3596
rect 129366 3544 129372 3596
rect 129424 3584 129430 3596
rect 130378 3584 130384 3596
rect 129424 3556 130384 3584
rect 129424 3544 129430 3556
rect 130378 3544 130384 3556
rect 130436 3544 130442 3596
rect 135438 3544 135444 3596
rect 135496 3584 135502 3596
rect 137646 3584 137652 3596
rect 135496 3556 137652 3584
rect 135496 3544 135502 3556
rect 137646 3544 137652 3556
rect 137704 3544 137710 3596
rect 138750 3544 138756 3596
rect 138808 3584 138814 3596
rect 151814 3584 151820 3596
rect 138808 3556 151820 3584
rect 138808 3544 138814 3556
rect 151814 3544 151820 3556
rect 151872 3544 151878 3596
rect 152458 3544 152464 3596
rect 152516 3584 152522 3596
rect 160094 3584 160100 3596
rect 152516 3556 160100 3584
rect 152516 3544 152522 3556
rect 160094 3544 160100 3556
rect 160152 3544 160158 3596
rect 172146 3544 172152 3596
rect 172204 3584 172210 3596
rect 475746 3584 475752 3596
rect 172204 3556 475752 3584
rect 172204 3544 172210 3556
rect 475746 3544 475752 3556
rect 475804 3544 475810 3596
rect 481634 3544 481640 3596
rect 481692 3584 481698 3596
rect 482462 3584 482468 3596
rect 481692 3556 482468 3584
rect 481692 3544 481698 3556
rect 482462 3544 482468 3556
rect 482520 3544 482526 3596
rect 506474 3544 506480 3596
rect 506532 3584 506538 3596
rect 507302 3584 507308 3596
rect 506532 3556 507308 3584
rect 506532 3544 506538 3556
rect 507302 3544 507308 3556
rect 507360 3544 507366 3596
rect 574738 3544 574744 3596
rect 574796 3584 574802 3596
rect 574796 3556 576854 3584
rect 574796 3544 574802 3556
rect 11054 3476 11060 3528
rect 11112 3516 11118 3528
rect 11974 3516 11980 3528
rect 11112 3488 11980 3516
rect 11112 3476 11118 3488
rect 11974 3476 11980 3488
rect 12032 3476 12038 3528
rect 124950 3516 124956 3528
rect 16546 3488 124956 3516
rect 7650 3408 7656 3460
rect 7708 3448 7714 3460
rect 16546 3448 16574 3488
rect 124950 3476 124956 3488
rect 125008 3476 125014 3528
rect 140130 3476 140136 3528
rect 140188 3516 140194 3528
rect 163682 3516 163688 3528
rect 140188 3488 163688 3516
rect 140188 3476 140194 3488
rect 163682 3476 163688 3488
rect 163740 3476 163746 3528
rect 171962 3476 171968 3528
rect 172020 3516 172026 3528
rect 174262 3516 174268 3528
rect 172020 3488 174268 3516
rect 172020 3476 172026 3488
rect 174262 3476 174268 3488
rect 174320 3476 174326 3528
rect 176654 3476 176660 3528
rect 176712 3516 176718 3528
rect 177850 3516 177856 3528
rect 176712 3488 177856 3516
rect 176712 3476 176718 3488
rect 177850 3476 177856 3488
rect 177908 3476 177914 3528
rect 177942 3476 177948 3528
rect 178000 3516 178006 3528
rect 519538 3516 519544 3528
rect 178000 3488 519544 3516
rect 178000 3476 178006 3488
rect 519538 3476 519544 3488
rect 519596 3476 519602 3528
rect 531314 3476 531320 3528
rect 531372 3516 531378 3528
rect 532142 3516 532148 3528
rect 531372 3488 532148 3516
rect 531372 3476 531378 3488
rect 532142 3476 532148 3488
rect 532200 3476 532206 3528
rect 539594 3476 539600 3528
rect 539652 3516 539658 3528
rect 540422 3516 540428 3528
rect 539652 3488 540428 3516
rect 539652 3476 539658 3488
rect 540422 3476 540428 3488
rect 540480 3476 540486 3528
rect 564434 3476 564440 3528
rect 564492 3516 564498 3528
rect 565262 3516 565268 3528
rect 564492 3488 565268 3516
rect 564492 3476 564498 3488
rect 565262 3476 565268 3488
rect 565320 3476 565326 3528
rect 7708 3420 16574 3448
rect 7708 3408 7714 3420
rect 62022 3408 62028 3460
rect 62080 3448 62086 3460
rect 62080 3420 99374 3448
rect 62080 3408 62086 3420
rect 69014 3340 69020 3392
rect 69072 3380 69078 3392
rect 69934 3380 69940 3392
rect 69072 3352 69940 3380
rect 69072 3340 69078 3352
rect 69934 3340 69940 3352
rect 69992 3340 69998 3392
rect 93854 3340 93860 3392
rect 93912 3380 93918 3392
rect 94774 3380 94780 3392
rect 93912 3352 94780 3380
rect 93912 3340 93918 3352
rect 94774 3340 94780 3352
rect 94832 3340 94838 3392
rect 99346 3380 99374 3420
rect 110414 3408 110420 3460
rect 110472 3448 110478 3460
rect 111610 3448 111616 3460
rect 110472 3420 111616 3448
rect 110472 3408 110478 3420
rect 111610 3408 111616 3420
rect 111668 3408 111674 3460
rect 118694 3408 118700 3460
rect 118752 3448 118758 3460
rect 119890 3448 119896 3460
rect 118752 3420 119896 3448
rect 118752 3408 118758 3420
rect 119890 3408 119896 3420
rect 119948 3408 119954 3460
rect 140222 3408 140228 3460
rect 140280 3448 140286 3460
rect 164878 3448 164884 3460
rect 140280 3420 164884 3448
rect 140280 3408 140286 3420
rect 164878 3408 164884 3420
rect 164936 3408 164942 3460
rect 173250 3408 173256 3460
rect 173308 3448 173314 3460
rect 526622 3448 526628 3460
rect 173308 3420 526628 3448
rect 173308 3408 173314 3420
rect 526622 3408 526628 3420
rect 526680 3408 526686 3460
rect 576826 3448 576854 3556
rect 580994 3448 581000 3460
rect 576826 3420 581000 3448
rect 580994 3408 581000 3420
rect 581052 3408 581058 3460
rect 119338 3380 119344 3392
rect 99346 3352 119344 3380
rect 119338 3340 119344 3352
rect 119396 3340 119402 3392
rect 144178 3340 144184 3392
rect 144236 3380 144242 3392
rect 149514 3380 149520 3392
rect 144236 3352 149520 3380
rect 144236 3340 144242 3352
rect 149514 3340 149520 3352
rect 149572 3340 149578 3392
rect 153010 3380 153016 3392
rect 151786 3352 153016 3380
rect 136542 3272 136548 3324
rect 136600 3312 136606 3324
rect 142430 3312 142436 3324
rect 136600 3284 142436 3312
rect 136600 3272 136606 3284
rect 142430 3272 142436 3284
rect 142488 3272 142494 3324
rect 142798 3272 142804 3324
rect 142856 3312 142862 3324
rect 150618 3312 150624 3324
rect 142856 3284 150624 3312
rect 142856 3272 142862 3284
rect 150618 3272 150624 3284
rect 150676 3272 150682 3324
rect 118786 3204 118792 3256
rect 118844 3244 118850 3256
rect 123570 3244 123576 3256
rect 118844 3216 123576 3244
rect 118844 3204 118850 3216
rect 123570 3204 123576 3216
rect 123628 3204 123634 3256
rect 140038 3204 140044 3256
rect 140096 3244 140102 3256
rect 144730 3244 144736 3256
rect 140096 3216 144736 3244
rect 140096 3204 140102 3216
rect 144730 3204 144736 3216
rect 144788 3204 144794 3256
rect 144454 3136 144460 3188
rect 144512 3176 144518 3188
rect 151786 3176 151814 3352
rect 153010 3340 153016 3352
rect 153068 3340 153074 3392
rect 166258 3340 166264 3392
rect 166316 3380 166322 3392
rect 170766 3380 170772 3392
rect 166316 3352 170772 3380
rect 166316 3340 166322 3352
rect 170766 3340 170772 3352
rect 170824 3340 170830 3392
rect 175918 3340 175924 3392
rect 175976 3380 175982 3392
rect 212166 3380 212172 3392
rect 175976 3352 212172 3380
rect 175976 3340 175982 3352
rect 212166 3340 212172 3352
rect 212224 3340 212230 3392
rect 307754 3340 307760 3392
rect 307812 3380 307818 3392
rect 309042 3380 309048 3392
rect 307812 3352 309048 3380
rect 307812 3340 307818 3352
rect 309042 3340 309048 3352
rect 309100 3340 309106 3392
rect 316034 3340 316040 3392
rect 316092 3380 316098 3392
rect 317322 3380 317328 3392
rect 316092 3352 317328 3380
rect 316092 3340 316098 3352
rect 317322 3340 317328 3352
rect 317380 3340 317386 3392
rect 324406 3340 324412 3392
rect 324464 3380 324470 3392
rect 325602 3380 325608 3392
rect 324464 3352 325608 3380
rect 324464 3340 324470 3352
rect 325602 3340 325608 3352
rect 325660 3340 325666 3392
rect 332594 3340 332600 3392
rect 332652 3380 332658 3392
rect 333882 3380 333888 3392
rect 332652 3352 333888 3380
rect 332652 3340 332658 3352
rect 333882 3340 333888 3352
rect 333940 3340 333946 3392
rect 340966 3340 340972 3392
rect 341024 3380 341030 3392
rect 342162 3380 342168 3392
rect 341024 3352 342168 3380
rect 341024 3340 341030 3352
rect 342162 3340 342168 3352
rect 342220 3340 342226 3392
rect 349246 3340 349252 3392
rect 349304 3380 349310 3392
rect 350442 3380 350448 3392
rect 349304 3352 350448 3380
rect 349304 3340 349310 3352
rect 350442 3340 350448 3352
rect 350500 3340 350506 3392
rect 365714 3340 365720 3392
rect 365772 3380 365778 3392
rect 367002 3380 367008 3392
rect 365772 3352 367008 3380
rect 365772 3340 365778 3352
rect 367002 3340 367008 3352
rect 367060 3340 367066 3392
rect 374086 3340 374092 3392
rect 374144 3380 374150 3392
rect 375282 3380 375288 3392
rect 374144 3352 375288 3380
rect 374144 3340 374150 3352
rect 375282 3340 375288 3352
rect 375340 3340 375346 3392
rect 382366 3340 382372 3392
rect 382424 3380 382430 3392
rect 383562 3380 383568 3392
rect 382424 3352 383568 3380
rect 382424 3340 382430 3352
rect 383562 3340 383568 3352
rect 383620 3340 383626 3392
rect 390646 3340 390652 3392
rect 390704 3380 390710 3392
rect 391842 3380 391848 3392
rect 390704 3352 391848 3380
rect 390704 3340 390710 3352
rect 391842 3340 391848 3352
rect 391900 3340 391906 3392
rect 398926 3340 398932 3392
rect 398984 3380 398990 3392
rect 400122 3380 400128 3392
rect 398984 3352 400128 3380
rect 398984 3340 398990 3352
rect 400122 3340 400128 3352
rect 400180 3340 400186 3392
rect 407114 3340 407120 3392
rect 407172 3380 407178 3392
rect 408402 3380 408408 3392
rect 407172 3352 408408 3380
rect 407172 3340 407178 3352
rect 408402 3340 408408 3352
rect 408460 3340 408466 3392
rect 415394 3340 415400 3392
rect 415452 3380 415458 3392
rect 416682 3380 416688 3392
rect 415452 3352 416688 3380
rect 415452 3340 415458 3352
rect 416682 3340 416688 3352
rect 416740 3340 416746 3392
rect 423766 3340 423772 3392
rect 423824 3380 423830 3392
rect 424962 3380 424968 3392
rect 423824 3352 424968 3380
rect 423824 3340 423830 3352
rect 424962 3340 424968 3352
rect 425020 3340 425026 3392
rect 432046 3340 432052 3392
rect 432104 3380 432110 3392
rect 433242 3380 433248 3392
rect 432104 3352 433248 3380
rect 432104 3340 432110 3352
rect 433242 3340 433248 3352
rect 433300 3340 433306 3392
rect 440234 3340 440240 3392
rect 440292 3380 440298 3392
rect 441522 3380 441528 3392
rect 440292 3352 441528 3380
rect 440292 3340 440298 3352
rect 441522 3340 441528 3352
rect 441580 3340 441586 3392
rect 448606 3340 448612 3392
rect 448664 3380 448670 3392
rect 449802 3380 449808 3392
rect 448664 3352 449808 3380
rect 448664 3340 448670 3352
rect 449802 3340 449808 3352
rect 449860 3340 449866 3392
rect 456886 3340 456892 3392
rect 456944 3380 456950 3392
rect 458082 3380 458088 3392
rect 456944 3352 458088 3380
rect 456944 3340 456950 3352
rect 458082 3340 458088 3352
rect 458140 3340 458146 3392
rect 174538 3272 174544 3324
rect 174596 3312 174602 3324
rect 195606 3312 195612 3324
rect 174596 3284 195612 3312
rect 174596 3272 174602 3284
rect 195606 3272 195612 3284
rect 195664 3272 195670 3324
rect 171870 3204 171876 3256
rect 171928 3244 171934 3256
rect 177942 3244 177948 3256
rect 171928 3216 177948 3244
rect 171928 3204 171934 3216
rect 177942 3204 177948 3216
rect 178000 3204 178006 3256
rect 144512 3148 151814 3176
rect 144512 3136 144518 3148
rect 165062 3068 165068 3120
rect 165120 3108 165126 3120
rect 171962 3108 171968 3120
rect 165120 3080 171968 3108
rect 165120 3068 165126 3080
rect 171962 3068 171968 3080
rect 172020 3068 172026 3120
<< via1 >>
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 201500 702992 201552 703044
rect 202788 702992 202840 703044
rect 331220 702992 331272 703044
rect 332508 702992 332560 703044
rect 196624 700612 196676 700664
rect 218980 700612 219032 700664
rect 193864 700544 193916 700596
rect 283840 700544 283892 700596
rect 192484 700476 192536 700528
rect 348792 700476 348844 700528
rect 189724 700408 189776 700460
rect 413652 700408 413704 700460
rect 89168 700340 89220 700392
rect 182548 700340 182600 700392
rect 188344 700340 188396 700392
rect 478512 700340 478564 700392
rect 8116 700272 8168 700324
rect 119344 700272 119396 700324
rect 137836 700272 137888 700324
rect 180800 700272 180852 700324
rect 185584 700272 185636 700324
rect 543464 700272 543516 700324
rect 105452 699660 105504 699712
rect 106924 699660 106976 699712
rect 266360 697552 266412 697604
rect 267648 697552 267700 697604
rect 2780 683680 2832 683732
rect 4804 683680 4856 683732
rect 184204 683136 184256 683188
rect 579620 683136 579672 683188
rect 3332 632068 3384 632120
rect 7564 632068 7616 632120
rect 184296 630640 184348 630692
rect 580172 630640 580224 630692
rect 120724 616836 120776 616888
rect 579988 616836 580040 616888
rect 3148 579640 3200 579692
rect 17224 579640 17276 579692
rect 184388 576852 184440 576904
rect 579988 576852 580040 576904
rect 120816 563048 120868 563100
rect 580172 563048 580224 563100
rect 3148 553392 3200 553444
rect 115204 553392 115256 553444
rect 182364 536800 182416 536852
rect 579620 536800 579672 536852
rect 3332 527824 3384 527876
rect 8944 527824 8996 527876
rect 214564 524424 214616 524476
rect 580172 524424 580224 524476
rect 3332 514768 3384 514820
rect 180892 514768 180944 514820
rect 120908 510620 120960 510672
rect 579620 510620 579672 510672
rect 2780 501032 2832 501084
rect 4896 501032 4948 501084
rect 182272 484372 182324 484424
rect 580172 484372 580224 484424
rect 211804 470568 211856 470620
rect 579988 470568 580040 470620
rect 3056 462340 3108 462392
rect 179420 462340 179472 462392
rect 3884 461592 3936 461644
rect 53104 461592 53156 461644
rect 121000 456764 121052 456816
rect 580172 456764 580224 456816
rect 2964 448536 3016 448588
rect 44824 448536 44876 448588
rect 118700 429836 118752 429888
rect 580632 429836 580684 429888
rect 3332 422288 3384 422340
rect 10324 422288 10376 422340
rect 182824 418140 182876 418192
rect 579712 418140 579764 418192
rect 118608 404336 118660 404388
rect 580172 404336 580224 404388
rect 3332 397468 3384 397520
rect 86224 397468 86276 397520
rect 3332 371220 3384 371272
rect 84844 371220 84896 371272
rect 224224 364352 224276 364404
rect 580172 364352 580224 364404
rect 3332 357416 3384 357468
rect 180984 357416 181036 357468
rect 118516 351908 118568 351960
rect 580172 351908 580224 351960
rect 3332 345040 3384 345092
rect 116584 345040 116636 345092
rect 3148 318792 3200 318844
rect 13084 318792 13136 318844
rect 221464 311856 221516 311908
rect 580172 311856 580224 311908
rect 3332 304988 3384 305040
rect 178684 304988 178736 305040
rect 124864 298120 124916 298172
rect 580172 298120 580224 298172
rect 3332 292544 3384 292596
rect 121092 292544 121144 292596
rect 180064 271872 180116 271924
rect 579620 271872 579672 271924
rect 3240 266364 3292 266416
rect 18604 266364 18656 266416
rect 220084 258068 220136 258120
rect 580172 258068 580224 258120
rect 2964 253920 3016 253972
rect 178776 253920 178828 253972
rect 129004 244264 129056 244316
rect 579620 244264 579672 244316
rect 182180 233792 182232 233844
rect 182548 233792 182600 233844
rect 182824 231548 182876 231600
rect 182824 230324 182876 230376
rect 207664 229780 207716 229832
rect 212540 229780 212592 229832
rect 161388 229712 161440 229764
rect 392492 229712 392544 229764
rect 180156 229100 180208 229152
rect 182548 229100 182600 229152
rect 123668 228352 123720 228404
rect 143540 228352 143592 228404
rect 166264 228352 166316 228404
rect 272524 228352 272576 228404
rect 2872 227740 2924 227792
rect 138664 227740 138716 227792
rect 182180 224204 182232 224256
rect 182548 224204 182600 224256
rect 217324 218016 217376 218068
rect 579988 218016 580040 218068
rect 3332 213936 3384 213988
rect 31024 213936 31076 213988
rect 144920 208360 144972 208412
rect 151820 208360 151872 208412
rect 126244 205640 126296 205692
rect 580172 205640 580224 205692
rect 154120 204892 154172 204944
rect 242900 204892 242952 204944
rect 146208 203532 146260 203584
rect 207664 203532 207716 203584
rect 147404 202104 147456 202156
rect 180156 202104 180208 202156
rect 3332 201492 3384 201544
rect 179604 201492 179656 201544
rect 159180 199384 159232 199436
rect 362960 199384 363012 199436
rect 154580 198024 154632 198076
rect 166264 198024 166316 198076
rect 157340 197956 157392 198008
rect 332600 197956 332652 198008
rect 138664 196732 138716 196784
rect 164240 196732 164292 196784
rect 153844 196664 153896 196716
rect 181076 196664 181128 196716
rect 157248 196596 157300 196648
rect 302240 196596 302292 196648
rect 152464 196460 152516 196512
rect 154580 196460 154632 196512
rect 62120 195916 62172 195968
rect 138112 195916 138164 195968
rect 153476 195916 153528 195968
rect 154120 195916 154172 195968
rect 92480 195848 92532 195900
rect 139400 195848 139452 195900
rect 148784 195644 148836 195696
rect 165528 195644 165580 195696
rect 151452 191088 151504 191140
rect 3332 187688 3384 187740
rect 121184 187688 121236 187740
rect 144460 180684 144512 180736
rect 146116 180684 146168 180736
rect 161480 180548 161532 180600
rect 162124 180888 162176 180940
rect 17868 180072 17920 180124
rect 136824 180276 136876 180328
rect 136640 180072 136692 180124
rect 141240 180072 141292 180124
rect 143540 179596 143592 179648
rect 122840 178780 122892 178832
rect 136640 178780 136692 178832
rect 121460 178644 121512 178696
rect 137008 178644 137060 178696
rect 144184 178644 144236 178696
rect 215944 178032 215996 178084
rect 580172 178032 580224 178084
rect 140780 177828 140832 177880
rect 141608 177828 141660 177880
rect 124220 177284 124272 177336
rect 137100 177284 137152 177336
rect 3332 176604 3384 176656
rect 17868 176604 17920 176656
rect 161388 176196 161440 176248
rect 125600 175992 125652 176044
rect 137192 175992 137244 176044
rect 128360 175924 128412 175976
rect 137284 175924 137336 175976
rect 159088 175584 159140 175636
rect 165436 174972 165488 175024
rect 165528 174972 165580 175024
rect 163136 174700 163188 174752
rect 165436 174700 165488 174752
rect 165528 174700 165580 174752
rect 133880 173884 133932 173936
rect 135260 173884 135312 173936
rect 140780 173816 140832 173868
rect 141608 173816 141660 173868
rect 131120 173272 131172 173324
rect 137376 173272 137428 173324
rect 126980 173204 127032 173256
rect 140780 173204 140832 173256
rect 3792 173136 3844 173188
rect 179696 173136 179748 173188
rect 135260 172388 135312 172440
rect 138940 172388 138992 172440
rect 132500 172184 132552 172236
rect 137468 172184 137520 172236
rect 138020 171368 138072 171420
rect 140964 171368 141016 171420
rect 122104 165588 122156 165640
rect 579804 165588 579856 165640
rect 162860 164704 162912 164756
rect 163596 164704 163648 164756
rect 165528 164160 165580 164212
rect 168380 164160 168432 164212
rect 3332 162868 3384 162920
rect 14464 162868 14516 162920
rect 165436 162800 165488 162852
rect 169852 162800 169904 162852
rect 182916 151784 182968 151836
rect 579988 151784 580040 151836
rect 3700 151036 3752 151088
rect 181260 151036 181312 151088
rect 3516 150016 3568 150068
rect 3700 150016 3752 150068
rect 3516 149064 3568 149116
rect 181168 149064 181220 149116
rect 3700 148316 3752 148368
rect 181352 148316 181404 148368
rect 119068 146956 119120 147008
rect 234620 146956 234672 147008
rect 23480 146888 23532 146940
rect 179788 146888 179840 146940
rect 119160 145528 119212 145580
rect 299480 145528 299532 145580
rect 118884 144168 118936 144220
rect 429200 144168 429252 144220
rect 151820 143488 151872 143540
rect 157432 143488 157484 143540
rect 164056 143488 164108 143540
rect 166172 143488 166224 143540
rect 162768 143216 162820 143268
rect 166080 143216 166132 143268
rect 137744 143148 137796 143200
rect 139400 143148 139452 143200
rect 164240 142944 164292 142996
rect 176200 142944 176252 142996
rect 150440 142876 150492 142928
rect 154580 142876 154632 142928
rect 162860 142876 162912 142928
rect 174636 142876 174688 142928
rect 163136 142808 163188 142860
rect 178040 142808 178092 142860
rect 118240 142128 118292 142180
rect 124864 142128 124916 142180
rect 149060 142128 149112 142180
rect 152740 142128 152792 142180
rect 118148 141516 118200 141568
rect 129004 141516 129056 141568
rect 118056 141448 118108 141500
rect 169760 141448 169812 141500
rect 118976 141380 119028 141432
rect 494060 141380 494112 141432
rect 118332 140224 118384 140276
rect 126244 140224 126296 140276
rect 3884 140156 3936 140208
rect 181444 140156 181496 140208
rect 119252 140088 119304 140140
rect 364340 140088 364392 140140
rect 118792 140020 118844 140072
rect 558920 140020 558972 140072
rect 118424 139476 118476 139528
rect 122104 139476 122156 139528
rect 3516 139408 3568 139460
rect 179512 139408 179564 139460
rect 178776 139340 178828 139392
rect 182180 139340 182232 139392
rect 178684 139272 178736 139324
rect 182456 139272 182508 139324
rect 193956 137980 194008 138032
rect 580172 137980 580224 138032
rect 7656 136688 7708 136740
rect 117320 136688 117372 136740
rect 2872 136620 2924 136672
rect 115296 136620 115348 136672
rect 9036 135260 9088 135312
rect 117320 135260 117372 135312
rect 21364 133900 21416 133952
rect 117320 133900 117372 133952
rect 14464 133832 14516 133884
rect 117412 133832 117464 133884
rect 31024 132404 31076 132456
rect 117320 132404 117372 132456
rect 18604 131044 18656 131096
rect 117320 131044 117372 131096
rect 13084 129684 13136 129736
rect 117320 129684 117372 129736
rect 84844 128256 84896 128308
rect 117320 128256 117372 128308
rect 10324 126896 10376 126948
rect 117320 126896 117372 126948
rect 53104 124108 53156 124160
rect 117320 124108 117372 124160
rect 8944 122748 8996 122800
rect 117320 122748 117372 122800
rect 17224 121388 17276 121440
rect 117320 121388 117372 121440
rect 7564 120028 7616 120080
rect 117320 120028 117372 120080
rect 4804 118600 4856 118652
rect 117320 118600 117372 118652
rect 40040 117240 40092 117292
rect 117320 117240 117372 117292
rect 106924 115880 106976 115932
rect 117320 115880 117372 115932
rect 180156 111800 180208 111852
rect 580080 111800 580132 111852
rect 3332 111732 3384 111784
rect 21364 111732 21416 111784
rect 183284 108944 183336 108996
rect 196624 108944 196676 108996
rect 183284 107584 183336 107636
rect 193864 107584 193916 107636
rect 183284 106224 183336 106276
rect 192484 106224 192536 106276
rect 183284 104592 183336 104644
rect 189724 104592 189776 104644
rect 183468 102892 183520 102944
rect 188344 102892 188396 102944
rect 182640 101260 182692 101312
rect 185584 101260 185636 101312
rect 182456 100444 182508 100496
rect 184204 100444 184256 100496
rect 192484 99356 192536 99408
rect 580080 99356 580132 99408
rect 182180 99288 182232 99340
rect 184296 99288 184348 99340
rect 182180 97384 182232 97436
rect 184388 97384 184440 97436
rect 183192 96568 183244 96620
rect 214564 96568 214616 96620
rect 183468 95140 183520 95192
rect 211804 95140 211856 95192
rect 183376 93100 183428 93152
rect 224224 93100 224276 93152
rect 183468 91740 183520 91792
rect 221464 91740 221516 91792
rect 183376 90312 183428 90364
rect 220084 90312 220136 90364
rect 580080 89360 580132 89412
rect 580540 89360 580592 89412
rect 580540 89224 580592 89276
rect 580724 89224 580776 89276
rect 183468 88952 183520 89004
rect 217324 88952 217376 89004
rect 183376 87592 183428 87644
rect 215944 87592 215996 87644
rect 183468 85484 183520 85536
rect 193956 85484 194008 85536
rect 183468 84124 183520 84176
rect 192484 84124 192536 84176
rect 118608 80724 118660 80776
rect 580908 80724 580960 80776
rect 121092 79976 121144 80028
rect 125416 80248 125468 80300
rect 125232 80044 125284 80096
rect 178592 80656 178644 80708
rect 580816 80656 580868 80708
rect 123852 79976 123904 80028
rect 124956 79908 125008 79960
rect 126106 79908 126158 79960
rect 126198 79908 126250 79960
rect 126382 79908 126434 79960
rect 126842 79908 126894 79960
rect 127210 79908 127262 79960
rect 127302 79908 127354 79960
rect 127486 79908 127538 79960
rect 127578 79908 127630 79960
rect 127670 79908 127722 79960
rect 127854 79908 127906 79960
rect 125830 79840 125882 79892
rect 126014 79840 126066 79892
rect 124772 79772 124824 79824
rect 116584 79704 116636 79756
rect 123576 79704 123628 79756
rect 125738 79772 125790 79824
rect 121184 79636 121236 79688
rect 125416 79636 125468 79688
rect 125600 79636 125652 79688
rect 125692 79636 125744 79688
rect 125968 79636 126020 79688
rect 126290 79840 126342 79892
rect 126244 79704 126296 79756
rect 126336 79704 126388 79756
rect 127026 79772 127078 79824
rect 127578 79772 127630 79824
rect 127256 79704 127308 79756
rect 126888 79636 126940 79688
rect 126980 79636 127032 79688
rect 127164 79636 127216 79688
rect 127946 79840 127998 79892
rect 128130 79908 128182 79960
rect 128590 79908 128642 79960
rect 128774 79908 128826 79960
rect 128866 79908 128918 79960
rect 128958 79908 129010 79960
rect 129234 79908 129286 79960
rect 130154 79908 130206 79960
rect 130246 79908 130298 79960
rect 130338 79908 130390 79960
rect 130430 79908 130482 79960
rect 128406 79772 128458 79824
rect 128636 79772 128688 79824
rect 128728 79772 128780 79824
rect 127900 79704 127952 79756
rect 127992 79704 128044 79756
rect 128084 79704 128136 79756
rect 128820 79704 128872 79756
rect 128360 79636 128412 79688
rect 128452 79636 128504 79688
rect 86224 79568 86276 79620
rect 115296 79432 115348 79484
rect 71780 79364 71832 79416
rect 3976 79296 4028 79348
rect 126060 79568 126112 79620
rect 126152 79568 126204 79620
rect 129142 79840 129194 79892
rect 129786 79840 129838 79892
rect 129602 79772 129654 79824
rect 129188 79636 129240 79688
rect 129556 79636 129608 79688
rect 129280 79568 129332 79620
rect 129464 79568 129516 79620
rect 130200 79704 130252 79756
rect 130292 79704 130344 79756
rect 128912 79500 128964 79552
rect 129096 79500 129148 79552
rect 129740 79500 129792 79552
rect 125508 79432 125560 79484
rect 130890 79908 130942 79960
rect 131718 79908 131770 79960
rect 131994 79908 132046 79960
rect 132270 79908 132322 79960
rect 130706 79772 130758 79824
rect 130660 79636 130712 79688
rect 130568 79568 130620 79620
rect 131074 79840 131126 79892
rect 131028 79704 131080 79756
rect 131856 79636 131908 79688
rect 131304 79568 131356 79620
rect 132316 79704 132368 79756
rect 130844 79500 130896 79552
rect 132224 79500 132276 79552
rect 130936 79432 130988 79484
rect 132914 79908 132966 79960
rect 133190 79908 133242 79960
rect 133926 79908 133978 79960
rect 132868 79636 132920 79688
rect 132960 79568 133012 79620
rect 133742 79840 133794 79892
rect 134662 79908 134714 79960
rect 134846 79908 134898 79960
rect 135122 79908 135174 79960
rect 135398 79908 135450 79960
rect 135582 79908 135634 79960
rect 135950 79908 136002 79960
rect 137238 79908 137290 79960
rect 137606 79908 137658 79960
rect 134202 79840 134254 79892
rect 133972 79772 134024 79824
rect 134708 79772 134760 79824
rect 133512 79568 133564 79620
rect 133788 79568 133840 79620
rect 133328 79500 133380 79552
rect 135306 79840 135358 79892
rect 135352 79636 135404 79688
rect 135260 79500 135312 79552
rect 135766 79840 135818 79892
rect 136042 79840 136094 79892
rect 136686 79840 136738 79892
rect 136870 79840 136922 79892
rect 135720 79704 135772 79756
rect 135536 79500 135588 79552
rect 129096 79364 129148 79416
rect 129832 79364 129884 79416
rect 130108 79364 130160 79416
rect 134800 79432 134852 79484
rect 132776 79364 132828 79416
rect 133880 79364 133932 79416
rect 135996 79364 136048 79416
rect 136824 79636 136876 79688
rect 137008 79568 137060 79620
rect 138526 79908 138578 79960
rect 138710 79908 138762 79960
rect 138894 79908 138946 79960
rect 139078 79908 139130 79960
rect 139446 79908 139498 79960
rect 138342 79840 138394 79892
rect 138572 79772 138624 79824
rect 138664 79772 138716 79824
rect 138802 79772 138854 79824
rect 139170 79840 139222 79892
rect 139032 79704 139084 79756
rect 138756 79636 138808 79688
rect 138848 79636 138900 79688
rect 137836 79568 137888 79620
rect 138204 79568 138256 79620
rect 138940 79568 138992 79620
rect 139906 79908 139958 79960
rect 140366 79908 140418 79960
rect 139492 79636 139544 79688
rect 140090 79840 140142 79892
rect 140274 79840 140326 79892
rect 137468 79500 137520 79552
rect 139676 79500 139728 79552
rect 140320 79500 140372 79552
rect 140504 79500 140556 79552
rect 141286 79908 141338 79960
rect 141562 79908 141614 79960
rect 140918 79840 140970 79892
rect 141010 79840 141062 79892
rect 141102 79840 141154 79892
rect 141470 79840 141522 79892
rect 141746 79840 141798 79892
rect 140964 79636 141016 79688
rect 141516 79704 141568 79756
rect 141148 79568 141200 79620
rect 140964 79500 141016 79552
rect 140044 79432 140096 79484
rect 141332 79568 141384 79620
rect 141700 79500 141752 79552
rect 142482 79908 142534 79960
rect 142574 79908 142626 79960
rect 142758 79908 142810 79960
rect 142850 79908 142902 79960
rect 142942 79908 142994 79960
rect 143034 79908 143086 79960
rect 144138 79908 144190 79960
rect 144230 79908 144282 79960
rect 144322 79908 144374 79960
rect 144414 79908 144466 79960
rect 144598 79908 144650 79960
rect 144690 79908 144742 79960
rect 142206 79840 142258 79892
rect 142528 79704 142580 79756
rect 142252 79568 142304 79620
rect 142344 79500 142396 79552
rect 142712 79568 142764 79620
rect 141884 79432 141936 79484
rect 142160 79432 142212 79484
rect 143862 79840 143914 79892
rect 143310 79772 143362 79824
rect 143402 79772 143454 79824
rect 143586 79772 143638 79824
rect 143678 79772 143730 79824
rect 143264 79636 143316 79688
rect 143540 79636 143592 79688
rect 143080 79568 143132 79620
rect 143448 79568 143500 79620
rect 143954 79772 144006 79824
rect 144000 79636 144052 79688
rect 144184 79636 144236 79688
rect 143356 79500 143408 79552
rect 144092 79568 144144 79620
rect 143724 79500 143776 79552
rect 143816 79432 143868 79484
rect 144368 79432 144420 79484
rect 144736 79568 144788 79620
rect 145702 79908 145754 79960
rect 145794 79908 145846 79960
rect 146254 79908 146306 79960
rect 146346 79908 146398 79960
rect 145150 79840 145202 79892
rect 145242 79840 145294 79892
rect 144920 79500 144972 79552
rect 145748 79772 145800 79824
rect 146438 79840 146490 79892
rect 146300 79704 146352 79756
rect 145288 79636 145340 79688
rect 146116 79636 146168 79688
rect 146392 79568 146444 79620
rect 147174 79908 147226 79960
rect 147358 79908 147410 79960
rect 147450 79908 147502 79960
rect 147542 79908 147594 79960
rect 147634 79908 147686 79960
rect 146990 79840 147042 79892
rect 146806 79772 146858 79824
rect 146852 79636 146904 79688
rect 147496 79704 147548 79756
rect 147312 79636 147364 79688
rect 147404 79636 147456 79688
rect 146668 79568 146720 79620
rect 146944 79568 146996 79620
rect 148278 79840 148330 79892
rect 148370 79840 148422 79892
rect 147910 79772 147962 79824
rect 148324 79704 148376 79756
rect 149198 79908 149250 79960
rect 149290 79908 149342 79960
rect 149566 79908 149618 79960
rect 148968 79636 149020 79688
rect 148140 79568 148192 79620
rect 147220 79500 147272 79552
rect 147680 79500 147732 79552
rect 149382 79840 149434 79892
rect 149474 79840 149526 79892
rect 149842 79840 149894 79892
rect 149520 79636 149572 79688
rect 149244 79568 149296 79620
rect 149428 79500 149480 79552
rect 148508 79432 148560 79484
rect 149060 79364 149112 79416
rect 149796 79636 149848 79688
rect 149980 79568 150032 79620
rect 151130 79908 151182 79960
rect 151498 79908 151550 79960
rect 151590 79908 151642 79960
rect 151958 79908 152010 79960
rect 150256 79568 150308 79620
rect 150670 79840 150722 79892
rect 150854 79840 150906 79892
rect 150440 79500 150492 79552
rect 150624 79500 150676 79552
rect 151222 79840 151274 79892
rect 151314 79840 151366 79892
rect 151268 79704 151320 79756
rect 151360 79568 151412 79620
rect 152234 79840 152286 79892
rect 151544 79772 151596 79824
rect 151866 79772 151918 79824
rect 151636 79704 151688 79756
rect 152004 79636 152056 79688
rect 151912 79568 151964 79620
rect 151268 79432 151320 79484
rect 152096 79364 152148 79416
rect 123576 79296 123628 79348
rect 125600 79160 125652 79212
rect 127624 79160 127676 79212
rect 128084 79160 128136 79212
rect 129648 79228 129700 79280
rect 133512 79228 133564 79280
rect 133880 79228 133932 79280
rect 145472 79160 145524 79212
rect 151912 79296 151964 79348
rect 152510 79908 152562 79960
rect 152372 79704 152424 79756
rect 152280 79636 152332 79688
rect 152694 79908 152746 79960
rect 152602 79840 152654 79892
rect 152970 79772 153022 79824
rect 152648 79704 152700 79756
rect 152556 79636 152608 79688
rect 153338 79908 153390 79960
rect 153522 79908 153574 79960
rect 153706 79908 153758 79960
rect 154902 79908 154954 79960
rect 155454 79908 155506 79960
rect 155822 79908 155874 79960
rect 155914 79908 155966 79960
rect 156282 79908 156334 79960
rect 156374 79908 156426 79960
rect 157018 79908 157070 79960
rect 153476 79568 153528 79620
rect 153890 79840 153942 79892
rect 154166 79840 154218 79892
rect 154718 79840 154770 79892
rect 153660 79636 153712 79688
rect 153844 79636 153896 79688
rect 154028 79568 154080 79620
rect 154304 79568 154356 79620
rect 154580 79568 154632 79620
rect 152832 79500 152884 79552
rect 153016 79500 153068 79552
rect 153292 79500 153344 79552
rect 155132 79500 155184 79552
rect 155408 79500 155460 79552
rect 155868 79772 155920 79824
rect 156466 79840 156518 79892
rect 157294 79840 157346 79892
rect 157386 79840 157438 79892
rect 156558 79772 156610 79824
rect 156742 79772 156794 79824
rect 157064 79772 157116 79824
rect 156512 79636 156564 79688
rect 156328 79568 156380 79620
rect 156420 79568 156472 79620
rect 152924 79432 152976 79484
rect 152464 79364 152516 79416
rect 155684 79364 155736 79416
rect 153108 79296 153160 79348
rect 154948 79296 155000 79348
rect 156420 79432 156472 79484
rect 157156 79636 157208 79688
rect 157340 79636 157392 79688
rect 157570 79908 157622 79960
rect 157662 79840 157714 79892
rect 157754 79840 157806 79892
rect 157432 79568 157484 79620
rect 158214 79908 158266 79960
rect 158122 79840 158174 79892
rect 158168 79704 158220 79756
rect 158490 79840 158542 79892
rect 158582 79840 158634 79892
rect 158444 79704 158496 79756
rect 158260 79636 158312 79688
rect 158352 79636 158404 79688
rect 158536 79636 158588 79688
rect 156972 79500 157024 79552
rect 157248 79500 157300 79552
rect 157708 79500 157760 79552
rect 157616 79432 157668 79484
rect 156972 79364 157024 79416
rect 174636 80588 174688 80640
rect 178040 80588 178092 80640
rect 580448 80588 580500 80640
rect 175740 80520 175792 80572
rect 580356 80520 580408 80572
rect 175924 80452 175976 80504
rect 158766 79908 158818 79960
rect 158858 79908 158910 79960
rect 159042 79908 159094 79960
rect 159318 79908 159370 79960
rect 159686 79908 159738 79960
rect 159778 79908 159830 79960
rect 160054 79908 160106 79960
rect 160146 79908 160198 79960
rect 160238 79908 160290 79960
rect 160330 79908 160382 79960
rect 160422 79908 160474 79960
rect 160606 79908 160658 79960
rect 160698 79908 160750 79960
rect 158812 79772 158864 79824
rect 158950 79772 159002 79824
rect 158904 79636 158956 79688
rect 159226 79840 159278 79892
rect 159594 79840 159646 79892
rect 159272 79568 159324 79620
rect 159180 79500 159232 79552
rect 159640 79704 159692 79756
rect 159548 79568 159600 79620
rect 159824 79500 159876 79552
rect 160192 79772 160244 79824
rect 160284 79772 160336 79824
rect 160606 79772 160658 79824
rect 160468 79636 160520 79688
rect 160560 79568 160612 79620
rect 161158 79908 161210 79960
rect 161066 79840 161118 79892
rect 160974 79772 161026 79824
rect 161342 79840 161394 79892
rect 161618 79840 161670 79892
rect 161894 79840 161946 79892
rect 162170 79840 162222 79892
rect 161204 79772 161256 79824
rect 161112 79704 161164 79756
rect 161020 79636 161072 79688
rect 161940 79636 161992 79688
rect 162032 79636 162084 79688
rect 160928 79568 160980 79620
rect 162262 79772 162314 79824
rect 161388 79500 161440 79552
rect 159732 79432 159784 79484
rect 159916 79432 159968 79484
rect 162124 79364 162176 79416
rect 162538 79908 162590 79960
rect 163274 79908 163326 79960
rect 163918 79908 163970 79960
rect 162722 79840 162774 79892
rect 163090 79840 163142 79892
rect 163182 79840 163234 79892
rect 162584 79772 162636 79824
rect 162676 79704 162728 79756
rect 163044 79704 163096 79756
rect 163136 79704 163188 79756
rect 162952 79636 163004 79688
rect 163734 79840 163786 79892
rect 163826 79840 163878 79892
rect 163550 79772 163602 79824
rect 163872 79568 163924 79620
rect 163504 79500 163556 79552
rect 163688 79500 163740 79552
rect 162860 79432 162912 79484
rect 164562 79908 164614 79960
rect 165022 79840 165074 79892
rect 164838 79772 164890 79824
rect 164148 79636 164200 79688
rect 165206 79908 165258 79960
rect 165942 79908 165994 79960
rect 166402 79908 166454 79960
rect 165666 79840 165718 79892
rect 166126 79840 166178 79892
rect 165252 79772 165304 79824
rect 164056 79568 164108 79620
rect 164792 79568 164844 79620
rect 165528 79568 165580 79620
rect 165712 79568 165764 79620
rect 166264 79568 166316 79620
rect 167506 79908 167558 79960
rect 167782 79908 167834 79960
rect 167046 79840 167098 79892
rect 166816 79636 166868 79688
rect 166632 79500 166684 79552
rect 167368 79568 167420 79620
rect 168334 79908 168386 79960
rect 168426 79840 168478 79892
rect 168288 79772 168340 79824
rect 168380 79704 168432 79756
rect 168886 79908 168938 79960
rect 169070 79908 169122 79960
rect 169438 79908 169490 79960
rect 169254 79840 169306 79892
rect 169024 79704 169076 79756
rect 168932 79636 168984 79688
rect 168840 79568 168892 79620
rect 164884 79432 164936 79484
rect 163964 79364 164016 79416
rect 164240 79364 164292 79416
rect 166908 79364 166960 79416
rect 164884 79296 164936 79348
rect 165528 79296 165580 79348
rect 167460 79296 167512 79348
rect 168656 79364 168708 79416
rect 169806 79772 169858 79824
rect 169208 79636 169260 79688
rect 169760 79636 169812 79688
rect 169990 79636 170042 79688
rect 170036 79500 170088 79552
rect 169300 79364 169352 79416
rect 170634 79908 170686 79960
rect 170312 79364 170364 79416
rect 170726 79840 170778 79892
rect 180156 80384 180208 80436
rect 231860 80248 231912 80300
rect 174452 80180 174504 80232
rect 249800 80180 249852 80232
rect 171094 79908 171146 79960
rect 175740 80112 175792 80164
rect 175832 80112 175884 80164
rect 284300 80112 284352 80164
rect 175096 80044 175148 80096
rect 175924 80044 175976 80096
rect 426440 80044 426492 80096
rect 171554 79908 171606 79960
rect 171830 79908 171882 79960
rect 171922 79908 171974 79960
rect 172106 79908 172158 79960
rect 172198 79908 172250 79960
rect 172566 79908 172618 79960
rect 171646 79840 171698 79892
rect 171600 79704 171652 79756
rect 170864 79636 170916 79688
rect 170772 79568 170824 79620
rect 172060 79772 172112 79824
rect 172152 79772 172204 79824
rect 172934 79840 172986 79892
rect 173302 79840 173354 79892
rect 173670 79908 173722 79960
rect 173624 79772 173676 79824
rect 173256 79704 173308 79756
rect 173946 79840 173998 79892
rect 174130 79772 174182 79824
rect 173992 79704 174044 79756
rect 171968 79636 172020 79688
rect 173072 79636 173124 79688
rect 174084 79636 174136 79688
rect 174544 79636 174596 79688
rect 374000 79636 374052 79688
rect 172612 79568 172664 79620
rect 179512 79568 179564 79620
rect 171692 79432 171744 79484
rect 171784 79432 171836 79484
rect 173164 79432 173216 79484
rect 173716 79432 173768 79484
rect 174636 79432 174688 79484
rect 171508 79364 171560 79416
rect 173348 79364 173400 79416
rect 177396 79500 177448 79552
rect 331220 79500 331272 79552
rect 175096 79432 175148 79484
rect 580264 79432 580316 79484
rect 580632 79364 580684 79416
rect 171692 79296 171744 79348
rect 173808 79296 173860 79348
rect 165160 79228 165212 79280
rect 165436 79228 165488 79280
rect 155684 79160 155736 79212
rect 128084 79024 128136 79076
rect 128636 79024 128688 79076
rect 129096 79024 129148 79076
rect 133880 79024 133932 79076
rect 130384 78956 130436 79008
rect 130568 78956 130620 79008
rect 152464 79092 152516 79144
rect 158352 79092 158404 79144
rect 158996 79092 159048 79144
rect 159732 79092 159784 79144
rect 165804 79160 165856 79212
rect 168012 79160 168064 79212
rect 168840 79160 168892 79212
rect 169576 79160 169628 79212
rect 169760 79160 169812 79212
rect 170128 79160 170180 79212
rect 171600 79228 171652 79280
rect 580540 79296 580592 79348
rect 171692 79160 171744 79212
rect 171876 79160 171928 79212
rect 175832 79160 175884 79212
rect 154028 79024 154080 79076
rect 163136 79024 163188 79076
rect 170956 79092 171008 79144
rect 171324 79092 171376 79144
rect 182916 79092 182968 79144
rect 165804 79024 165856 79076
rect 166080 79024 166132 79076
rect 200120 79024 200172 79076
rect 153108 78956 153160 79008
rect 159180 78956 159232 79008
rect 252560 78956 252612 79008
rect 44824 78752 44876 78804
rect 145472 78888 145524 78940
rect 152924 78888 152976 78940
rect 154948 78888 155000 78940
rect 165436 78888 165488 78940
rect 165528 78888 165580 78940
rect 213920 78888 213972 78940
rect 154672 78752 154724 78804
rect 155040 78752 155092 78804
rect 157984 78752 158036 78804
rect 158260 78752 158312 78804
rect 125968 78684 126020 78736
rect 126336 78684 126388 78736
rect 155960 78684 156012 78736
rect 156236 78684 156288 78736
rect 159732 78752 159784 78804
rect 306380 78820 306432 78872
rect 164240 78752 164292 78804
rect 164700 78752 164752 78804
rect 164884 78752 164936 78804
rect 173900 78752 173952 78804
rect 124036 78616 124088 78668
rect 128084 78616 128136 78668
rect 135352 78616 135404 78668
rect 135812 78616 135864 78668
rect 147588 78616 147640 78668
rect 165160 78684 165212 78736
rect 170956 78684 171008 78736
rect 171232 78684 171284 78736
rect 172428 78684 172480 78736
rect 172612 78684 172664 78736
rect 201500 78752 201552 78804
rect 93124 78548 93176 78600
rect 127992 78548 128044 78600
rect 155868 78548 155920 78600
rect 157984 78548 158036 78600
rect 126152 78480 126204 78532
rect 126336 78480 126388 78532
rect 130016 78480 130068 78532
rect 130752 78480 130804 78532
rect 141240 78480 141292 78532
rect 164700 78548 164752 78600
rect 166908 78548 166960 78600
rect 171692 78548 171744 78600
rect 171968 78616 172020 78668
rect 182272 78616 182324 78668
rect 173532 78548 173584 78600
rect 170864 78480 170916 78532
rect 170956 78480 171008 78532
rect 171140 78480 171192 78532
rect 172888 78480 172940 78532
rect 180800 78480 180852 78532
rect 123668 78412 123720 78464
rect 134892 78412 134944 78464
rect 153200 78412 153252 78464
rect 156236 78412 156288 78464
rect 157708 78412 157760 78464
rect 158076 78412 158128 78464
rect 161664 78412 161716 78464
rect 127072 78344 127124 78396
rect 135260 78344 135312 78396
rect 149520 78344 149572 78396
rect 159732 78344 159784 78396
rect 162124 78344 162176 78396
rect 165160 78344 165212 78396
rect 167644 78412 167696 78464
rect 242164 78412 242216 78464
rect 315304 78344 315356 78396
rect 113824 78208 113876 78260
rect 125876 78276 125928 78328
rect 142252 78276 142304 78328
rect 165528 78276 165580 78328
rect 165804 78276 165856 78328
rect 430580 78276 430632 78328
rect 110420 78140 110472 78192
rect 129648 78208 129700 78260
rect 89720 78004 89772 78056
rect 132500 78072 132552 78124
rect 144920 78208 144972 78260
rect 154764 78208 154816 78260
rect 161296 78208 161348 78260
rect 162768 78208 162820 78260
rect 436744 78208 436796 78260
rect 145288 78140 145340 78192
rect 150808 78140 150860 78192
rect 151176 78140 151228 78192
rect 155316 78140 155368 78192
rect 159732 78140 159784 78192
rect 164700 78140 164752 78192
rect 159180 78072 159232 78124
rect 164424 78072 164476 78124
rect 164976 78072 165028 78124
rect 165436 78140 165488 78192
rect 480260 78140 480312 78192
rect 171508 78072 171560 78124
rect 171692 78072 171744 78124
rect 498200 78072 498252 78124
rect 145288 78004 145340 78056
rect 150716 78004 150768 78056
rect 157248 78004 157300 78056
rect 168380 78004 168432 78056
rect 170772 78004 170824 78056
rect 170864 78004 170916 78056
rect 53840 77936 53892 77988
rect 129740 77936 129792 77988
rect 137836 77936 137888 77988
rect 138020 77936 138072 77988
rect 139492 77936 139544 77988
rect 145840 77936 145892 77988
rect 154212 77936 154264 77988
rect 162768 77936 162820 77988
rect 166816 77936 166868 77988
rect 171876 77936 171928 77988
rect 171968 77936 172020 77988
rect 174084 77936 174136 77988
rect 174544 78004 174596 78056
rect 574744 78004 574796 78056
rect 581092 77936 581144 77988
rect 125324 77868 125376 77920
rect 133052 77868 133104 77920
rect 141148 77868 141200 77920
rect 152832 77868 152884 77920
rect 154764 77868 154816 77920
rect 155592 77868 155644 77920
rect 157064 77868 157116 77920
rect 171324 77868 171376 77920
rect 116584 77800 116636 77852
rect 129188 77800 129240 77852
rect 129924 77800 129976 77852
rect 131672 77800 131724 77852
rect 152004 77800 152056 77852
rect 152556 77800 152608 77852
rect 157432 77800 157484 77852
rect 171784 77800 171836 77852
rect 143540 77732 143592 77784
rect 125416 77664 125468 77716
rect 133696 77664 133748 77716
rect 154580 77732 154632 77784
rect 158628 77732 158680 77784
rect 159272 77732 159324 77784
rect 159180 77664 159232 77716
rect 164884 77732 164936 77784
rect 172152 77732 172204 77784
rect 171692 77664 171744 77716
rect 122380 77596 122432 77648
rect 125232 77596 125284 77648
rect 145012 77596 145064 77648
rect 159272 77596 159324 77648
rect 120816 77528 120868 77580
rect 128268 77528 128320 77580
rect 141884 77528 141936 77580
rect 166080 77596 166132 77648
rect 169300 77596 169352 77648
rect 170312 77596 170364 77648
rect 179144 77596 179196 77648
rect 580080 77596 580132 77648
rect 164884 77528 164936 77580
rect 174452 77528 174504 77580
rect 3516 77460 3568 77512
rect 173992 77460 174044 77512
rect 125692 77392 125744 77444
rect 135444 77392 135496 77444
rect 151452 77392 151504 77444
rect 153844 77392 153896 77444
rect 159180 77392 159232 77444
rect 168840 77392 168892 77444
rect 171600 77392 171652 77444
rect 171784 77392 171836 77444
rect 125232 77324 125284 77376
rect 132408 77324 132460 77376
rect 158352 77324 158404 77376
rect 166816 77324 166868 77376
rect 126244 77256 126296 77308
rect 130568 77256 130620 77308
rect 151820 77256 151872 77308
rect 152740 77256 152792 77308
rect 158812 77256 158864 77308
rect 158996 77256 159048 77308
rect 159272 77256 159324 77308
rect 164884 77256 164936 77308
rect 166632 77256 166684 77308
rect 170496 77256 170548 77308
rect 125876 77188 125928 77240
rect 126796 77188 126848 77240
rect 127164 77188 127216 77240
rect 127440 77188 127492 77240
rect 127532 77188 127584 77240
rect 127808 77188 127860 77240
rect 128084 77188 128136 77240
rect 128360 77188 128412 77240
rect 152004 77188 152056 77240
rect 152464 77188 152516 77240
rect 154304 77188 154356 77240
rect 155776 77188 155828 77240
rect 160284 77188 160336 77240
rect 160836 77188 160888 77240
rect 163044 77188 163096 77240
rect 163596 77188 163648 77240
rect 163964 77188 164016 77240
rect 169300 77188 169352 77240
rect 172336 77188 172388 77240
rect 527180 77188 527232 77240
rect 143632 77120 143684 77172
rect 143908 77120 143960 77172
rect 152740 77120 152792 77172
rect 226340 77120 226392 77172
rect 149244 77052 149296 77104
rect 149520 77052 149572 77104
rect 152464 77052 152516 77104
rect 240140 77052 240192 77104
rect 129096 76984 129148 77036
rect 130200 76984 130252 77036
rect 145932 76984 145984 77036
rect 260840 76984 260892 77036
rect 146116 76916 146168 76968
rect 267740 76916 267792 76968
rect 133052 76848 133104 76900
rect 135536 76848 135588 76900
rect 144000 76848 144052 76900
rect 144184 76848 144236 76900
rect 146576 76848 146628 76900
rect 147036 76848 147088 76900
rect 148048 76848 148100 76900
rect 288440 76848 288492 76900
rect 122840 76780 122892 76832
rect 133328 76780 133380 76832
rect 143908 76780 143960 76832
rect 144092 76780 144144 76832
rect 148600 76780 148652 76832
rect 296720 76780 296772 76832
rect 118700 76712 118752 76764
rect 133788 76712 133840 76764
rect 136916 76712 136968 76764
rect 137100 76712 137152 76764
rect 138848 76712 138900 76764
rect 139308 76712 139360 76764
rect 139492 76712 139544 76764
rect 140044 76712 140096 76764
rect 143816 76712 143868 76764
rect 144000 76712 144052 76764
rect 146208 76712 146260 76764
rect 146668 76712 146720 76764
rect 149152 76712 149204 76764
rect 302240 76712 302292 76764
rect 93860 76644 93912 76696
rect 130936 76644 130988 76696
rect 132408 76644 132460 76696
rect 140504 76644 140556 76696
rect 142896 76644 142948 76696
rect 70400 76576 70452 76628
rect 131028 76576 131080 76628
rect 131764 76576 131816 76628
rect 132040 76576 132092 76628
rect 132684 76576 132736 76628
rect 133236 76576 133288 76628
rect 133420 76576 133472 76628
rect 133696 76576 133748 76628
rect 135812 76576 135864 76628
rect 136456 76576 136508 76628
rect 138296 76576 138348 76628
rect 138848 76576 138900 76628
rect 140780 76576 140832 76628
rect 141700 76576 141752 76628
rect 143816 76576 143868 76628
rect 144460 76576 144512 76628
rect 145012 76576 145064 76628
rect 145380 76576 145432 76628
rect 146392 76576 146444 76628
rect 146668 76576 146720 76628
rect 148048 76576 148100 76628
rect 148324 76576 148376 76628
rect 149336 76644 149388 76696
rect 149888 76644 149940 76696
rect 150256 76644 150308 76696
rect 152464 76644 152516 76696
rect 154396 76644 154448 76696
rect 356060 76644 356112 76696
rect 152740 76576 152792 76628
rect 159272 76576 159324 76628
rect 159548 76576 159600 76628
rect 160192 76576 160244 76628
rect 160376 76576 160428 76628
rect 160468 76576 160520 76628
rect 160652 76576 160704 76628
rect 161572 76576 161624 76628
rect 162216 76576 162268 76628
rect 163044 76576 163096 76628
rect 163504 76576 163556 76628
rect 165804 76576 165856 76628
rect 166356 76576 166408 76628
rect 166448 76576 166500 76628
rect 166632 76576 166684 76628
rect 167644 76576 167696 76628
rect 167828 76576 167880 76628
rect 168656 76576 168708 76628
rect 169392 76576 169444 76628
rect 69020 76508 69072 76560
rect 131120 76508 131172 76560
rect 139584 76508 139636 76560
rect 139952 76508 140004 76560
rect 141240 76508 141292 76560
rect 141516 76508 141568 76560
rect 142252 76508 142304 76560
rect 142804 76508 142856 76560
rect 146852 76508 146904 76560
rect 147128 76508 147180 76560
rect 149244 76508 149296 76560
rect 149704 76508 149756 76560
rect 152464 76508 152516 76560
rect 152924 76508 152976 76560
rect 161664 76508 161716 76560
rect 162308 76508 162360 76560
rect 164332 76508 164384 76560
rect 164792 76508 164844 76560
rect 168380 76508 168432 76560
rect 169116 76508 169168 76560
rect 169300 76508 169352 76560
rect 171784 76576 171836 76628
rect 172152 76576 172204 76628
rect 557540 76576 557592 76628
rect 170312 76508 170364 76560
rect 558920 76508 558972 76560
rect 131028 76440 131080 76492
rect 132592 76440 132644 76492
rect 137928 76440 137980 76492
rect 138664 76440 138716 76492
rect 139768 76440 139820 76492
rect 182180 76440 182232 76492
rect 124864 76372 124916 76424
rect 131580 76372 131632 76424
rect 145380 76372 145432 76424
rect 145656 76372 145708 76424
rect 145840 76372 145892 76424
rect 178040 76372 178092 76424
rect 139768 76304 139820 76356
rect 140228 76304 140280 76356
rect 147772 76304 147824 76356
rect 148324 76304 148376 76356
rect 150900 76304 150952 76356
rect 151452 76304 151504 76356
rect 160376 76304 160428 76356
rect 160744 76304 160796 76356
rect 161480 76304 161532 76356
rect 167828 76304 167880 76356
rect 168472 76304 168524 76356
rect 168840 76304 168892 76356
rect 171508 76304 171560 76356
rect 195980 76304 196032 76356
rect 125140 76236 125192 76288
rect 126704 76236 126756 76288
rect 131580 76236 131632 76288
rect 131948 76236 132000 76288
rect 135628 76236 135680 76288
rect 136640 76236 136692 76288
rect 164148 76236 164200 76288
rect 164424 76236 164476 76288
rect 167000 76236 167052 76288
rect 167920 76236 167972 76288
rect 160468 76168 160520 76220
rect 161020 76168 161072 76220
rect 168472 76168 168524 76220
rect 169024 76168 169076 76220
rect 128728 76100 128780 76152
rect 129464 76100 129516 76152
rect 136640 76100 136692 76152
rect 137744 76100 137796 76152
rect 144920 76100 144972 76152
rect 146024 76100 146076 76152
rect 159456 76100 159508 76152
rect 159824 76100 159876 76152
rect 160744 76100 160796 76152
rect 160928 76100 160980 76152
rect 165712 76100 165764 76152
rect 166264 76100 166316 76152
rect 125048 76032 125100 76084
rect 126980 76032 127032 76084
rect 129740 76032 129792 76084
rect 135904 76032 135956 76084
rect 131488 75964 131540 76016
rect 132132 75964 132184 76016
rect 163136 75964 163188 76016
rect 163872 75964 163924 76016
rect 137376 75896 137428 75948
rect 144460 75896 144512 75948
rect 153384 75896 153436 75948
rect 153568 75896 153620 75948
rect 170956 75896 171008 75948
rect 173348 75896 173400 75948
rect 134064 75828 134116 75880
rect 134708 75828 134760 75880
rect 130384 75760 130436 75812
rect 133052 75760 133104 75812
rect 129188 75692 129240 75744
rect 129556 75692 129608 75744
rect 159640 75692 159692 75744
rect 164884 75692 164936 75744
rect 155040 75624 155092 75676
rect 155316 75624 155368 75676
rect 157340 75624 157392 75676
rect 157892 75624 157944 75676
rect 125784 75488 125836 75540
rect 126612 75488 126664 75540
rect 128544 75488 128596 75540
rect 129924 75488 129976 75540
rect 135536 75488 135588 75540
rect 136272 75488 136324 75540
rect 142528 75488 142580 75540
rect 142712 75488 142764 75540
rect 152832 75488 152884 75540
rect 167460 75556 167512 75608
rect 167828 75556 167880 75608
rect 197360 75488 197412 75540
rect 123576 75420 123628 75472
rect 130108 75420 130160 75472
rect 153660 75420 153712 75472
rect 155592 75420 155644 75472
rect 167092 75420 167144 75472
rect 167460 75420 167512 75472
rect 171140 75420 171192 75472
rect 358820 75420 358872 75472
rect 107660 75352 107712 75404
rect 132224 75352 132276 75404
rect 142528 75352 142580 75404
rect 143080 75352 143132 75404
rect 157340 75352 157392 75404
rect 157708 75352 157760 75404
rect 164884 75352 164936 75404
rect 438860 75352 438912 75404
rect 51080 75284 51132 75336
rect 125508 75284 125560 75336
rect 49700 75216 49752 75268
rect 129280 75284 129332 75336
rect 134340 75284 134392 75336
rect 134616 75284 134668 75336
rect 150716 75284 150768 75336
rect 151084 75284 151136 75336
rect 154580 75284 154632 75336
rect 155500 75284 155552 75336
rect 156052 75284 156104 75336
rect 156604 75284 156656 75336
rect 163780 75284 163832 75336
rect 489920 75284 489972 75336
rect 150808 75216 150860 75268
rect 151268 75216 151320 75268
rect 154948 75216 155000 75268
rect 155224 75216 155276 75268
rect 156328 75216 156380 75268
rect 156512 75216 156564 75268
rect 157708 75216 157760 75268
rect 158168 75216 158220 75268
rect 167828 75216 167880 75268
rect 506480 75216 506532 75268
rect 46940 75148 46992 75200
rect 134156 75148 134208 75200
rect 135168 75148 135220 75200
rect 150900 75148 150952 75200
rect 151360 75148 151412 75200
rect 155040 75148 155092 75200
rect 155408 75148 155460 75200
rect 156052 75148 156104 75200
rect 156972 75148 157024 75200
rect 157524 75148 157576 75200
rect 158260 75148 158312 75200
rect 168012 75148 168064 75200
rect 517520 75148 517572 75200
rect 147772 75080 147824 75132
rect 148416 75080 148468 75132
rect 152188 75080 152240 75132
rect 152648 75080 152700 75132
rect 153568 75080 153620 75132
rect 154120 75080 154172 75132
rect 169944 75080 169996 75132
rect 170220 75080 170272 75132
rect 124036 75012 124088 75064
rect 135444 75012 135496 75064
rect 136180 75012 136232 75064
rect 156236 75012 156288 75064
rect 156788 75012 156840 75064
rect 163228 75012 163280 75064
rect 163688 75012 163740 75064
rect 156144 74944 156196 74996
rect 156880 74944 156932 74996
rect 136732 74604 136784 74656
rect 137008 74604 137060 74656
rect 139492 74604 139544 74656
rect 140320 74604 140372 74656
rect 138480 74536 138532 74588
rect 138756 74536 138808 74588
rect 144092 74536 144144 74588
rect 144368 74536 144420 74588
rect 171232 74468 171284 74520
rect 171692 74468 171744 74520
rect 149152 74400 149204 74452
rect 150072 74400 150124 74452
rect 145472 74264 145524 74316
rect 145748 74264 145800 74316
rect 141792 74128 141844 74180
rect 209780 74128 209832 74180
rect 146300 74060 146352 74112
rect 216680 74060 216732 74112
rect 119344 73992 119396 74044
rect 130476 73992 130528 74044
rect 131120 73992 131172 74044
rect 134984 73992 135036 74044
rect 143356 73992 143408 74044
rect 223580 73992 223632 74044
rect 93952 73924 94004 73976
rect 131028 73924 131080 73976
rect 147220 73924 147272 73976
rect 251180 73924 251232 73976
rect 69112 73856 69164 73908
rect 130844 73856 130896 73908
rect 137468 73856 137520 73908
rect 139216 73856 139268 73908
rect 153292 73856 153344 73908
rect 347780 73856 347832 73908
rect 30380 73788 30432 73840
rect 127900 73788 127952 73840
rect 141332 73788 141384 73840
rect 141608 73788 141660 73840
rect 157984 73788 158036 73840
rect 390560 73788 390612 73840
rect 136732 73720 136784 73772
rect 137560 73720 137612 73772
rect 138020 73244 138072 73296
rect 142988 73244 143040 73296
rect 171048 73108 171100 73160
rect 580172 73108 580224 73160
rect 150072 72768 150124 72820
rect 307760 72768 307812 72820
rect 122288 72700 122340 72752
rect 130568 72700 130620 72752
rect 149704 72700 149756 72752
rect 311900 72700 311952 72752
rect 114560 72632 114612 72684
rect 134524 72632 134576 72684
rect 151452 72632 151504 72684
rect 325700 72632 325752 72684
rect 96620 72564 96672 72616
rect 133144 72564 133196 72616
rect 151728 72564 151780 72616
rect 332600 72564 332652 72616
rect 85580 72496 85632 72548
rect 132316 72496 132368 72548
rect 154488 72496 154540 72548
rect 340880 72496 340932 72548
rect 26240 72428 26292 72480
rect 127808 72428 127860 72480
rect 152464 72428 152516 72480
rect 343640 72428 343692 72480
rect 166632 72360 166684 72412
rect 173256 72360 173308 72412
rect 132592 71680 132644 71732
rect 135352 71680 135404 71732
rect 3424 71612 3476 71664
rect 9036 71612 9088 71664
rect 121460 71408 121512 71460
rect 134892 71408 134944 71460
rect 100760 71340 100812 71392
rect 133696 71340 133748 71392
rect 82820 71272 82872 71324
rect 131304 71272 131356 71324
rect 155316 71272 155368 71324
rect 382280 71272 382332 71324
rect 48320 71204 48372 71256
rect 129372 71204 129424 71256
rect 157892 71204 157944 71256
rect 408500 71204 408552 71256
rect 29000 71136 29052 71188
rect 128084 71136 128136 71188
rect 165252 71136 165304 71188
rect 500960 71136 501012 71188
rect 16580 71068 16632 71120
rect 126612 71068 126664 71120
rect 164884 71068 164936 71120
rect 507860 71068 507912 71120
rect 11060 71000 11112 71052
rect 126520 71000 126572 71052
rect 139308 71000 139360 71052
rect 165068 71000 165120 71052
rect 166172 71000 166224 71052
rect 523040 71000 523092 71052
rect 141516 69980 141568 70032
rect 209872 69980 209924 70032
rect 159364 69912 159416 69964
rect 431960 69912 432012 69964
rect 103520 69844 103572 69896
rect 133052 69844 133104 69896
rect 159272 69844 159324 69896
rect 437480 69844 437532 69896
rect 78680 69776 78732 69828
rect 131856 69776 131908 69828
rect 160836 69776 160888 69828
rect 447140 69776 447192 69828
rect 60740 69708 60792 69760
rect 129096 69708 129148 69760
rect 167920 69708 167972 69760
rect 536840 69708 536892 69760
rect 44180 69640 44232 69692
rect 128912 69640 128964 69692
rect 169484 69640 169536 69692
rect 564440 69640 564492 69692
rect 137284 68960 137336 69012
rect 138756 68960 138808 69012
rect 138664 68892 138716 68944
rect 140136 68892 140188 68944
rect 141424 68552 141476 68604
rect 202880 68552 202932 68604
rect 144276 68484 144328 68536
rect 238760 68484 238812 68536
rect 157156 68416 157208 68468
rect 320180 68416 320232 68468
rect 162124 68348 162176 68400
rect 467840 68348 467892 68400
rect 115940 68280 115992 68332
rect 134248 68280 134300 68332
rect 169024 68280 169076 68332
rect 561680 68280 561732 68332
rect 145564 67056 145616 67108
rect 256700 67056 256752 67108
rect 156696 66988 156748 67040
rect 396080 66988 396132 67040
rect 167736 66920 167788 66972
rect 539600 66920 539652 66972
rect 33140 66852 33192 66904
rect 127532 66852 127584 66904
rect 167644 66852 167696 66904
rect 543740 66852 543792 66904
rect 138572 66172 138624 66224
rect 140228 66172 140280 66224
rect 142712 65628 142764 65680
rect 218060 65628 218112 65680
rect 144184 65560 144236 65612
rect 234620 65560 234672 65612
rect 155776 65492 155828 65544
rect 367100 65492 367152 65544
rect 141332 64404 141384 64456
rect 207020 64404 207072 64456
rect 142620 64336 142672 64388
rect 220820 64336 220872 64388
rect 153660 64268 153712 64320
rect 362960 64268 363012 64320
rect 158352 64200 158404 64252
rect 374092 64200 374144 64252
rect 155132 64132 155184 64184
rect 376760 64132 376812 64184
rect 144092 62908 144144 62960
rect 242900 62908 242952 62960
rect 151084 62840 151136 62892
rect 324320 62840 324372 62892
rect 137192 62772 137244 62824
rect 144184 62772 144236 62824
rect 163596 62772 163648 62824
rect 481640 62772 481692 62824
rect 142528 61616 142580 61668
rect 224960 61616 225012 61668
rect 162308 61548 162360 61600
rect 368480 61548 368532 61600
rect 156604 61480 156656 61532
rect 390652 61480 390704 61532
rect 157892 61412 157944 61464
rect 412640 61412 412692 61464
rect 102140 61344 102192 61396
rect 125416 61344 125468 61396
rect 159180 61344 159232 61396
rect 440240 61344 440292 61396
rect 137100 60664 137152 60716
rect 142804 60664 142856 60716
rect 183008 60664 183060 60716
rect 580172 60664 580224 60716
rect 140044 60324 140096 60376
rect 180800 60324 180852 60376
rect 120080 60256 120132 60308
rect 123668 60256 123720 60308
rect 145472 60256 145524 60308
rect 259460 60256 259512 60308
rect 150992 60188 151044 60240
rect 327080 60188 327132 60240
rect 160744 60120 160796 60172
rect 444380 60120 444432 60172
rect 163504 60052 163556 60104
rect 481732 60052 481784 60104
rect 164792 59984 164844 60036
rect 498292 59984 498344 60036
rect 3056 59304 3108 59356
rect 181536 59304 181588 59356
rect 149612 58760 149664 58812
rect 309140 58760 309192 58812
rect 152464 58692 152516 58744
rect 340972 58692 341024 58744
rect 155040 58624 155092 58676
rect 383660 58624 383712 58676
rect 137008 57876 137060 57928
rect 140044 57876 140096 57928
rect 139952 57536 140004 57588
rect 179420 57536 179472 57588
rect 152372 57468 152424 57520
rect 345020 57468 345072 57520
rect 156512 57400 156564 57452
rect 394700 57400 394752 57452
rect 159088 57332 159140 57384
rect 433340 57332 433392 57384
rect 164700 57264 164752 57316
rect 505100 57264 505152 57316
rect 95240 57196 95292 57248
rect 125324 57196 125376 57248
rect 168932 57196 168984 57248
rect 564532 57196 564584 57248
rect 153568 55904 153620 55956
rect 365720 55904 365772 55956
rect 88340 55836 88392 55888
rect 125232 55836 125284 55888
rect 157800 55836 157852 55888
rect 415400 55836 415452 55888
rect 150900 54748 150952 54800
rect 331220 54748 331272 54800
rect 154948 54680 155000 54732
rect 380900 54680 380952 54732
rect 156420 54612 156472 54664
rect 398840 54612 398892 54664
rect 160652 54544 160704 54596
rect 448520 54544 448572 54596
rect 163412 54476 163464 54528
rect 487160 54476 487212 54528
rect 157708 53320 157760 53372
rect 419540 53320 419592 53372
rect 160560 53252 160612 53304
rect 451280 53252 451332 53304
rect 167552 53184 167604 53236
rect 538220 53184 538272 53236
rect 168840 53116 168892 53168
rect 552020 53116 552072 53168
rect 170128 53048 170180 53100
rect 571340 53048 571392 53100
rect 141240 51824 141292 51876
rect 204260 51824 204312 51876
rect 166080 51756 166132 51808
rect 527180 51756 527232 51808
rect 13820 51688 13872 51740
rect 125140 51688 125192 51740
rect 138480 51688 138532 51740
rect 166264 51688 166316 51740
rect 167460 51688 167512 51740
rect 534080 51688 534132 51740
rect 144000 50600 144052 50652
rect 233240 50600 233292 50652
rect 165988 50532 166040 50584
rect 520280 50532 520332 50584
rect 165804 50464 165856 50516
rect 523132 50464 523184 50516
rect 170772 50396 170824 50448
rect 550640 50396 550692 50448
rect 170036 50328 170088 50380
rect 569960 50328 570012 50380
rect 139860 49240 139912 49292
rect 183560 49240 183612 49292
rect 153476 49172 153528 49224
rect 357440 49172 357492 49224
rect 159732 49104 159784 49156
rect 382372 49104 382424 49156
rect 171600 49036 171652 49088
rect 432052 49036 432104 49088
rect 138388 48968 138440 49020
rect 165804 48968 165856 49020
rect 165896 48968 165948 49020
rect 516140 48968 516192 49020
rect 142436 47676 142488 47728
rect 215300 47676 215352 47728
rect 164608 47608 164660 47660
rect 502340 47608 502392 47660
rect 168656 47540 168708 47592
rect 563060 47540 563112 47592
rect 118516 46860 118568 46912
rect 580172 46860 580224 46912
rect 139768 46316 139820 46368
rect 187700 46316 187752 46368
rect 143908 46248 143960 46300
rect 236000 46248 236052 46300
rect 158996 46180 159048 46232
rect 427820 46180 427872 46232
rect 3424 45500 3476 45552
rect 173992 45500 174044 45552
rect 141148 45024 141200 45076
rect 208400 45024 208452 45076
rect 152280 44956 152332 45008
rect 339500 44956 339552 45008
rect 138296 44888 138348 44940
rect 168656 44888 168708 44940
rect 171692 44888 171744 44940
rect 425060 44888 425112 44940
rect 81440 44820 81492 44872
rect 131580 44820 131632 44872
rect 163320 44820 163372 44872
rect 485780 44820 485832 44872
rect 139676 43528 139728 43580
rect 185032 43528 185084 43580
rect 152188 43460 152240 43512
rect 349160 43460 349212 43512
rect 168748 43392 168800 43444
rect 556160 43392 556212 43444
rect 142344 42168 142396 42220
rect 218152 42168 218204 42220
rect 148324 42100 148376 42152
rect 285680 42100 285732 42152
rect 150808 42032 150860 42084
rect 328460 42032 328512 42084
rect 145380 37952 145432 38004
rect 258080 37952 258132 38004
rect 45560 37884 45612 37936
rect 116584 37884 116636 37936
rect 152096 37884 152148 37936
rect 338120 37884 338172 37936
rect 7564 36524 7616 36576
rect 124220 36524 124272 36576
rect 166632 36524 166684 36576
rect 418160 36524 418212 36576
rect 148232 35368 148284 35420
rect 291200 35368 291252 35420
rect 149520 35300 149572 35352
rect 305000 35300 305052 35352
rect 160928 35232 160980 35284
rect 375380 35232 375432 35284
rect 38660 35164 38712 35216
rect 122380 35164 122432 35216
rect 163228 35164 163280 35216
rect 490012 35164 490064 35216
rect 145288 33940 145340 33992
rect 259552 33940 259604 33992
rect 148140 33872 148192 33924
rect 287060 33872 287112 33924
rect 158904 33804 158956 33856
rect 429200 33804 429252 33856
rect 169944 33736 169996 33788
rect 572720 33736 572772 33788
rect 3148 33056 3200 33108
rect 7656 33056 7708 33108
rect 173348 33056 173400 33108
rect 580172 33056 580224 33108
rect 31760 32376 31812 32428
rect 120816 32376 120868 32428
rect 142252 32376 142304 32428
rect 219440 32376 219492 32428
rect 154120 31152 154172 31204
rect 332692 31152 332744 31204
rect 150716 31084 150768 31136
rect 329840 31084 329892 31136
rect 167368 31016 167420 31068
rect 542360 31016 542412 31068
rect 145104 29928 145156 29980
rect 251272 29928 251324 29980
rect 145196 29860 145248 29912
rect 253940 29860 253992 29912
rect 150624 29792 150676 29844
rect 324412 29792 324464 29844
rect 156328 29724 156380 29776
rect 391940 29724 391992 29776
rect 160008 29656 160060 29708
rect 434720 29656 434772 29708
rect 167276 29588 167328 29640
rect 535460 29588 535512 29640
rect 141056 28500 141108 28552
rect 201500 28500 201552 28552
rect 143816 28432 143868 28484
rect 242992 28432 243044 28484
rect 152004 28364 152056 28416
rect 346400 28364 346452 28416
rect 154856 28296 154908 28348
rect 378140 28296 378192 28348
rect 171416 28228 171468 28280
rect 397460 28228 397512 28280
rect 139584 27072 139636 27124
rect 186320 27072 186372 27124
rect 171508 27004 171560 27056
rect 411260 27004 411312 27056
rect 156236 26936 156288 26988
rect 398932 26936 398984 26988
rect 165712 26868 165764 26920
rect 524420 26868 524472 26920
rect 140964 25848 141016 25900
rect 201592 25848 201644 25900
rect 149428 25780 149480 25832
rect 303620 25780 303672 25832
rect 156144 25712 156196 25764
rect 401600 25712 401652 25764
rect 157616 25644 157668 25696
rect 414020 25644 414072 25696
rect 167184 25576 167236 25628
rect 540980 25576 541032 25628
rect 167092 25508 167144 25560
rect 545120 25508 545172 25560
rect 135812 24964 135864 25016
rect 140964 24964 141016 25016
rect 140872 24352 140924 24404
rect 198740 24352 198792 24404
rect 148048 24284 148100 24336
rect 292672 24284 292724 24336
rect 98000 24216 98052 24268
rect 132868 24216 132920 24268
rect 149336 24216 149388 24268
rect 313280 24216 313332 24268
rect 27620 24148 27672 24200
rect 127440 24148 127492 24200
rect 157524 24148 157576 24200
rect 416780 24148 416832 24200
rect 3332 24080 3384 24132
rect 179880 24080 179932 24132
rect 182824 24080 182876 24132
rect 579620 24080 579672 24132
rect 135720 23876 135772 23928
rect 139584 23876 139636 23928
rect 3424 23060 3476 23112
rect 174084 23060 174136 23112
rect 172060 22992 172112 23044
rect 404360 22992 404412 23044
rect 42800 22924 42852 22976
rect 128636 22924 128688 22976
rect 157432 22924 157484 22976
rect 409880 22924 409932 22976
rect 11152 22856 11204 22908
rect 125968 22856 126020 22908
rect 160468 22856 160520 22908
rect 455420 22856 455472 22908
rect 9680 22788 9732 22840
rect 126060 22788 126112 22840
rect 136916 22788 136968 22840
rect 148048 22788 148100 22840
rect 164516 22788 164568 22840
rect 499580 22788 499632 22840
rect 118332 22720 118384 22772
rect 580264 22720 580316 22772
rect 138848 22040 138900 22092
rect 143816 22040 143868 22092
rect 160376 21428 160428 21480
rect 454040 21428 454092 21480
rect 170496 21360 170548 21412
rect 514852 21360 514904 21412
rect 144920 20136 144972 20188
rect 262220 20136 262272 20188
rect 145012 20068 145064 20120
rect 255320 20068 255372 20120
rect 255964 20068 256016 20120
rect 456892 20068 456944 20120
rect 124220 20000 124272 20052
rect 134156 20000 134208 20052
rect 143724 20000 143776 20052
rect 241520 20000 241572 20052
rect 242164 20000 242216 20052
rect 449900 20000 449952 20052
rect 67640 19932 67692 19984
rect 130016 19932 130068 19984
rect 157340 19932 157392 19984
rect 415492 19932 415544 19984
rect 143632 18844 143684 18896
rect 234712 18844 234764 18896
rect 164424 18776 164476 18828
rect 509240 18776 509292 18828
rect 168564 18708 168616 18760
rect 553400 18708 553452 18760
rect 168472 18640 168524 18692
rect 556252 18640 556304 18692
rect 168380 18572 168432 18624
rect 560300 18572 560352 18624
rect 160284 17348 160336 17400
rect 445760 17348 445812 17400
rect 160192 17280 160244 17332
rect 448612 17280 448664 17332
rect 164332 17212 164384 17264
rect 506572 17212 506624 17264
rect 144552 16056 144604 16108
rect 237656 16056 237708 16108
rect 151912 15988 151964 16040
rect 342904 15988 342956 16040
rect 153384 15920 153436 15972
rect 361120 15920 361172 15972
rect 163136 15852 163188 15904
rect 492312 15852 492364 15904
rect 147956 14696 148008 14748
rect 289820 14696 289872 14748
rect 149244 14628 149296 14680
rect 311440 14628 311492 14680
rect 154764 14560 154816 14612
rect 386696 14560 386748 14612
rect 160100 14492 160152 14544
rect 453304 14492 453356 14544
rect 163044 14424 163096 14476
rect 488816 14424 488868 14476
rect 151820 13200 151872 13252
rect 349252 13200 349304 13252
rect 155684 13132 155736 13184
rect 361856 13132 361908 13184
rect 162952 13064 163004 13116
rect 484768 13064 484820 13116
rect 106464 11772 106516 11824
rect 132776 11772 132828 11824
rect 136824 11772 136876 11824
rect 145472 11772 145524 11824
rect 156052 11772 156104 11824
rect 400864 11772 400916 11824
rect 63224 11704 63276 11756
rect 129924 11704 129976 11756
rect 138204 11704 138256 11756
rect 167184 11704 167236 11756
rect 169852 11704 169904 11756
rect 574652 11704 574704 11756
rect 234620 11636 234672 11688
rect 235816 11636 235868 11688
rect 259460 11636 259512 11688
rect 260656 11636 260708 11688
rect 150532 10412 150584 10464
rect 322112 10412 322164 10464
rect 117320 10344 117372 10396
rect 134064 10344 134116 10396
rect 154672 10344 154724 10396
rect 379520 10344 379572 10396
rect 25320 10276 25372 10328
rect 93124 10276 93176 10328
rect 99840 10276 99892 10328
rect 132684 10276 132736 10328
rect 168196 10276 168248 10328
rect 539692 10276 539744 10328
rect 147036 9392 147088 9444
rect 270040 9392 270092 9444
rect 146852 9324 146904 9376
rect 277124 9324 277176 9376
rect 146944 9256 146996 9308
rect 276020 9256 276072 9308
rect 149152 9188 149204 9240
rect 315028 9188 315080 9240
rect 315304 9188 315356 9240
rect 465172 9188 465224 9240
rect 153292 9120 153344 9172
rect 358728 9120 358780 9172
rect 85672 9052 85724 9104
rect 131488 9052 131540 9104
rect 161940 9052 161992 9104
rect 463976 9052 464028 9104
rect 78588 8984 78640 9036
rect 128360 8984 128412 9036
rect 162032 8984 162084 9036
rect 467472 8984 467524 9036
rect 64328 8916 64380 8968
rect 126244 8916 126296 8968
rect 165620 8916 165672 8968
rect 521844 8916 521896 8968
rect 142160 7896 142212 7948
rect 222752 7896 222804 7948
rect 53748 7828 53800 7880
rect 129188 7828 129240 7880
rect 149060 7828 149112 7880
rect 307944 7828 307996 7880
rect 45468 7760 45520 7812
rect 128820 7760 128872 7812
rect 150440 7760 150492 7812
rect 323308 7760 323360 7812
rect 35992 7692 36044 7744
rect 127256 7692 127308 7744
rect 154580 7692 154632 7744
rect 385960 7692 386012 7744
rect 34796 7624 34848 7676
rect 127808 7624 127860 7676
rect 172244 7624 172296 7676
rect 440332 7624 440384 7676
rect 24216 7556 24268 7608
rect 122196 7556 122248 7608
rect 164240 7556 164292 7608
rect 504180 7556 504232 7608
rect 102140 7488 102192 7540
rect 103336 7488 103388 7540
rect 146668 6808 146720 6860
rect 268844 6808 268896 6860
rect 146576 6740 146628 6792
rect 272432 6740 272484 6792
rect 146760 6672 146812 6724
rect 273628 6672 273680 6724
rect 147864 6604 147916 6656
rect 296076 6604 296128 6656
rect 105728 6536 105780 6588
rect 133052 6536 133104 6588
rect 155960 6536 156012 6588
rect 394240 6536 394292 6588
rect 84476 6468 84528 6520
rect 131764 6468 131816 6520
rect 161756 6468 161808 6520
rect 462780 6468 462832 6520
rect 80888 6400 80940 6452
rect 131672 6400 131724 6452
rect 161848 6400 161900 6452
rect 466276 6400 466328 6452
rect 77392 6332 77444 6384
rect 131396 6332 131448 6384
rect 161572 6332 161624 6384
rect 469864 6332 469916 6384
rect 52552 6264 52604 6316
rect 128728 6264 128780 6316
rect 161480 6264 161532 6316
rect 471060 6264 471112 6316
rect 19432 6196 19484 6248
rect 125048 6196 125100 6248
rect 161664 6196 161716 6248
rect 473452 6196 473504 6248
rect 18236 6128 18288 6180
rect 125876 6128 125928 6180
rect 169760 6128 169812 6180
rect 572720 6128 572772 6180
rect 132408 6060 132460 6112
rect 190828 6060 190880 6112
rect 136732 5176 136784 5228
rect 154212 5176 154264 5228
rect 101404 5108 101456 5160
rect 113824 5108 113876 5160
rect 114008 5108 114060 5160
rect 134432 5108 134484 5160
rect 138020 5108 138072 5160
rect 169576 5108 169628 5160
rect 66720 5040 66772 5092
rect 103520 5040 103572 5092
rect 103704 5040 103756 5092
rect 130292 5040 130344 5092
rect 140780 5040 140832 5092
rect 206192 5040 206244 5092
rect 15936 4972 15988 5024
rect 101404 4972 101456 5024
rect 147772 4972 147824 5024
rect 294880 4972 294932 5024
rect 436744 4972 436796 5024
rect 28908 4904 28960 4956
rect 127716 4904 127768 4956
rect 154396 4904 154448 4956
rect 364616 4904 364668 4956
rect 6460 4836 6512 4888
rect 10324 4836 10376 4888
rect 13544 4836 13596 4888
rect 125784 4836 125836 4888
rect 136640 4836 136692 4888
rect 157800 4836 157852 4888
rect 159824 4836 159876 4888
rect 436744 4836 436796 4888
rect 479340 4836 479392 4888
rect 8760 4768 8812 4820
rect 126428 4768 126480 4820
rect 138112 4768 138164 4820
rect 162492 4768 162544 4820
rect 162860 4768 162912 4820
rect 493508 4768 493560 4820
rect 572 4088 624 4140
rect 7564 4088 7616 4140
rect 135628 4088 135680 4140
rect 136548 4088 136600 4140
rect 140320 4088 140372 4140
rect 186136 4088 186188 4140
rect 139492 4020 139544 4072
rect 189724 4020 189776 4072
rect 251180 4020 251232 4072
rect 252376 4020 252428 4072
rect 146392 3952 146444 4004
rect 271236 3952 271288 4004
rect 146484 3884 146536 3936
rect 274824 3884 274876 3936
rect 102232 3816 102284 3868
rect 124864 3816 124916 3868
rect 146300 3816 146352 3868
rect 278320 3816 278372 3868
rect 284300 3816 284352 3868
rect 285036 3816 285088 3868
rect 87972 3748 88024 3800
rect 123484 3748 123536 3800
rect 147680 3748 147732 3800
rect 292580 3748 292632 3800
rect 65524 3680 65576 3732
rect 122380 3680 122432 3732
rect 173164 3680 173216 3732
rect 461584 3748 461636 3800
rect 462228 3680 462280 3732
rect 577412 3680 577464 3732
rect 2872 3612 2924 3664
rect 120724 3612 120776 3664
rect 135536 3612 135588 3664
rect 138848 3612 138900 3664
rect 142988 3612 143040 3664
rect 155408 3612 155460 3664
rect 171784 3612 171836 3664
rect 472256 3612 472308 3664
rect 5264 3544 5316 3596
rect 122104 3544 122156 3596
rect 129372 3544 129424 3596
rect 130384 3544 130436 3596
rect 135444 3544 135496 3596
rect 137652 3544 137704 3596
rect 138756 3544 138808 3596
rect 151820 3544 151872 3596
rect 152464 3544 152516 3596
rect 160100 3544 160152 3596
rect 172152 3544 172204 3596
rect 475752 3544 475804 3596
rect 481640 3544 481692 3596
rect 482468 3544 482520 3596
rect 506480 3544 506532 3596
rect 507308 3544 507360 3596
rect 574744 3544 574796 3596
rect 11060 3476 11112 3528
rect 11980 3476 12032 3528
rect 7656 3408 7708 3460
rect 124956 3476 125008 3528
rect 140136 3476 140188 3528
rect 163688 3476 163740 3528
rect 171968 3476 172020 3528
rect 174268 3476 174320 3528
rect 176660 3476 176712 3528
rect 177856 3476 177908 3528
rect 177948 3476 178000 3528
rect 519544 3476 519596 3528
rect 531320 3476 531372 3528
rect 532148 3476 532200 3528
rect 539600 3476 539652 3528
rect 540428 3476 540480 3528
rect 564440 3476 564492 3528
rect 565268 3476 565320 3528
rect 62028 3408 62080 3460
rect 69020 3340 69072 3392
rect 69940 3340 69992 3392
rect 93860 3340 93912 3392
rect 94780 3340 94832 3392
rect 110420 3408 110472 3460
rect 111616 3408 111668 3460
rect 118700 3408 118752 3460
rect 119896 3408 119948 3460
rect 140228 3408 140280 3460
rect 164884 3408 164936 3460
rect 173256 3408 173308 3460
rect 526628 3408 526680 3460
rect 581000 3408 581052 3460
rect 119344 3340 119396 3392
rect 144184 3340 144236 3392
rect 149520 3340 149572 3392
rect 136548 3272 136600 3324
rect 142436 3272 142488 3324
rect 142804 3272 142856 3324
rect 150624 3272 150676 3324
rect 118792 3204 118844 3256
rect 123576 3204 123628 3256
rect 140044 3204 140096 3256
rect 144736 3204 144788 3256
rect 144460 3136 144512 3188
rect 153016 3340 153068 3392
rect 166264 3340 166316 3392
rect 170772 3340 170824 3392
rect 175924 3340 175976 3392
rect 212172 3340 212224 3392
rect 307760 3340 307812 3392
rect 309048 3340 309100 3392
rect 316040 3340 316092 3392
rect 317328 3340 317380 3392
rect 324412 3340 324464 3392
rect 325608 3340 325660 3392
rect 332600 3340 332652 3392
rect 333888 3340 333940 3392
rect 340972 3340 341024 3392
rect 342168 3340 342220 3392
rect 349252 3340 349304 3392
rect 350448 3340 350500 3392
rect 365720 3340 365772 3392
rect 367008 3340 367060 3392
rect 374092 3340 374144 3392
rect 375288 3340 375340 3392
rect 382372 3340 382424 3392
rect 383568 3340 383620 3392
rect 390652 3340 390704 3392
rect 391848 3340 391900 3392
rect 398932 3340 398984 3392
rect 400128 3340 400180 3392
rect 407120 3340 407172 3392
rect 408408 3340 408460 3392
rect 415400 3340 415452 3392
rect 416688 3340 416740 3392
rect 423772 3340 423824 3392
rect 424968 3340 425020 3392
rect 432052 3340 432104 3392
rect 433248 3340 433300 3392
rect 440240 3340 440292 3392
rect 441528 3340 441580 3392
rect 448612 3340 448664 3392
rect 449808 3340 449860 3392
rect 456892 3340 456944 3392
rect 458088 3340 458140 3392
rect 174544 3272 174596 3324
rect 195612 3272 195664 3324
rect 171876 3204 171928 3256
rect 177948 3204 178000 3256
rect 165068 3068 165120 3120
rect 171968 3068 172020 3120
<< metal2 >>
rect 8086 703520 8198 704960
rect 23492 703582 24164 703610
rect 8128 700330 8156 703520
rect 8116 700324 8168 700330
rect 8116 700266 8168 700272
rect 2778 684312 2834 684321
rect 2778 684247 2834 684256
rect 2792 683738 2820 684247
rect 2780 683732 2832 683738
rect 2780 683674 2832 683680
rect 4804 683732 4856 683738
rect 4804 683674 4856 683680
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3332 632120 3384 632126
rect 3330 632088 3332 632097
rect 3384 632088 3386 632097
rect 3330 632023 3386 632032
rect 3146 580000 3202 580009
rect 3146 579935 3202 579944
rect 3160 579698 3188 579935
rect 3148 579692 3200 579698
rect 3148 579634 3200 579640
rect 3146 553888 3202 553897
rect 3146 553823 3202 553832
rect 3160 553450 3188 553823
rect 3148 553444 3200 553450
rect 3148 553386 3200 553392
rect 3330 527912 3386 527921
rect 3330 527847 3332 527856
rect 3384 527847 3386 527856
rect 3332 527818 3384 527824
rect 3330 514856 3386 514865
rect 3330 514791 3332 514800
rect 3384 514791 3386 514800
rect 3332 514762 3384 514768
rect 2778 501800 2834 501809
rect 2778 501735 2834 501744
rect 2792 501090 2820 501735
rect 2780 501084 2832 501090
rect 2780 501026 2832 501032
rect 3054 462632 3110 462641
rect 3054 462567 3110 462576
rect 3068 462398 3096 462567
rect 3056 462392 3108 462398
rect 3056 462334 3108 462340
rect 2962 449576 3018 449585
rect 2962 449511 3018 449520
rect 2976 448594 3004 449511
rect 2964 448588 3016 448594
rect 2964 448530 3016 448536
rect 3330 423600 3386 423609
rect 3330 423535 3386 423544
rect 3344 422346 3372 423535
rect 3332 422340 3384 422346
rect 3332 422282 3384 422288
rect 3332 397520 3384 397526
rect 3330 397488 3332 397497
rect 3384 397488 3386 397497
rect 3330 397423 3386 397432
rect 3330 371376 3386 371385
rect 3330 371311 3386 371320
rect 3344 371278 3372 371311
rect 3332 371272 3384 371278
rect 3332 371214 3384 371220
rect 3330 358456 3386 358465
rect 3330 358391 3386 358400
rect 3344 357474 3372 358391
rect 3332 357468 3384 357474
rect 3332 357410 3384 357416
rect 3330 345400 3386 345409
rect 3330 345335 3386 345344
rect 3344 345098 3372 345335
rect 3332 345092 3384 345098
rect 3332 345034 3384 345040
rect 3146 319288 3202 319297
rect 3146 319223 3202 319232
rect 3160 318850 3188 319223
rect 3148 318844 3200 318850
rect 3148 318786 3200 318792
rect 3330 306232 3386 306241
rect 3330 306167 3386 306176
rect 3344 305046 3372 306167
rect 3332 305040 3384 305046
rect 3332 304982 3384 304988
rect 3330 293176 3386 293185
rect 3330 293111 3386 293120
rect 3344 292602 3372 293111
rect 3332 292596 3384 292602
rect 3332 292538 3384 292544
rect 3238 267200 3294 267209
rect 3238 267135 3294 267144
rect 3252 266422 3280 267135
rect 3240 266416 3292 266422
rect 3240 266358 3292 266364
rect 2962 254144 3018 254153
rect 2962 254079 3018 254088
rect 2976 253978 3004 254079
rect 2964 253972 3016 253978
rect 2964 253914 3016 253920
rect 2870 228032 2926 228041
rect 2870 227967 2926 227976
rect 2884 227798 2912 227967
rect 2872 227792 2924 227798
rect 2872 227734 2924 227740
rect 3330 214976 3386 214985
rect 3330 214911 3386 214920
rect 3344 213994 3372 214911
rect 3332 213988 3384 213994
rect 3332 213930 3384 213936
rect 3330 201920 3386 201929
rect 3330 201855 3386 201864
rect 3344 201550 3372 201855
rect 3332 201544 3384 201550
rect 3332 201486 3384 201492
rect 3330 188864 3386 188873
rect 3330 188799 3386 188808
rect 3344 187746 3372 188799
rect 3332 187740 3384 187746
rect 3332 187682 3384 187688
rect 3332 176656 3384 176662
rect 3332 176598 3384 176604
rect 3344 175953 3372 176598
rect 3330 175944 3386 175953
rect 3330 175879 3386 175888
rect 3332 162920 3384 162926
rect 3330 162888 3332 162897
rect 3384 162888 3386 162897
rect 3330 162823 3386 162832
rect 2870 136776 2926 136785
rect 2870 136711 2926 136720
rect 2884 136678 2912 136711
rect 2872 136672 2924 136678
rect 2872 136614 2924 136620
rect 3332 111784 3384 111790
rect 3332 111726 3384 111732
rect 3344 110673 3372 111726
rect 3330 110664 3386 110673
rect 3330 110599 3386 110608
rect 3436 78985 3464 658135
rect 3528 150074 3556 671191
rect 3698 619168 3754 619177
rect 3698 619103 3754 619112
rect 3606 606112 3662 606121
rect 3606 606047 3662 606056
rect 3516 150068 3568 150074
rect 3516 150010 3568 150016
rect 3514 149832 3570 149841
rect 3514 149767 3570 149776
rect 3528 149122 3556 149767
rect 3516 149116 3568 149122
rect 3516 149058 3568 149064
rect 3516 139460 3568 139466
rect 3516 139402 3568 139408
rect 3528 97617 3556 139402
rect 3514 97608 3570 97617
rect 3514 97543 3570 97552
rect 3514 84688 3570 84697
rect 3514 84623 3570 84632
rect 3422 78976 3478 78985
rect 3422 78911 3478 78920
rect 3528 77518 3556 84623
rect 3620 79121 3648 606047
rect 3712 151094 3740 619103
rect 3790 566944 3846 566953
rect 3790 566879 3846 566888
rect 3804 173194 3832 566879
rect 3882 475688 3938 475697
rect 3882 475623 3938 475632
rect 3896 461650 3924 475623
rect 3884 461644 3936 461650
rect 3884 461586 3936 461592
rect 3882 410544 3938 410553
rect 3882 410479 3938 410488
rect 3792 173188 3844 173194
rect 3792 173130 3844 173136
rect 3700 151088 3752 151094
rect 3700 151030 3752 151036
rect 3700 150068 3752 150074
rect 3700 150010 3752 150016
rect 3712 148374 3740 150010
rect 3700 148368 3752 148374
rect 3700 148310 3752 148316
rect 3896 140214 3924 410479
rect 3974 241088 4030 241097
rect 3974 241023 4030 241032
rect 3884 140208 3936 140214
rect 3884 140150 3936 140156
rect 3988 79354 4016 241023
rect 4816 118658 4844 683674
rect 7564 632120 7616 632126
rect 7564 632062 7616 632068
rect 4896 501084 4948 501090
rect 4896 501026 4948 501032
rect 4804 118652 4856 118658
rect 4804 118594 4856 118600
rect 3976 79348 4028 79354
rect 3976 79290 4028 79296
rect 4908 79257 4936 501026
rect 7576 120086 7604 632062
rect 17224 579692 17276 579698
rect 17224 579634 17276 579640
rect 8944 527876 8996 527882
rect 8944 527818 8996 527824
rect 7656 136740 7708 136746
rect 7656 136682 7708 136688
rect 7564 120080 7616 120086
rect 7564 120022 7616 120028
rect 4894 79248 4950 79257
rect 4894 79183 4950 79192
rect 3606 79112 3662 79121
rect 3606 79047 3662 79056
rect 3516 77512 3568 77518
rect 3516 77454 3568 77460
rect 1398 72448 1454 72457
rect 1398 72383 1454 72392
rect 572 4140 624 4146
rect 572 4082 624 4088
rect 584 480 612 4082
rect 542 -960 654 480
rect 1412 354 1440 72383
rect 3424 71664 3476 71670
rect 3422 71632 3424 71641
rect 3476 71632 3478 71641
rect 3422 71567 3478 71576
rect 3056 59356 3108 59362
rect 3056 59298 3108 59304
rect 3068 58585 3096 59298
rect 3054 58576 3110 58585
rect 3054 58511 3110 58520
rect 3424 45552 3476 45558
rect 3422 45520 3424 45529
rect 3476 45520 3478 45529
rect 3422 45455 3478 45464
rect 7564 36576 7616 36582
rect 7564 36518 7616 36524
rect 3148 33108 3200 33114
rect 3148 33050 3200 33056
rect 3160 32473 3188 33050
rect 3146 32464 3202 32473
rect 3146 32399 3202 32408
rect 3332 24132 3384 24138
rect 3332 24074 3384 24080
rect 3344 19417 3372 24074
rect 3424 23112 3476 23118
rect 3424 23054 3476 23060
rect 3330 19408 3386 19417
rect 3330 19343 3386 19352
rect 3436 6497 3464 23054
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 6460 4888 6512 4894
rect 4066 4856 4122 4865
rect 6460 4830 6512 4836
rect 4066 4791 4122 4800
rect 2872 3664 2924 3670
rect 2872 3606 2924 3612
rect 2884 480 2912 3606
rect 4080 480 4108 4791
rect 5264 3596 5316 3602
rect 5264 3538 5316 3544
rect 5276 480 5304 3538
rect 6472 480 6500 4830
rect 7576 4146 7604 36518
rect 7668 33114 7696 136682
rect 8956 122806 8984 527818
rect 10324 422340 10376 422346
rect 10324 422282 10376 422288
rect 9036 135312 9088 135318
rect 9036 135254 9088 135260
rect 8944 122800 8996 122806
rect 8944 122742 8996 122748
rect 9048 71670 9076 135254
rect 10336 126954 10364 422282
rect 13084 318844 13136 318850
rect 13084 318786 13136 318792
rect 13096 129742 13124 318786
rect 14464 162920 14516 162926
rect 14464 162862 14516 162868
rect 14476 133890 14504 162862
rect 14464 133884 14516 133890
rect 14464 133826 14516 133832
rect 13084 129736 13136 129742
rect 13084 129678 13136 129684
rect 10324 126948 10376 126954
rect 10324 126890 10376 126896
rect 17236 121446 17264 579634
rect 18604 266416 18656 266422
rect 18604 266358 18656 266364
rect 17868 180124 17920 180130
rect 17868 180066 17920 180072
rect 17880 176662 17908 180066
rect 17868 176656 17920 176662
rect 17868 176598 17920 176604
rect 18616 131102 18644 266358
rect 23492 146946 23520 703582
rect 24136 703474 24164 703582
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 24320 703474 24348 703520
rect 24136 703446 24348 703474
rect 31024 213988 31076 213994
rect 31024 213930 31076 213936
rect 23480 146940 23532 146946
rect 23480 146882 23532 146888
rect 21364 133952 21416 133958
rect 21364 133894 21416 133900
rect 18604 131096 18656 131102
rect 18604 131038 18656 131044
rect 17224 121440 17276 121446
rect 17224 121382 17276 121388
rect 21376 111790 21404 133894
rect 31036 132462 31064 213930
rect 31024 132456 31076 132462
rect 31024 132398 31076 132404
rect 40052 117298 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 234632 703582 235028 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 703050 73016 703520
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 53104 461644 53156 461650
rect 53104 461586 53156 461592
rect 44824 448588 44876 448594
rect 44824 448530 44876 448536
rect 40040 117292 40092 117298
rect 40040 117234 40092 117240
rect 21364 111784 21416 111790
rect 21364 111726 21416 111732
rect 44836 78810 44864 448530
rect 53116 124166 53144 461586
rect 62132 230574 62514 230602
rect 62132 195974 62160 230574
rect 62120 195968 62172 195974
rect 62120 195910 62172 195916
rect 53104 124160 53156 124166
rect 53104 124102 53156 124108
rect 71792 79422 71820 702986
rect 89180 700398 89208 703520
rect 89168 700392 89220 700398
rect 89168 700334 89220 700340
rect 105464 699718 105492 703520
rect 137848 700330 137876 703520
rect 154132 702434 154160 703520
rect 170324 702434 170352 703520
rect 202800 703050 202828 703520
rect 201500 703044 201552 703050
rect 201500 702986 201552 702992
rect 202788 703044 202840 703050
rect 202788 702986 202840 702992
rect 153856 702406 154160 702434
rect 169772 702406 170352 702434
rect 119344 700324 119396 700330
rect 119344 700266 119396 700272
rect 137836 700324 137888 700330
rect 137836 700266 137888 700272
rect 105452 699712 105504 699718
rect 105452 699654 105504 699660
rect 106924 699712 106976 699718
rect 106924 699654 106976 699660
rect 86224 397520 86276 397526
rect 86224 397462 86276 397468
rect 84844 371272 84896 371278
rect 84844 371214 84896 371220
rect 84856 128314 84884 371214
rect 84844 128308 84896 128314
rect 84844 128250 84896 128256
rect 86236 79626 86264 397462
rect 92492 195906 92520 230588
rect 92480 195900 92532 195906
rect 92480 195842 92532 195848
rect 106936 115938 106964 699654
rect 115204 553444 115256 553450
rect 115204 553386 115256 553392
rect 106924 115932 106976 115938
rect 106924 115874 106976 115880
rect 86224 79620 86276 79626
rect 86224 79562 86276 79568
rect 71780 79416 71832 79422
rect 115216 79393 115244 553386
rect 118700 429888 118752 429894
rect 118700 429830 118752 429836
rect 118608 404388 118660 404394
rect 118608 404330 118660 404336
rect 118516 351960 118568 351966
rect 118516 351902 118568 351908
rect 116584 345092 116636 345098
rect 116584 345034 116636 345040
rect 115296 136672 115348 136678
rect 115296 136614 115348 136620
rect 115308 79490 115336 136614
rect 116596 79762 116624 345034
rect 118240 142180 118292 142186
rect 118240 142122 118292 142128
rect 118148 141568 118200 141574
rect 118148 141510 118200 141516
rect 118056 141500 118108 141506
rect 118056 141442 118108 141448
rect 117318 137592 117374 137601
rect 117318 137527 117374 137536
rect 117332 136746 117360 137527
rect 117320 136740 117372 136746
rect 117320 136682 117372 136688
rect 117318 136096 117374 136105
rect 117318 136031 117374 136040
rect 117332 135318 117360 136031
rect 117320 135312 117372 135318
rect 117320 135254 117372 135260
rect 117318 134600 117374 134609
rect 117318 134535 117374 134544
rect 117332 133958 117360 134535
rect 117320 133952 117372 133958
rect 117320 133894 117372 133900
rect 117412 133884 117464 133890
rect 117412 133826 117464 133832
rect 117424 133113 117452 133826
rect 117410 133104 117466 133113
rect 117410 133039 117466 133048
rect 117320 132456 117372 132462
rect 117320 132398 117372 132404
rect 117332 131617 117360 132398
rect 117318 131608 117374 131617
rect 117318 131543 117374 131552
rect 117320 131096 117372 131102
rect 117320 131038 117372 131044
rect 117332 130121 117360 131038
rect 117318 130112 117374 130121
rect 117318 130047 117374 130056
rect 117320 129736 117372 129742
rect 117320 129678 117372 129684
rect 117332 128625 117360 129678
rect 117318 128616 117374 128625
rect 117318 128551 117374 128560
rect 117320 128308 117372 128314
rect 117320 128250 117372 128256
rect 117332 127129 117360 128250
rect 117318 127120 117374 127129
rect 117318 127055 117374 127064
rect 117320 126948 117372 126954
rect 117320 126890 117372 126896
rect 117332 125633 117360 126890
rect 117318 125624 117374 125633
rect 117318 125559 117374 125568
rect 117320 124160 117372 124166
rect 117318 124128 117320 124137
rect 117372 124128 117374 124137
rect 117318 124063 117374 124072
rect 117320 122800 117372 122806
rect 117320 122742 117372 122748
rect 117332 122641 117360 122742
rect 117318 122632 117374 122641
rect 117318 122567 117374 122576
rect 117320 121440 117372 121446
rect 117320 121382 117372 121388
rect 117332 121145 117360 121382
rect 117318 121136 117374 121145
rect 117318 121071 117374 121080
rect 117320 120080 117372 120086
rect 117320 120022 117372 120028
rect 117332 119649 117360 120022
rect 117318 119640 117374 119649
rect 117318 119575 117374 119584
rect 117320 118652 117372 118658
rect 117320 118594 117372 118600
rect 117332 118153 117360 118594
rect 117318 118144 117374 118153
rect 117318 118079 117374 118088
rect 117320 117292 117372 117298
rect 117320 117234 117372 117240
rect 117332 116657 117360 117234
rect 117318 116648 117374 116657
rect 117318 116583 117374 116592
rect 117320 115932 117372 115938
rect 117320 115874 117372 115880
rect 117332 115161 117360 115874
rect 117318 115152 117374 115161
rect 117318 115087 117374 115096
rect 118068 113665 118096 141442
rect 118054 113656 118110 113665
rect 118054 113591 118110 113600
rect 118160 91225 118188 141510
rect 118252 92721 118280 142122
rect 118332 140276 118384 140282
rect 118332 140218 118384 140224
rect 118238 92712 118294 92721
rect 118238 92647 118294 92656
rect 118146 91216 118202 91225
rect 118146 91151 118202 91160
rect 118344 89729 118372 140218
rect 118424 139528 118476 139534
rect 118424 139470 118476 139476
rect 118330 89720 118386 89729
rect 118330 89655 118386 89664
rect 118436 88233 118464 139470
rect 118528 94217 118556 351902
rect 118620 95713 118648 404330
rect 118712 103193 118740 429830
rect 119068 147008 119120 147014
rect 119068 146950 119120 146956
rect 118884 144220 118936 144226
rect 118884 144162 118936 144168
rect 118792 140072 118844 140078
rect 118792 140014 118844 140020
rect 118804 104689 118832 140014
rect 118896 107681 118924 144162
rect 118976 141432 119028 141438
rect 118976 141374 119028 141380
rect 118882 107672 118938 107681
rect 118882 107607 118938 107616
rect 118988 106185 119016 141374
rect 119080 112169 119108 146950
rect 119160 145580 119212 145586
rect 119160 145522 119212 145528
rect 119066 112160 119122 112169
rect 119066 112095 119122 112104
rect 119172 110673 119200 145522
rect 119252 140140 119304 140146
rect 119252 140082 119304 140088
rect 119158 110664 119214 110673
rect 119158 110599 119214 110608
rect 119264 109177 119292 140082
rect 119250 109168 119306 109177
rect 119250 109103 119306 109112
rect 118974 106176 119030 106185
rect 118974 106111 119030 106120
rect 118790 104680 118846 104689
rect 118790 104615 118846 104624
rect 118698 103184 118754 103193
rect 118698 103119 118754 103128
rect 118606 95704 118662 95713
rect 118606 95639 118662 95648
rect 118514 94208 118570 94217
rect 118514 94143 118570 94152
rect 118422 88224 118478 88233
rect 118422 88159 118478 88168
rect 118422 86728 118478 86737
rect 118422 86663 118478 86672
rect 118330 82240 118386 82249
rect 118330 82175 118386 82184
rect 116584 79756 116636 79762
rect 116584 79698 116636 79704
rect 115296 79484 115348 79490
rect 115296 79426 115348 79432
rect 71780 79358 71832 79364
rect 115202 79384 115258 79393
rect 115202 79319 115258 79328
rect 44824 78804 44876 78810
rect 44824 78746 44876 78752
rect 93124 78600 93176 78606
rect 93124 78542 93176 78548
rect 89720 78056 89772 78062
rect 89720 77998 89772 78004
rect 53840 77988 53892 77994
rect 53840 77930 53892 77936
rect 10322 77888 10378 77897
rect 10322 77823 10378 77832
rect 9036 71664 9088 71670
rect 9036 71606 9088 71612
rect 7656 33108 7708 33114
rect 7656 33050 7708 33056
rect 9680 22840 9732 22846
rect 9680 22782 9732 22788
rect 8760 4820 8812 4826
rect 8760 4762 8812 4768
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 7656 3460 7708 3466
rect 7656 3402 7708 3408
rect 7668 480 7696 3402
rect 8772 480 8800 4762
rect 1646 354 1758 480
rect 1412 326 1758 354
rect 1646 -960 1758 326
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9692 354 9720 22782
rect 10336 4894 10364 77823
rect 37278 76664 37334 76673
rect 37278 76599 37334 76608
rect 20718 76528 20774 76537
rect 20718 76463 20774 76472
rect 16580 71120 16632 71126
rect 16580 71062 16632 71068
rect 11060 71052 11112 71058
rect 11060 70994 11112 71000
rect 10324 4888 10376 4894
rect 10324 4830 10376 4836
rect 11072 3534 11100 70994
rect 13820 51740 13872 51746
rect 13820 51682 13872 51688
rect 11152 22908 11204 22914
rect 11152 22850 11204 22856
rect 11060 3528 11112 3534
rect 11060 3470 11112 3476
rect 11164 480 11192 22850
rect 13832 16574 13860 51682
rect 16592 16574 16620 71062
rect 19338 25528 19394 25537
rect 19338 25463 19394 25472
rect 19352 16574 19380 25463
rect 20732 16574 20760 76463
rect 30380 73840 30432 73846
rect 30380 73782 30432 73788
rect 35898 73808 35954 73817
rect 26240 72480 26292 72486
rect 26240 72422 26292 72428
rect 22098 68232 22154 68241
rect 22098 68167 22154 68176
rect 22112 16574 22140 68167
rect 13832 16546 14320 16574
rect 16592 16546 17080 16574
rect 19352 16546 20208 16574
rect 20732 16546 21864 16574
rect 22112 16546 22600 16574
rect 13544 4888 13596 4894
rect 13544 4830 13596 4836
rect 11980 3528 12032 3534
rect 11980 3470 12032 3476
rect 9926 354 10038 480
rect 9692 326 10038 354
rect 9926 -960 10038 326
rect 11122 -960 11234 480
rect 11992 354 12020 3470
rect 13556 480 13584 4830
rect 12318 354 12430 480
rect 11992 326 12430 354
rect 12318 -960 12430 326
rect 13514 -960 13626 480
rect 14292 354 14320 16546
rect 15936 5024 15988 5030
rect 15936 4966 15988 4972
rect 15948 480 15976 4966
rect 17052 480 17080 16546
rect 19432 6248 19484 6254
rect 19432 6190 19484 6196
rect 18236 6180 18288 6186
rect 18236 6122 18288 6128
rect 18248 480 18276 6122
rect 19444 480 19472 6190
rect 14710 354 14822 480
rect 14292 326 14822 354
rect 14710 -960 14822 326
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20180 354 20208 16546
rect 21836 480 21864 16546
rect 20598 354 20710 480
rect 20180 326 20710 354
rect 20598 -960 20710 326
rect 21794 -960 21906 480
rect 22572 354 22600 16546
rect 25320 10328 25372 10334
rect 25320 10270 25372 10276
rect 24216 7608 24268 7614
rect 24216 7550 24268 7556
rect 24228 480 24256 7550
rect 25332 480 25360 10270
rect 22990 354 23102 480
rect 22572 326 23102 354
rect 22990 -960 23102 326
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 72422
rect 29000 71188 29052 71194
rect 29000 71130 29052 71136
rect 27620 24200 27672 24206
rect 27620 24142 27672 24148
rect 27632 16574 27660 24142
rect 29012 16574 29040 71130
rect 30392 16574 30420 73782
rect 35898 73743 35954 73752
rect 33140 66904 33192 66910
rect 33140 66846 33192 66852
rect 31760 32428 31812 32434
rect 31760 32370 31812 32376
rect 31772 16574 31800 32370
rect 33152 16574 33180 66846
rect 35912 16574 35940 73743
rect 37292 16574 37320 76599
rect 51080 75336 51132 75342
rect 51080 75278 51132 75284
rect 49700 75268 49752 75274
rect 49700 75210 49752 75216
rect 46940 75200 46992 75206
rect 46940 75142 46992 75148
rect 40038 72584 40094 72593
rect 40038 72519 40094 72528
rect 38660 35216 38712 35222
rect 38660 35158 38712 35164
rect 38672 16574 38700 35158
rect 40052 16574 40080 72519
rect 44180 69692 44232 69698
rect 44180 69634 44232 69640
rect 42800 22976 42852 22982
rect 42800 22918 42852 22924
rect 27632 16546 27752 16574
rect 29012 16546 30144 16574
rect 30392 16546 30880 16574
rect 31772 16546 31984 16574
rect 33152 16546 33640 16574
rect 35912 16546 36768 16574
rect 37292 16546 38424 16574
rect 38672 16546 39160 16574
rect 40052 16546 40264 16574
rect 27724 480 27752 16546
rect 28908 4956 28960 4962
rect 28908 4898 28960 4904
rect 28920 480 28948 4898
rect 30116 480 30144 16546
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 30852 354 30880 16546
rect 31270 354 31382 480
rect 30852 326 31382 354
rect 31956 354 31984 16546
rect 33612 480 33640 16546
rect 35992 7744 36044 7750
rect 35992 7686 36044 7692
rect 34796 7676 34848 7682
rect 34796 7618 34848 7624
rect 34808 480 34836 7618
rect 36004 480 36032 7686
rect 32374 354 32486 480
rect 31956 326 32486 354
rect 31270 -960 31382 326
rect 32374 -960 32486 326
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 36740 354 36768 16546
rect 38396 480 38424 16546
rect 37158 354 37270 480
rect 36740 326 37270 354
rect 37158 -960 37270 326
rect 38354 -960 38466 480
rect 39132 354 39160 16546
rect 39550 354 39662 480
rect 39132 326 39662 354
rect 40236 354 40264 16546
rect 41878 7576 41934 7585
rect 41878 7511 41934 7520
rect 41892 480 41920 7511
rect 40654 354 40766 480
rect 40236 326 40766 354
rect 39550 -960 39662 326
rect 40654 -960 40766 326
rect 41850 -960 41962 480
rect 42812 354 42840 22918
rect 44192 16574 44220 69634
rect 45560 37936 45612 37942
rect 45560 37878 45612 37884
rect 45572 16574 45600 37878
rect 46952 16574 46980 75142
rect 48320 71256 48372 71262
rect 48320 71198 48372 71204
rect 48332 16574 48360 71198
rect 49712 16574 49740 75210
rect 44192 16546 44312 16574
rect 45572 16546 46704 16574
rect 46952 16546 47440 16574
rect 48332 16546 48544 16574
rect 49712 16546 50200 16574
rect 44284 480 44312 16546
rect 45468 7812 45520 7818
rect 45468 7754 45520 7760
rect 45480 480 45508 7754
rect 46676 480 46704 16546
rect 43046 354 43158 480
rect 42812 326 43158 354
rect 43046 -960 43158 326
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47412 354 47440 16546
rect 47830 354 47942 480
rect 47412 326 47942 354
rect 48516 354 48544 16546
rect 50172 480 50200 16546
rect 48934 354 49046 480
rect 48516 326 49046 354
rect 47830 -960 47942 326
rect 48934 -960 49046 326
rect 50130 -960 50242 480
rect 51092 354 51120 75278
rect 53852 16574 53880 77930
rect 70400 76628 70452 76634
rect 70400 76570 70452 76576
rect 69020 76560 69072 76566
rect 69020 76502 69072 76508
rect 60740 69760 60792 69766
rect 60740 69702 60792 69708
rect 55218 69592 55274 69601
rect 55218 69527 55274 69536
rect 55232 16574 55260 69527
rect 57978 68368 58034 68377
rect 57978 68303 58034 68312
rect 57992 16574 58020 68303
rect 60752 16574 60780 69702
rect 67640 19984 67692 19990
rect 67640 19926 67692 19932
rect 53852 16546 54984 16574
rect 55232 16546 56088 16574
rect 57992 16546 58480 16574
rect 60752 16546 60872 16574
rect 53748 7880 53800 7886
rect 53748 7822 53800 7828
rect 52552 6316 52604 6322
rect 52552 6258 52604 6264
rect 52564 480 52592 6258
rect 53760 480 53788 7822
rect 54956 480 54984 16546
rect 56060 480 56088 16546
rect 57242 8936 57298 8945
rect 57242 8871 57298 8880
rect 57256 480 57284 8871
rect 58452 480 58480 16546
rect 59634 9072 59690 9081
rect 59634 9007 59690 9016
rect 59648 480 59676 9007
rect 60844 480 60872 16546
rect 63224 11756 63276 11762
rect 63224 11698 63276 11704
rect 62028 3460 62080 3466
rect 62028 3402 62080 3408
rect 62040 480 62068 3402
rect 63236 480 63264 11698
rect 64328 8968 64380 8974
rect 64328 8910 64380 8916
rect 64340 480 64368 8910
rect 66720 5092 66772 5098
rect 66720 5034 66772 5040
rect 65524 3732 65576 3738
rect 65524 3674 65576 3680
rect 65536 480 65564 3674
rect 66732 480 66760 5034
rect 51326 354 51438 480
rect 51092 326 51438 354
rect 51326 -960 51438 326
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67652 354 67680 19926
rect 69032 3398 69060 76502
rect 69112 73908 69164 73914
rect 69112 73850 69164 73856
rect 69020 3392 69072 3398
rect 69020 3334 69072 3340
rect 69124 480 69152 73850
rect 70412 16574 70440 76570
rect 75918 75168 75974 75177
rect 75918 75103 75974 75112
rect 71778 73944 71834 73953
rect 71778 73879 71834 73888
rect 71792 16574 71820 73879
rect 73158 65512 73214 65521
rect 73158 65447 73214 65456
rect 73172 16574 73200 65447
rect 74538 44840 74594 44849
rect 74538 44775 74594 44784
rect 74552 16574 74580 44775
rect 70412 16546 71544 16574
rect 71792 16546 72648 16574
rect 73172 16546 73384 16574
rect 74552 16546 75040 16574
rect 69940 3392 69992 3398
rect 69940 3334 69992 3340
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 69952 354 69980 3334
rect 71516 480 71544 16546
rect 72620 480 72648 16546
rect 70278 354 70390 480
rect 69952 326 70390 354
rect 70278 -960 70390 326
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73356 354 73384 16546
rect 75012 480 75040 16546
rect 73774 354 73886 480
rect 73356 326 73886 354
rect 73774 -960 73886 326
rect 74970 -960 75082 480
rect 75932 354 75960 75103
rect 85580 72548 85632 72554
rect 85580 72490 85632 72496
rect 82820 71324 82872 71330
rect 82820 71266 82872 71272
rect 78680 69828 78732 69834
rect 78680 69770 78732 69776
rect 78692 16574 78720 69770
rect 81440 44872 81492 44878
rect 81440 44814 81492 44820
rect 81452 16574 81480 44814
rect 82832 16574 82860 71266
rect 85592 16574 85620 72490
rect 88340 55888 88392 55894
rect 88340 55830 88392 55836
rect 88352 16574 88380 55830
rect 89732 16574 89760 77998
rect 91098 69728 91154 69737
rect 91098 69663 91154 69672
rect 91112 16574 91140 69663
rect 78692 16546 79272 16574
rect 81452 16546 81664 16574
rect 82832 16546 83320 16574
rect 85592 16546 86448 16574
rect 88352 16546 89208 16574
rect 89732 16546 89944 16574
rect 91112 16546 91600 16574
rect 78588 9036 78640 9042
rect 78588 8978 78640 8984
rect 77392 6384 77444 6390
rect 77392 6326 77444 6332
rect 77404 480 77432 6326
rect 78600 480 78628 8978
rect 76166 354 76278 480
rect 75932 326 76278 354
rect 76166 -960 76278 326
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79244 354 79272 16546
rect 80888 6452 80940 6458
rect 80888 6394 80940 6400
rect 80900 480 80928 6394
rect 79662 354 79774 480
rect 79244 326 79774 354
rect 79662 -960 79774 326
rect 80858 -960 80970 480
rect 81636 354 81664 16546
rect 83292 480 83320 16546
rect 85672 9104 85724 9110
rect 85672 9046 85724 9052
rect 84476 6520 84528 6526
rect 84476 6462 84528 6468
rect 84488 480 84516 6462
rect 85684 480 85712 9046
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86420 354 86448 16546
rect 87972 3800 88024 3806
rect 87972 3742 88024 3748
rect 87984 480 88012 3742
rect 89180 480 89208 16546
rect 86838 354 86950 480
rect 86420 326 86950 354
rect 86838 -960 86950 326
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 89916 354 89944 16546
rect 91572 480 91600 16546
rect 93136 10334 93164 78542
rect 113824 78260 113876 78266
rect 113824 78202 113876 78208
rect 110420 78192 110472 78198
rect 110420 78134 110472 78140
rect 93860 76696 93912 76702
rect 93860 76638 93912 76644
rect 93124 10328 93176 10334
rect 93124 10270 93176 10276
rect 92754 9208 92810 9217
rect 92754 9143 92810 9152
rect 92768 480 92796 9143
rect 93872 3398 93900 76638
rect 107660 75404 107712 75410
rect 107660 75346 107712 75352
rect 93952 73976 94004 73982
rect 93952 73918 94004 73924
rect 93860 3392 93912 3398
rect 93860 3334 93912 3340
rect 93964 480 93992 73918
rect 96620 72616 96672 72622
rect 96620 72558 96672 72564
rect 95240 57248 95292 57254
rect 95240 57190 95292 57196
rect 95252 16574 95280 57190
rect 96632 16574 96660 72558
rect 100760 71392 100812 71398
rect 100760 71334 100812 71340
rect 98000 24268 98052 24274
rect 98000 24210 98052 24216
rect 98012 16574 98040 24210
rect 95252 16546 95832 16574
rect 96632 16546 97488 16574
rect 98012 16546 98224 16574
rect 94780 3392 94832 3398
rect 94780 3334 94832 3340
rect 90334 354 90446 480
rect 89916 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 94792 354 94820 3334
rect 95118 354 95230 480
rect 94792 326 95230 354
rect 95804 354 95832 16546
rect 97460 480 97488 16546
rect 96222 354 96334 480
rect 95804 326 96334 354
rect 95118 -960 95230 326
rect 96222 -960 96334 326
rect 97418 -960 97530 480
rect 98196 354 98224 16546
rect 99840 10328 99892 10334
rect 99840 10270 99892 10276
rect 99852 480 99880 10270
rect 98614 354 98726 480
rect 98196 326 98726 354
rect 98614 -960 98726 326
rect 99810 -960 99922 480
rect 100772 354 100800 71334
rect 103520 69896 103572 69902
rect 103520 69838 103572 69844
rect 102140 61396 102192 61402
rect 102140 61338 102192 61344
rect 102152 7546 102180 61338
rect 103532 16574 103560 69838
rect 107672 16574 107700 75346
rect 103532 16546 104112 16574
rect 107672 16546 108160 16574
rect 102140 7540 102192 7546
rect 102140 7482 102192 7488
rect 103336 7540 103388 7546
rect 103336 7482 103388 7488
rect 101404 5160 101456 5166
rect 101404 5102 101456 5108
rect 101416 5030 101444 5102
rect 101404 5024 101456 5030
rect 101404 4966 101456 4972
rect 102232 3868 102284 3874
rect 102232 3810 102284 3816
rect 102244 480 102272 3810
rect 103348 480 103376 7482
rect 103532 5098 103744 5114
rect 103520 5092 103756 5098
rect 103572 5086 103704 5092
rect 103520 5034 103572 5040
rect 103704 5034 103756 5040
rect 101006 354 101118 480
rect 100772 326 101118 354
rect 101006 -960 101118 326
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104084 354 104112 16546
rect 106464 11824 106516 11830
rect 106464 11766 106516 11772
rect 105728 6588 105780 6594
rect 105728 6530 105780 6536
rect 105740 480 105768 6530
rect 104502 354 104614 480
rect 104084 326 104614 354
rect 104502 -960 104614 326
rect 105698 -960 105810 480
rect 106476 354 106504 11766
rect 108132 480 108160 16546
rect 109314 7712 109370 7721
rect 109314 7647 109370 7656
rect 109328 480 109356 7647
rect 110432 3466 110460 78134
rect 111798 76800 111854 76809
rect 111798 76735 111854 76744
rect 111812 16574 111840 76735
rect 111812 16546 112392 16574
rect 110510 10296 110566 10305
rect 110510 10231 110566 10240
rect 110420 3460 110472 3466
rect 110420 3402 110472 3408
rect 110524 480 110552 10231
rect 111616 3460 111668 3466
rect 111616 3402 111668 3408
rect 111628 480 111656 3402
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112364 354 112392 16546
rect 113836 5166 113864 78202
rect 116584 77852 116636 77858
rect 116584 77794 116636 77800
rect 114560 72684 114612 72690
rect 114560 72626 114612 72632
rect 114572 16574 114600 72626
rect 115940 68332 115992 68338
rect 115940 68274 115992 68280
rect 115952 16574 115980 68274
rect 116596 37942 116624 77794
rect 116584 37936 116636 37942
rect 116584 37878 116636 37884
rect 118344 22778 118372 82175
rect 118436 80617 118464 86663
rect 118606 85232 118662 85241
rect 118606 85167 118662 85176
rect 118514 83736 118570 83745
rect 118514 83671 118570 83680
rect 118422 80608 118478 80617
rect 118422 80543 118478 80552
rect 118528 46918 118556 83671
rect 118620 80782 118648 85167
rect 118608 80776 118660 80782
rect 118608 80718 118660 80724
rect 119356 79529 119384 700266
rect 120724 616888 120776 616894
rect 120724 616830 120776 616836
rect 120736 102105 120764 616830
rect 120816 563100 120868 563106
rect 120816 563042 120868 563048
rect 120722 102096 120778 102105
rect 120722 102031 120778 102040
rect 120828 100745 120856 563042
rect 120908 510672 120960 510678
rect 120908 510614 120960 510620
rect 120814 100736 120870 100745
rect 120814 100671 120870 100680
rect 120920 98705 120948 510614
rect 121000 456816 121052 456822
rect 121000 456758 121052 456764
rect 120906 98696 120962 98705
rect 120906 98631 120962 98640
rect 121012 97209 121040 456758
rect 124864 298172 124916 298178
rect 124864 298114 124916 298120
rect 121092 292596 121144 292602
rect 121092 292538 121144 292544
rect 120998 97200 121054 97209
rect 120998 97135 121054 97144
rect 121104 80034 121132 292538
rect 123680 228410 123708 230588
rect 123668 228404 123720 228410
rect 123668 228346 123720 228352
rect 121184 187740 121236 187746
rect 121184 187682 121236 187688
rect 121092 80028 121144 80034
rect 121092 79970 121144 79976
rect 121196 79694 121224 187682
rect 122840 178832 122892 178838
rect 122840 178774 122892 178780
rect 121460 178696 121512 178702
rect 121460 178638 121512 178644
rect 121472 139890 121500 178638
rect 122104 165640 122156 165646
rect 122104 165582 122156 165588
rect 121472 139862 121808 139890
rect 122116 139534 122144 165582
rect 122852 151814 122880 178774
rect 124220 177336 124272 177342
rect 124220 177278 124272 177284
rect 124232 151814 124260 177278
rect 122852 151786 122972 151814
rect 124232 151786 124536 151814
rect 122944 139890 122972 151786
rect 124508 139890 124536 151786
rect 124876 142186 124904 298114
rect 129004 244316 129056 244322
rect 129004 244258 129056 244264
rect 126244 205692 126296 205698
rect 126244 205634 126296 205640
rect 125600 176044 125652 176050
rect 125600 175986 125652 175992
rect 125612 151814 125640 175986
rect 125612 151786 126100 151814
rect 124864 142180 124916 142186
rect 124864 142122 124916 142128
rect 126072 139890 126100 151786
rect 126256 140282 126284 205634
rect 128360 175976 128412 175982
rect 128360 175918 128412 175924
rect 126980 173256 127032 173262
rect 126980 173198 127032 173204
rect 126992 151814 127020 173198
rect 128372 151814 128400 175918
rect 126992 151786 127664 151814
rect 128372 151786 128952 151814
rect 126244 140276 126296 140282
rect 126244 140218 126296 140224
rect 127636 139890 127664 151786
rect 128924 140026 128952 151786
rect 129016 141574 129044 244258
rect 151832 230574 152582 230602
rect 143540 228404 143592 228410
rect 143540 228346 143592 228352
rect 138664 227792 138716 227798
rect 138664 227734 138716 227740
rect 138676 196790 138704 227734
rect 143552 200705 143580 228346
rect 151832 208418 151860 230574
rect 144920 208412 144972 208418
rect 144920 208354 144972 208360
rect 151820 208412 151872 208418
rect 151820 208354 151872 208360
rect 143538 200696 143594 200705
rect 143538 200631 143594 200640
rect 138664 196784 138716 196790
rect 138664 196726 138716 196732
rect 144932 196466 144960 208354
rect 146208 203584 146260 203590
rect 146208 203526 146260 203532
rect 144932 196438 145774 196466
rect 138112 195968 138164 195974
rect 138112 195910 138164 195916
rect 139398 195936 139454 195945
rect 138124 195809 138152 195910
rect 139398 195871 139400 195880
rect 139452 195871 139454 195880
rect 142342 195936 142398 195945
rect 142398 195894 142554 195922
rect 142342 195871 142398 195880
rect 139400 195842 139452 195848
rect 146220 195809 146248 203526
rect 147404 202156 147456 202162
rect 147404 202098 147456 202104
rect 147416 196452 147444 202098
rect 153856 196722 153884 702406
rect 161388 229764 161440 229770
rect 161388 229706 161440 229712
rect 154120 204944 154172 204950
rect 154120 204886 154172 204892
rect 153844 196716 153896 196722
rect 153844 196658 153896 196664
rect 152464 196512 152516 196518
rect 152214 196460 152464 196466
rect 152214 196454 152516 196460
rect 152214 196438 152504 196454
rect 153198 196208 153254 196217
rect 153198 196143 153254 196152
rect 138110 195800 138166 195809
rect 138110 195735 138166 195744
rect 140778 195800 140834 195809
rect 146206 195800 146262 195809
rect 140834 195758 140990 195786
rect 140778 195735 140834 195744
rect 146206 195735 146262 195744
rect 148784 195696 148836 195702
rect 148784 195638 148836 195644
rect 148796 194721 148824 195638
rect 148782 194712 148838 194721
rect 148782 194647 148838 194656
rect 153212 193633 153240 196143
rect 154132 195974 154160 204886
rect 159180 199436 159232 199442
rect 159180 199378 159232 199384
rect 154580 198076 154632 198082
rect 154580 198018 154632 198024
rect 154592 196518 154620 198018
rect 157340 198008 157392 198014
rect 157340 197950 157392 197956
rect 157248 196648 157300 196654
rect 157248 196590 157300 196596
rect 154580 196512 154632 196518
rect 154580 196454 154632 196460
rect 153476 195968 153528 195974
rect 153474 195936 153476 195945
rect 154120 195968 154172 195974
rect 153528 195936 153530 195945
rect 153934 195936 153990 195945
rect 153778 195894 153934 195922
rect 153474 195871 153530 195880
rect 157260 195945 157288 196590
rect 154120 195910 154172 195916
rect 157246 195936 157302 195945
rect 153934 195871 153990 195880
rect 157246 195871 157302 195880
rect 157154 195528 157210 195537
rect 157352 195514 157380 197950
rect 158902 195936 158958 195945
rect 158562 195894 158902 195922
rect 158902 195871 158958 195880
rect 159192 195809 159220 199378
rect 161400 195945 161428 229706
rect 166264 228404 166316 228410
rect 166264 228346 166316 228352
rect 166276 198082 166304 228346
rect 166264 198076 166316 198082
rect 166264 198018 166316 198024
rect 164240 196784 164292 196790
rect 164240 196726 164292 196732
rect 161386 195936 161442 195945
rect 161386 195871 161442 195880
rect 159178 195800 159234 195809
rect 159178 195735 159234 195744
rect 157210 195486 157380 195514
rect 157154 195463 157210 195472
rect 151450 193624 151506 193633
rect 151450 193559 151506 193568
rect 153198 193624 153254 193633
rect 153198 193559 153254 193568
rect 151464 191146 151492 193559
rect 151452 191140 151504 191146
rect 151452 191082 151504 191088
rect 148782 191040 148838 191049
rect 148782 190975 148838 190984
rect 148796 190876 148824 190975
rect 149794 190632 149850 190641
rect 149638 190590 149794 190618
rect 149794 190567 149850 190576
rect 164252 189394 164280 196726
rect 165434 196344 165490 196353
rect 165434 196279 165490 196288
rect 164252 189366 164634 189394
rect 144642 186960 144698 186969
rect 144578 186918 144642 186946
rect 144642 186895 144698 186904
rect 162136 184198 162426 184226
rect 136836 182974 137494 183002
rect 136836 180334 136864 182974
rect 137020 182022 137494 182050
rect 136824 180328 136876 180334
rect 136824 180270 136876 180276
rect 136640 180124 136692 180130
rect 136640 180066 136692 180072
rect 136652 178838 136680 180066
rect 136640 178832 136692 178838
rect 136640 178774 136692 178780
rect 137020 178702 137048 182022
rect 141252 180130 141280 181084
rect 162136 180946 162164 184198
rect 162124 180940 162176 180946
rect 162124 180882 162176 180888
rect 144460 180736 144512 180742
rect 146116 180736 146168 180742
rect 144460 180678 144512 180684
rect 146114 180704 146116 180713
rect 146168 180704 146170 180713
rect 144472 180676 144500 180678
rect 146114 180639 146170 180648
rect 161480 180600 161532 180606
rect 161480 180542 161532 180548
rect 141240 180124 141292 180130
rect 141240 180066 141292 180072
rect 137112 179982 137494 180010
rect 137008 178696 137060 178702
rect 137008 178638 137060 178644
rect 137112 177342 137140 179982
rect 143540 179648 143592 179654
rect 143540 179590 143592 179596
rect 143552 179588 143580 179590
rect 137204 179030 137494 179058
rect 137100 177336 137152 177342
rect 137100 177278 137152 177284
rect 137204 176050 137232 179030
rect 140792 177886 140820 179452
rect 148046 179072 148102 179081
rect 147982 179030 148046 179058
rect 148046 179007 148102 179016
rect 142666 178800 142722 178809
rect 142666 178735 142722 178744
rect 144184 178696 144236 178702
rect 144184 178638 144236 178644
rect 140780 177880 140832 177886
rect 140780 177822 140832 177828
rect 141608 177880 141660 177886
rect 141608 177822 141660 177828
rect 137296 176990 137494 177018
rect 137192 176044 137244 176050
rect 137192 175986 137244 175992
rect 137296 175982 137324 176990
rect 137388 176038 137494 176066
rect 137284 175976 137336 175982
rect 137284 175918 137336 175924
rect 135258 174040 135314 174049
rect 135258 173975 135314 173984
rect 135272 173942 135300 173975
rect 133880 173936 133932 173942
rect 133880 173878 133932 173884
rect 135260 173936 135312 173942
rect 135260 173878 135312 173884
rect 131120 173324 131172 173330
rect 131120 173266 131172 173272
rect 129004 141568 129056 141574
rect 129004 141510 129056 141516
rect 128924 139998 129228 140026
rect 129200 139890 129228 139998
rect 131132 139890 131160 173266
rect 132500 172236 132552 172242
rect 132500 172178 132552 172184
rect 132512 139890 132540 172178
rect 133892 139890 133920 173878
rect 137388 173330 137416 176038
rect 137376 173324 137428 173330
rect 137376 173266 137428 173272
rect 135260 172440 135312 172446
rect 135260 172382 135312 172388
rect 135272 151814 135300 172382
rect 137480 172242 137508 174964
rect 137834 174040 137890 174049
rect 137890 173998 137954 174026
rect 137834 173975 137890 173984
rect 141620 173874 141648 177822
rect 142066 176760 142122 176769
rect 142066 176695 142122 176704
rect 140780 173868 140832 173874
rect 140780 173810 140832 173816
rect 141608 173868 141660 173874
rect 141608 173810 141660 173816
rect 138952 172446 138980 173740
rect 139412 173726 139978 173754
rect 138940 172440 138992 172446
rect 138940 172382 138992 172388
rect 137468 172236 137520 172242
rect 137468 172178 137520 172184
rect 138020 171420 138072 171426
rect 138020 171362 138072 171368
rect 138032 151814 138060 171362
rect 135272 151786 135484 151814
rect 138032 151786 138612 151814
rect 135456 139890 135484 151786
rect 137744 143200 137796 143206
rect 137744 143142 137796 143148
rect 137756 139890 137784 143142
rect 122944 139862 123372 139890
rect 124508 139862 124936 139890
rect 126072 139862 126500 139890
rect 127636 139862 128064 139890
rect 129200 139862 129628 139890
rect 131132 139862 131192 139890
rect 132512 139862 132756 139890
rect 133892 139862 134320 139890
rect 135456 139862 135884 139890
rect 137448 139862 137784 139890
rect 138584 139890 138612 151786
rect 139412 143206 139440 173726
rect 140792 173262 140820 173810
rect 140780 173256 140832 173262
rect 140780 173198 140832 173204
rect 140976 171426 141004 173740
rect 141252 173726 142002 173754
rect 140964 171420 141016 171426
rect 140964 171362 141016 171368
rect 141252 161474 141280 173726
rect 142080 171193 142108 176695
rect 144196 174593 144224 178638
rect 161492 178106 161520 180542
rect 161400 178078 161520 178106
rect 161400 176254 161428 178078
rect 161388 176248 161440 176254
rect 161388 176190 161440 176196
rect 159088 175636 159140 175642
rect 159088 175578 159140 175584
rect 144182 174584 144238 174593
rect 144182 174519 144238 174528
rect 156050 174584 156106 174593
rect 156050 174519 156106 174528
rect 145562 173904 145618 173913
rect 145618 173862 145958 173890
rect 145562 173839 145618 173848
rect 142710 173768 142766 173777
rect 148690 173768 148746 173777
rect 142766 173726 142922 173754
rect 142710 173703 142766 173712
rect 142066 171184 142122 171193
rect 142066 171119 142122 171128
rect 142066 171048 142122 171057
rect 142066 170983 142122 170992
rect 142080 162217 142108 170983
rect 142066 162208 142122 162217
rect 142066 162143 142122 162152
rect 140976 161446 141280 161474
rect 139400 143200 139452 143206
rect 139400 143142 139452 143148
rect 140976 142154 141004 161446
rect 143538 142488 143594 142497
rect 143538 142423 143594 142432
rect 140700 142126 141004 142154
rect 142066 142216 142122 142225
rect 142066 142151 142122 142160
rect 140700 139890 140728 142126
rect 138584 139862 139012 139890
rect 140576 139862 140728 139890
rect 142080 139890 142108 142151
rect 143552 139890 143580 142423
rect 144932 139890 144960 173740
rect 146772 173726 146970 173754
rect 146772 173641 146800 173726
rect 148746 173726 148994 173754
rect 149072 173726 149914 173754
rect 150452 173726 150926 173754
rect 152476 173726 152950 173754
rect 148690 173703 148746 173712
rect 146758 173632 146814 173641
rect 146758 173567 146814 173576
rect 146482 143440 146538 143449
rect 146482 143375 146538 143384
rect 146496 139890 146524 143375
rect 148046 143304 148102 143313
rect 148046 143239 148102 143248
rect 148060 139890 148088 143239
rect 149072 142186 149100 173726
rect 149610 143168 149666 143177
rect 149610 143103 149666 143112
rect 149060 142180 149112 142186
rect 149060 142122 149112 142128
rect 149624 139890 149652 143103
rect 150452 142934 150480 173726
rect 152476 161474 152504 173726
rect 151832 161446 152504 161474
rect 151832 143546 151860 161446
rect 151820 143540 151872 143546
rect 151820 143482 151872 143488
rect 151174 143032 151230 143041
rect 151174 142967 151230 142976
rect 151358 143032 151414 143041
rect 151358 142967 151414 142976
rect 150440 142928 150492 142934
rect 150440 142870 150492 142876
rect 151188 139890 151216 142967
rect 151372 142633 151400 142967
rect 154580 142928 154632 142934
rect 154580 142870 154632 142876
rect 151358 142624 151414 142633
rect 151358 142559 151414 142568
rect 152740 142180 152792 142186
rect 152740 142122 152792 142128
rect 152752 139890 152780 142122
rect 154592 139890 154620 142870
rect 156064 139890 156092 174519
rect 157432 143540 157484 143546
rect 157432 143482 157484 143488
rect 157444 139890 157472 143482
rect 159100 139890 159128 175578
rect 165448 175030 165476 196279
rect 166170 196208 166226 196217
rect 166170 196143 166226 196152
rect 166078 196072 166134 196081
rect 166078 196007 166134 196016
rect 165528 195696 165580 195702
rect 165528 195638 165580 195644
rect 165540 175030 165568 195638
rect 165436 175024 165488 175030
rect 165436 174966 165488 174972
rect 165528 175024 165580 175030
rect 165528 174966 165580 174972
rect 163136 174752 163188 174758
rect 163136 174694 163188 174700
rect 165436 174752 165488 174758
rect 165436 174694 165488 174700
rect 165528 174752 165580 174758
rect 165528 174694 165580 174700
rect 162860 164756 162912 164762
rect 162860 164698 162912 164704
rect 162768 143268 162820 143274
rect 162768 143210 162820 143216
rect 160558 143032 160614 143041
rect 160558 142967 160614 142976
rect 160572 139890 160600 142967
rect 162780 139890 162808 143210
rect 162872 142934 162900 164698
rect 162860 142928 162912 142934
rect 162860 142870 162912 142876
rect 163148 142866 163176 174694
rect 163608 173726 163990 173754
rect 164252 173726 165002 173754
rect 163608 164762 163636 173726
rect 163596 164756 163648 164762
rect 163596 164698 163648 164704
rect 164056 143540 164108 143546
rect 164056 143482 164108 143488
rect 163136 142860 163188 142866
rect 163136 142802 163188 142808
rect 164068 140162 164096 143482
rect 164252 143002 164280 173726
rect 164330 166424 164386 166433
rect 164330 166359 164386 166368
rect 164344 151814 164372 166359
rect 165448 162858 165476 174694
rect 165540 164218 165568 174694
rect 165528 164212 165580 164218
rect 165528 164154 165580 164160
rect 165436 162852 165488 162858
rect 165436 162794 165488 162800
rect 164344 151786 165200 151814
rect 164240 142996 164292 143002
rect 164240 142938 164292 142944
rect 142080 139862 142140 139890
rect 143552 139862 143704 139890
rect 144932 139862 145268 139890
rect 146496 139862 146832 139890
rect 148060 139862 148396 139890
rect 149624 139862 149960 139890
rect 151188 139862 151524 139890
rect 152752 139862 153088 139890
rect 154592 139862 154652 139890
rect 156064 139862 156216 139890
rect 157444 139862 157780 139890
rect 159100 139862 159344 139890
rect 160572 139862 160908 139890
rect 162472 139862 162808 139890
rect 164022 140134 164096 140162
rect 164022 139876 164050 140134
rect 165172 139890 165200 151786
rect 166092 143274 166120 196007
rect 166184 143546 166212 196143
rect 166998 166288 167054 166297
rect 166998 166223 167054 166232
rect 166172 143540 166224 143546
rect 166172 143482 166224 143488
rect 166080 143268 166132 143274
rect 166080 143210 166132 143216
rect 167012 139890 167040 166223
rect 168380 164212 168432 164218
rect 168380 164154 168432 164160
rect 168392 139890 168420 164154
rect 169772 141506 169800 702406
rect 196624 700664 196676 700670
rect 196624 700606 196676 700612
rect 193864 700596 193916 700602
rect 193864 700538 193916 700544
rect 192484 700528 192536 700534
rect 192484 700470 192536 700476
rect 189724 700460 189776 700466
rect 189724 700402 189776 700408
rect 182548 700392 182600 700398
rect 182548 700334 182600 700340
rect 188344 700392 188396 700398
rect 188344 700334 188396 700340
rect 180800 700324 180852 700330
rect 180800 700266 180852 700272
rect 179420 462392 179472 462398
rect 179420 462334 179472 462340
rect 178684 305040 178736 305046
rect 178684 304982 178736 304988
rect 169852 162852 169904 162858
rect 169852 162794 169904 162800
rect 169760 141500 169812 141506
rect 169760 141442 169812 141448
rect 169864 139890 169892 162794
rect 176200 142996 176252 143002
rect 176200 142938 176252 142944
rect 174636 142928 174688 142934
rect 171506 142896 171562 142905
rect 174636 142870 174688 142876
rect 171506 142831 171562 142840
rect 171520 139890 171548 142831
rect 173070 142760 173126 142769
rect 173070 142695 173126 142704
rect 173084 139890 173112 142695
rect 174648 139890 174676 142870
rect 176212 139890 176240 142938
rect 178040 142860 178092 142866
rect 178040 142802 178092 142808
rect 178052 139890 178080 142802
rect 165172 139862 165600 139890
rect 167012 139862 167164 139890
rect 168392 139862 168728 139890
rect 169864 139862 170292 139890
rect 171520 139862 171856 139890
rect 173084 139862 173420 139890
rect 174648 139862 174984 139890
rect 176212 139862 176548 139890
rect 178052 139862 178112 139890
rect 122104 139528 122156 139534
rect 122104 139470 122156 139476
rect 178696 139330 178724 304982
rect 178776 253972 178828 253978
rect 178776 253914 178828 253920
rect 178788 139398 178816 253914
rect 178776 139392 178828 139398
rect 178776 139334 178828 139340
rect 178684 139324 178736 139330
rect 178684 139266 178736 139272
rect 179432 119377 179460 462334
rect 180064 271924 180116 271930
rect 180064 271866 180116 271872
rect 179604 201544 179656 201550
rect 179604 201486 179656 201492
rect 179512 139460 179564 139466
rect 179512 139402 179564 139408
rect 179524 128217 179552 139402
rect 179510 128208 179566 128217
rect 179510 128143 179566 128152
rect 179616 126177 179644 201486
rect 179696 173188 179748 173194
rect 179696 173130 179748 173136
rect 179602 126168 179658 126177
rect 179602 126103 179658 126112
rect 179418 119368 179474 119377
rect 179418 119303 179474 119312
rect 179708 116657 179736 173130
rect 179788 146940 179840 146946
rect 179788 146882 179840 146888
rect 179694 116648 179750 116657
rect 179694 116583 179750 116592
rect 179800 112577 179828 146882
rect 179878 130520 179934 130529
rect 179878 130455 179934 130464
rect 179786 112568 179842 112577
rect 179786 112503 179842 112512
rect 178592 80708 178644 80714
rect 178592 80650 178644 80656
rect 174636 80640 174688 80646
rect 174636 80582 174688 80588
rect 178040 80640 178092 80646
rect 178040 80582 178092 80588
rect 125416 80300 125468 80306
rect 125416 80242 125468 80248
rect 123482 80200 123538 80209
rect 123482 80135 123538 80144
rect 121184 79688 121236 79694
rect 121184 79630 121236 79636
rect 119342 79520 119398 79529
rect 119342 79455 119398 79464
rect 122194 78296 122250 78305
rect 122194 78231 122250 78240
rect 120816 77580 120868 77586
rect 120816 77522 120868 77528
rect 118700 76764 118752 76770
rect 118700 76706 118752 76712
rect 118516 46912 118568 46918
rect 118516 46854 118568 46860
rect 118332 22772 118384 22778
rect 118332 22714 118384 22720
rect 114572 16546 114784 16574
rect 115952 16546 116440 16574
rect 113824 5160 113876 5166
rect 113824 5102 113876 5108
rect 114008 5160 114060 5166
rect 114008 5102 114060 5108
rect 114020 480 114048 5102
rect 112782 354 112894 480
rect 112364 326 112894 354
rect 112782 -960 112894 326
rect 113978 -960 114090 480
rect 114756 354 114784 16546
rect 116412 480 116440 16546
rect 117320 10396 117372 10402
rect 117320 10338 117372 10344
rect 115174 354 115286 480
rect 114756 326 115286 354
rect 115174 -960 115286 326
rect 116370 -960 116482 480
rect 117332 354 117360 10338
rect 118712 3466 118740 76706
rect 120722 75848 120778 75857
rect 120722 75783 120778 75792
rect 119344 74044 119396 74050
rect 119344 73986 119396 73992
rect 118700 3460 118752 3466
rect 118700 3402 118752 3408
rect 119356 3398 119384 73986
rect 120080 60308 120132 60314
rect 120080 60250 120132 60256
rect 120092 16574 120120 60250
rect 120092 16546 120672 16574
rect 119896 3460 119948 3466
rect 119896 3402 119948 3408
rect 119344 3392 119396 3398
rect 119344 3334 119396 3340
rect 118792 3256 118844 3262
rect 118792 3198 118844 3204
rect 118804 480 118832 3198
rect 119908 480 119936 3402
rect 117566 354 117678 480
rect 117332 326 117678 354
rect 117566 -960 117678 326
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 120644 354 120672 16546
rect 120736 3670 120764 75783
rect 120828 32434 120856 77522
rect 122102 74488 122158 74497
rect 122102 74423 122158 74432
rect 121460 71460 121512 71466
rect 121460 71402 121512 71408
rect 120816 32428 120868 32434
rect 120816 32370 120868 32376
rect 121472 16574 121500 71402
rect 121472 16546 122052 16574
rect 120724 3664 120776 3670
rect 120724 3606 120776 3612
rect 122024 3482 122052 16546
rect 122116 3602 122144 74423
rect 122208 7614 122236 78231
rect 122380 77648 122432 77654
rect 122380 77590 122432 77596
rect 122288 72752 122340 72758
rect 122288 72694 122340 72700
rect 122300 16574 122328 72694
rect 122392 35222 122420 77590
rect 122840 76832 122892 76838
rect 122840 76774 122892 76780
rect 122380 35216 122432 35222
rect 122380 35158 122432 35164
rect 122852 16574 122880 76774
rect 122300 16546 122420 16574
rect 122852 16546 123064 16574
rect 122196 7608 122248 7614
rect 122196 7550 122248 7556
rect 122392 3738 122420 16546
rect 122380 3732 122432 3738
rect 122380 3674 122432 3680
rect 122104 3596 122156 3602
rect 122104 3538 122156 3544
rect 122024 3454 122328 3482
rect 122300 480 122328 3454
rect 121062 354 121174 480
rect 120644 326 121174 354
rect 121062 -960 121174 326
rect 122258 -960 122370 480
rect 123036 354 123064 16546
rect 123496 3806 123524 80135
rect 125232 80096 125284 80102
rect 125232 80038 125284 80044
rect 123852 80028 123904 80034
rect 123852 79970 123904 79976
rect 123576 79756 123628 79762
rect 123576 79698 123628 79704
rect 123588 79354 123616 79698
rect 123576 79348 123628 79354
rect 123576 79290 123628 79296
rect 123668 78464 123720 78470
rect 123668 78406 123720 78412
rect 123576 75472 123628 75478
rect 123576 75414 123628 75420
rect 123484 3800 123536 3806
rect 123484 3742 123536 3748
rect 123588 3262 123616 75414
rect 123680 60314 123708 78406
rect 123864 76537 123892 79970
rect 124956 79960 125008 79966
rect 124956 79902 125008 79908
rect 124772 79824 124824 79830
rect 124772 79766 124824 79772
rect 124036 78668 124088 78674
rect 124036 78610 124088 78616
rect 123850 76528 123906 76537
rect 123850 76463 123906 76472
rect 124048 75070 124076 78610
rect 124036 75064 124088 75070
rect 124036 75006 124088 75012
rect 124784 70394 124812 79766
rect 124864 76424 124916 76430
rect 124864 76366 124916 76372
rect 124232 70366 124812 70394
rect 123668 60308 123720 60314
rect 123668 60250 123720 60256
rect 124232 36582 124260 70366
rect 124220 36576 124272 36582
rect 124220 36518 124272 36524
rect 124220 20052 124272 20058
rect 124220 19994 124272 20000
rect 124232 16574 124260 19994
rect 124232 16546 124720 16574
rect 123576 3256 123628 3262
rect 123576 3198 123628 3204
rect 124692 480 124720 16546
rect 124876 3874 124904 76366
rect 124864 3868 124916 3874
rect 124864 3810 124916 3816
rect 124968 3534 124996 79902
rect 125244 77654 125272 80038
rect 125428 79694 125456 80242
rect 174452 80232 174504 80238
rect 174452 80174 174504 80180
rect 125566 79971 125594 80036
rect 125552 79962 125608 79971
rect 125552 79897 125608 79906
rect 125658 79812 125686 80036
rect 125750 79971 125778 80036
rect 125736 79962 125792 79971
rect 125736 79897 125792 79906
rect 125842 79898 125870 80036
rect 125934 79971 125962 80036
rect 125920 79962 125976 79971
rect 125830 79892 125882 79898
rect 125920 79897 125976 79906
rect 126026 79898 126054 80036
rect 126118 79966 126146 80036
rect 126210 79966 126238 80036
rect 126106 79960 126158 79966
rect 126106 79902 126158 79908
rect 126198 79960 126250 79966
rect 126198 79902 126250 79908
rect 126302 79898 126330 80036
rect 126394 79966 126422 80036
rect 126382 79960 126434 79966
rect 126382 79902 126434 79908
rect 125830 79834 125882 79840
rect 126014 79892 126066 79898
rect 126014 79834 126066 79840
rect 126290 79892 126342 79898
rect 126290 79834 126342 79840
rect 125738 79824 125790 79830
rect 125658 79784 125738 79812
rect 125738 79766 125790 79772
rect 125874 79792 125930 79801
rect 125874 79727 125930 79736
rect 126244 79756 126296 79762
rect 125416 79688 125468 79694
rect 125600 79688 125652 79694
rect 125416 79630 125468 79636
rect 125598 79656 125600 79665
rect 125692 79688 125744 79694
rect 125652 79656 125654 79665
rect 125692 79630 125744 79636
rect 125782 79656 125838 79665
rect 125598 79591 125654 79600
rect 125508 79484 125560 79490
rect 125508 79426 125560 79432
rect 125324 77920 125376 77926
rect 125324 77862 125376 77868
rect 125232 77648 125284 77654
rect 125232 77590 125284 77596
rect 125232 77376 125284 77382
rect 125232 77318 125284 77324
rect 125140 76288 125192 76294
rect 125140 76230 125192 76236
rect 125048 76084 125100 76090
rect 125048 76026 125100 76032
rect 125060 6254 125088 76026
rect 125152 51746 125180 76230
rect 125244 55894 125272 77318
rect 125336 57254 125364 77862
rect 125416 77716 125468 77722
rect 125416 77658 125468 77664
rect 125428 61402 125456 77658
rect 125520 75342 125548 79426
rect 125600 79212 125652 79218
rect 125600 79154 125652 79160
rect 125612 78577 125640 79154
rect 125704 78713 125732 79630
rect 125782 79591 125838 79600
rect 125690 78704 125746 78713
rect 125690 78639 125746 78648
rect 125598 78568 125654 78577
rect 125598 78503 125654 78512
rect 125692 77444 125744 77450
rect 125692 77386 125744 77392
rect 125508 75336 125560 75342
rect 125508 75278 125560 75284
rect 125704 70394 125732 77386
rect 125796 75857 125824 79591
rect 125888 78334 125916 79727
rect 126244 79698 126296 79704
rect 126336 79756 126388 79762
rect 126336 79698 126388 79704
rect 125968 79688 126020 79694
rect 125968 79630 126020 79636
rect 125980 78849 126008 79630
rect 126060 79620 126112 79626
rect 126060 79562 126112 79568
rect 126152 79620 126204 79626
rect 126152 79562 126204 79568
rect 125966 78840 126022 78849
rect 125966 78775 126022 78784
rect 125968 78736 126020 78742
rect 125968 78678 126020 78684
rect 125876 78328 125928 78334
rect 125876 78270 125928 78276
rect 125876 77240 125928 77246
rect 125876 77182 125928 77188
rect 125782 75848 125838 75857
rect 125782 75783 125838 75792
rect 125784 75540 125836 75546
rect 125784 75482 125836 75488
rect 125612 70366 125732 70394
rect 125416 61396 125468 61402
rect 125416 61338 125468 61344
rect 125324 57248 125376 57254
rect 125324 57190 125376 57196
rect 125232 55888 125284 55894
rect 125232 55830 125284 55836
rect 125140 51740 125192 51746
rect 125140 51682 125192 51688
rect 125048 6248 125100 6254
rect 125048 6190 125100 6196
rect 124956 3528 125008 3534
rect 124956 3470 125008 3476
rect 123454 354 123566 480
rect 123036 326 123566 354
rect 123454 -960 123566 326
rect 124650 -960 124762 480
rect 125612 354 125640 70366
rect 125796 4894 125824 75482
rect 125888 6186 125916 77182
rect 125980 22914 126008 78678
rect 126072 77897 126100 79562
rect 126164 78538 126192 79562
rect 126152 78532 126204 78538
rect 126152 78474 126204 78480
rect 126256 78418 126284 79698
rect 126348 78742 126376 79698
rect 126486 79540 126514 80036
rect 126578 79642 126606 80036
rect 126670 79812 126698 80036
rect 126762 79937 126790 80036
rect 126854 79966 126882 80036
rect 126946 79971 126974 80036
rect 126842 79960 126894 79966
rect 126748 79928 126804 79937
rect 126842 79902 126894 79908
rect 126932 79962 126988 79971
rect 126932 79897 126988 79906
rect 126748 79863 126804 79872
rect 127038 79830 127066 80036
rect 127026 79824 127078 79830
rect 126670 79784 126744 79812
rect 126578 79614 126652 79642
rect 126486 79512 126560 79540
rect 126336 78736 126388 78742
rect 126336 78678 126388 78684
rect 126336 78532 126388 78538
rect 126336 78474 126388 78480
rect 126164 78390 126284 78418
rect 126058 77888 126114 77897
rect 126058 77823 126114 77832
rect 126164 70394 126192 78390
rect 126244 77308 126296 77314
rect 126244 77250 126296 77256
rect 126072 70366 126192 70394
rect 125968 22908 126020 22914
rect 125968 22850 126020 22856
rect 126072 22846 126100 70366
rect 126060 22840 126112 22846
rect 126060 22782 126112 22788
rect 126256 8974 126284 77250
rect 126348 70394 126376 78474
rect 126532 71058 126560 79512
rect 126624 75546 126652 79614
rect 126716 76294 126744 79784
rect 126886 79792 126942 79801
rect 126808 79750 126886 79778
rect 126808 77246 126836 79750
rect 127130 79801 127158 80036
rect 127222 79966 127250 80036
rect 127314 79966 127342 80036
rect 127406 79971 127434 80036
rect 127210 79960 127262 79966
rect 127210 79902 127262 79908
rect 127302 79960 127354 79966
rect 127302 79902 127354 79908
rect 127392 79962 127448 79971
rect 127498 79966 127526 80036
rect 127590 79966 127618 80036
rect 127682 79966 127710 80036
rect 127774 79971 127802 80036
rect 127392 79897 127448 79906
rect 127486 79960 127538 79966
rect 127486 79902 127538 79908
rect 127578 79960 127630 79966
rect 127578 79902 127630 79908
rect 127670 79960 127722 79966
rect 127670 79902 127722 79908
rect 127760 79962 127816 79971
rect 127866 79966 127894 80036
rect 127760 79897 127816 79906
rect 127854 79960 127906 79966
rect 127854 79902 127906 79908
rect 127958 79898 127986 80036
rect 128050 79971 128078 80036
rect 128036 79962 128092 79971
rect 128142 79966 128170 80036
rect 127946 79892 127998 79898
rect 128036 79897 128092 79906
rect 128130 79960 128182 79966
rect 128130 79902 128182 79908
rect 127946 79834 127998 79840
rect 127578 79824 127630 79830
rect 127026 79766 127078 79772
rect 127116 79792 127172 79801
rect 126886 79727 126942 79736
rect 127578 79766 127630 79772
rect 127714 79792 127770 79801
rect 127116 79727 127172 79736
rect 127256 79756 127308 79762
rect 127256 79698 127308 79704
rect 126888 79688 126940 79694
rect 126888 79630 126940 79636
rect 126980 79688 127032 79694
rect 126980 79630 127032 79636
rect 127164 79688 127216 79694
rect 127164 79630 127216 79636
rect 126796 77240 126848 77246
rect 126796 77182 126848 77188
rect 126704 76288 126756 76294
rect 126704 76230 126756 76236
rect 126612 75540 126664 75546
rect 126612 75482 126664 75488
rect 126900 74534 126928 79630
rect 126992 76090 127020 79630
rect 127072 78396 127124 78402
rect 127072 78338 127124 78344
rect 126980 76084 127032 76090
rect 126980 76026 127032 76032
rect 126624 74506 126928 74534
rect 126624 71126 126652 74506
rect 126612 71120 126664 71126
rect 126612 71062 126664 71068
rect 126520 71052 126572 71058
rect 126520 70994 126572 71000
rect 127084 70394 127112 78338
rect 127176 77246 127204 79630
rect 127268 78713 127296 79698
rect 127590 79540 127618 79766
rect 127714 79727 127770 79736
rect 127900 79756 127952 79762
rect 127452 79512 127618 79540
rect 127254 78704 127310 78713
rect 127254 78639 127310 78648
rect 127452 78674 127480 79512
rect 127624 79212 127676 79218
rect 127624 79154 127676 79160
rect 127452 78646 127572 78674
rect 127346 78160 127402 78169
rect 127346 78095 127402 78104
rect 127164 77240 127216 77246
rect 127164 77182 127216 77188
rect 127360 70394 127388 78095
rect 127544 77246 127572 78646
rect 127440 77240 127492 77246
rect 127440 77182 127492 77188
rect 127532 77240 127584 77246
rect 127532 77182 127584 77188
rect 126348 70366 126468 70394
rect 126244 8968 126296 8974
rect 126244 8910 126296 8916
rect 125876 6180 125928 6186
rect 125876 6122 125928 6128
rect 125784 4888 125836 4894
rect 125784 4830 125836 4836
rect 126440 4826 126468 70366
rect 126992 70366 127112 70394
rect 127268 70366 127388 70394
rect 126428 4820 126480 4826
rect 126428 4762 126480 4768
rect 126992 480 127020 70366
rect 127268 7750 127296 70366
rect 127346 68232 127402 68241
rect 127346 68167 127402 68176
rect 127360 16574 127388 68167
rect 127452 24206 127480 77182
rect 127636 74534 127664 79154
rect 127544 74506 127664 74534
rect 127544 66910 127572 74506
rect 127532 66904 127584 66910
rect 127532 66846 127584 66852
rect 127440 24200 127492 24206
rect 127440 24142 127492 24148
rect 127360 16546 127664 16574
rect 127256 7744 127308 7750
rect 127256 7686 127308 7692
rect 127636 3482 127664 16546
rect 127728 4962 127756 79727
rect 127900 79698 127952 79704
rect 127992 79756 128044 79762
rect 127992 79698 128044 79704
rect 128084 79756 128136 79762
rect 128234 79744 128262 80036
rect 128326 79971 128354 80036
rect 128312 79962 128368 79971
rect 128312 79897 128368 79906
rect 128418 79830 128446 80036
rect 128406 79824 128458 79830
rect 128406 79766 128458 79772
rect 128510 79778 128538 80036
rect 128602 79966 128630 80036
rect 128590 79960 128642 79966
rect 128694 79937 128722 80036
rect 128786 79966 128814 80036
rect 128878 79966 128906 80036
rect 128970 79966 128998 80036
rect 128774 79960 128826 79966
rect 128590 79902 128642 79908
rect 128680 79928 128736 79937
rect 128774 79902 128826 79908
rect 128866 79960 128918 79966
rect 128866 79902 128918 79908
rect 128958 79960 129010 79966
rect 129062 79937 129090 80036
rect 128958 79902 129010 79908
rect 129048 79928 129104 79937
rect 128680 79863 128736 79872
rect 129154 79898 129182 80036
rect 129246 79966 129274 80036
rect 129234 79960 129286 79966
rect 129234 79902 129286 79908
rect 129048 79863 129104 79872
rect 129142 79892 129194 79898
rect 129142 79834 129194 79840
rect 128636 79824 128688 79830
rect 128510 79750 128584 79778
rect 128636 79766 128688 79772
rect 128728 79824 128780 79830
rect 128728 79766 128780 79772
rect 129094 79792 129150 79801
rect 128084 79698 128136 79704
rect 128188 79716 128262 79744
rect 127808 77240 127860 77246
rect 127808 77182 127860 77188
rect 127820 72486 127848 77182
rect 127912 73846 127940 79698
rect 128004 78606 128032 79698
rect 128096 79218 128124 79698
rect 128084 79212 128136 79218
rect 128084 79154 128136 79160
rect 128084 79076 128136 79082
rect 128084 79018 128136 79024
rect 128096 78674 128124 79018
rect 128084 78668 128136 78674
rect 128084 78610 128136 78616
rect 127992 78600 128044 78606
rect 127992 78542 128044 78548
rect 128084 77240 128136 77246
rect 128084 77182 128136 77188
rect 127900 73840 127952 73846
rect 127900 73782 127952 73788
rect 127808 72480 127860 72486
rect 127808 72422 127860 72428
rect 128096 71194 128124 77182
rect 128084 71188 128136 71194
rect 128084 71130 128136 71136
rect 128188 64874 128216 79716
rect 128360 79688 128412 79694
rect 128266 79656 128322 79665
rect 128360 79630 128412 79636
rect 128452 79688 128504 79694
rect 128452 79630 128504 79636
rect 128266 79591 128322 79600
rect 128280 77586 128308 79591
rect 128268 77580 128320 77586
rect 128268 77522 128320 77528
rect 128372 77246 128400 79630
rect 128464 77353 128492 79630
rect 128450 77344 128506 77353
rect 128450 77279 128506 77288
rect 128360 77240 128412 77246
rect 128360 77182 128412 77188
rect 128556 76673 128584 79750
rect 128648 79082 128676 79766
rect 128636 79076 128688 79082
rect 128636 79018 128688 79024
rect 128740 78169 128768 79766
rect 128820 79756 128872 79762
rect 129094 79727 129150 79736
rect 129338 79744 129366 80036
rect 129430 79812 129458 80036
rect 129522 79937 129550 80036
rect 129508 79928 129564 79937
rect 129508 79863 129564 79872
rect 129614 79830 129642 80036
rect 129602 79824 129654 79830
rect 129430 79784 129504 79812
rect 128820 79698 128872 79704
rect 128726 78160 128782 78169
rect 128726 78095 128782 78104
rect 128832 77330 128860 79698
rect 129108 79558 129136 79727
rect 129338 79716 129412 79744
rect 129188 79688 129240 79694
rect 129188 79630 129240 79636
rect 128912 79552 128964 79558
rect 128912 79494 128964 79500
rect 129096 79552 129148 79558
rect 129096 79494 129148 79500
rect 128648 77302 128860 77330
rect 128542 76664 128598 76673
rect 128542 76599 128598 76608
rect 128544 75540 128596 75546
rect 128544 75482 128596 75488
rect 128556 70394 128584 75482
rect 127820 64846 128216 64874
rect 128372 70366 128584 70394
rect 127820 7682 127848 64846
rect 128372 9042 128400 70366
rect 128648 22982 128676 77302
rect 128728 76152 128780 76158
rect 128728 76094 128780 76100
rect 128636 22976 128688 22982
rect 128636 22918 128688 22924
rect 128360 9036 128412 9042
rect 128360 8978 128412 8984
rect 127808 7676 127860 7682
rect 127808 7618 127860 7624
rect 128740 6322 128768 76094
rect 128818 75984 128874 75993
rect 128818 75919 128874 75928
rect 128832 7818 128860 75919
rect 128924 69698 128952 79494
rect 129096 79416 129148 79422
rect 129096 79358 129148 79364
rect 129108 79082 129136 79358
rect 129096 79076 129148 79082
rect 129096 79018 129148 79024
rect 129200 77858 129228 79630
rect 129280 79620 129332 79626
rect 129280 79562 129332 79568
rect 129188 77852 129240 77858
rect 129188 77794 129240 77800
rect 129096 77036 129148 77042
rect 129096 76978 129148 76984
rect 129108 69766 129136 76978
rect 129188 75744 129240 75750
rect 129188 75686 129240 75692
rect 129096 69760 129148 69766
rect 129096 69702 129148 69708
rect 128912 69692 128964 69698
rect 128912 69634 128964 69640
rect 129200 7886 129228 75686
rect 129292 75342 129320 79562
rect 129280 75336 129332 75342
rect 129280 75278 129332 75284
rect 129384 71262 129412 79716
rect 129476 79626 129504 79784
rect 129706 79801 129734 80036
rect 129798 79898 129826 80036
rect 129786 79892 129838 79898
rect 129786 79834 129838 79840
rect 129602 79766 129654 79772
rect 129692 79792 129748 79801
rect 129692 79727 129748 79736
rect 129556 79688 129608 79694
rect 129738 79656 129794 79665
rect 129556 79630 129608 79636
rect 129464 79620 129516 79626
rect 129464 79562 129516 79568
rect 129568 79472 129596 79630
rect 129476 79444 129596 79472
rect 129660 79614 129738 79642
rect 129476 76158 129504 79444
rect 129660 79370 129688 79614
rect 129738 79591 129794 79600
rect 129740 79552 129792 79558
rect 129890 79540 129918 80036
rect 129982 79971 130010 80036
rect 129968 79962 130024 79971
rect 129968 79897 130024 79906
rect 130074 79744 130102 80036
rect 130166 79966 130194 80036
rect 130258 79966 130286 80036
rect 130350 79966 130378 80036
rect 130442 79966 130470 80036
rect 130154 79960 130206 79966
rect 130154 79902 130206 79908
rect 130246 79960 130298 79966
rect 130246 79902 130298 79908
rect 130338 79960 130390 79966
rect 130338 79902 130390 79908
rect 130430 79960 130482 79966
rect 130430 79902 130482 79908
rect 130534 79778 130562 80036
rect 130626 79812 130654 80036
rect 130718 79971 130746 80036
rect 130704 79962 130760 79971
rect 130704 79897 130760 79906
rect 130706 79824 130758 79830
rect 130626 79784 130706 79812
rect 130200 79756 130252 79762
rect 130074 79716 130148 79744
rect 130120 79665 130148 79716
rect 130200 79698 130252 79704
rect 130292 79756 130344 79762
rect 130292 79698 130344 79704
rect 130488 79750 130562 79778
rect 130706 79766 130758 79772
rect 130106 79656 130162 79665
rect 130106 79591 130162 79600
rect 129890 79512 129964 79540
rect 129740 79494 129792 79500
rect 129568 79342 129688 79370
rect 129464 76152 129516 76158
rect 129464 76094 129516 76100
rect 129568 75750 129596 79342
rect 129648 79280 129700 79286
rect 129648 79222 129700 79228
rect 129660 78266 129688 79222
rect 129648 78260 129700 78266
rect 129648 78202 129700 78208
rect 129752 77994 129780 79494
rect 129832 79416 129884 79422
rect 129832 79358 129884 79364
rect 129740 77988 129792 77994
rect 129740 77930 129792 77936
rect 129740 76084 129792 76090
rect 129740 76026 129792 76032
rect 129556 75744 129608 75750
rect 129556 75686 129608 75692
rect 129372 71256 129424 71262
rect 129372 71198 129424 71204
rect 129188 7880 129240 7886
rect 129188 7822 129240 7828
rect 128820 7812 128872 7818
rect 128820 7754 128872 7760
rect 129752 6914 129780 76026
rect 129844 70394 129872 79358
rect 129936 78713 129964 79512
rect 130108 79416 130160 79422
rect 130108 79358 130160 79364
rect 129922 78704 129978 78713
rect 129922 78639 129978 78648
rect 130016 78532 130068 78538
rect 130016 78474 130068 78480
rect 129924 77852 129976 77858
rect 129924 77794 129976 77800
rect 129936 75546 129964 77794
rect 129924 75540 129976 75546
rect 129924 75482 129976 75488
rect 129844 70366 129964 70394
rect 129936 11762 129964 70366
rect 130028 19990 130056 78474
rect 130120 75478 130148 79358
rect 130212 78849 130240 79698
rect 130198 78840 130254 78849
rect 130198 78775 130254 78784
rect 130304 78674 130332 79698
rect 130488 79608 130516 79750
rect 130660 79688 130712 79694
rect 130658 79656 130660 79665
rect 130712 79656 130714 79665
rect 130810 79642 130838 80036
rect 130902 79966 130930 80036
rect 130994 79971 131022 80036
rect 130890 79960 130942 79966
rect 130890 79902 130942 79908
rect 130980 79962 131036 79971
rect 130980 79897 131036 79906
rect 131086 79898 131114 80036
rect 131074 79892 131126 79898
rect 131074 79834 131126 79840
rect 131028 79756 131080 79762
rect 131178 79744 131206 80036
rect 131270 79937 131298 80036
rect 131256 79928 131312 79937
rect 131256 79863 131312 79872
rect 131362 79744 131390 80036
rect 131454 79971 131482 80036
rect 131440 79962 131496 79971
rect 131440 79897 131496 79906
rect 131546 79744 131574 80036
rect 131178 79716 131252 79744
rect 131362 79716 131436 79744
rect 131028 79698 131080 79704
rect 130396 79580 130516 79608
rect 130568 79620 130620 79626
rect 130396 79014 130424 79580
rect 130658 79591 130714 79600
rect 130764 79614 130838 79642
rect 130568 79562 130620 79568
rect 130580 79370 130608 79562
rect 130488 79342 130608 79370
rect 130384 79008 130436 79014
rect 130384 78950 130436 78956
rect 130212 78646 130332 78674
rect 130212 77042 130240 78646
rect 130200 77036 130252 77042
rect 130200 76978 130252 76984
rect 130290 76528 130346 76537
rect 130290 76463 130346 76472
rect 130108 75472 130160 75478
rect 130108 75414 130160 75420
rect 130016 19984 130068 19990
rect 130016 19926 130068 19932
rect 129924 11756 129976 11762
rect 129924 11698 129976 11704
rect 129752 6886 130240 6914
rect 128728 6316 128780 6322
rect 128728 6258 128780 6264
rect 127716 4956 127768 4962
rect 127716 4898 127768 4904
rect 129372 3596 129424 3602
rect 129372 3538 129424 3544
rect 127636 3454 128216 3482
rect 128188 480 128216 3454
rect 129384 480 129412 3538
rect 130212 3482 130240 6886
rect 130304 5098 130332 76463
rect 130384 75812 130436 75818
rect 130384 75754 130436 75760
rect 130292 5092 130344 5098
rect 130292 5034 130344 5040
rect 130396 3602 130424 75754
rect 130488 74050 130516 79342
rect 130568 79008 130620 79014
rect 130568 78950 130620 78956
rect 130580 77314 130608 78950
rect 130658 78840 130714 78849
rect 130658 78775 130714 78784
rect 130568 77308 130620 77314
rect 130568 77250 130620 77256
rect 130672 74534 130700 78775
rect 130764 78538 130792 79614
rect 130844 79552 130896 79558
rect 130844 79494 130896 79500
rect 130752 78532 130804 78538
rect 130752 78474 130804 78480
rect 130580 74506 130700 74534
rect 130476 74044 130528 74050
rect 130476 73986 130528 73992
rect 130580 72758 130608 74506
rect 130856 73914 130884 79494
rect 130936 79484 130988 79490
rect 130936 79426 130988 79432
rect 130948 76702 130976 79426
rect 130936 76696 130988 76702
rect 130936 76638 130988 76644
rect 131040 76634 131068 79698
rect 131118 79656 131174 79665
rect 131118 79591 131174 79600
rect 131028 76628 131080 76634
rect 131028 76570 131080 76576
rect 131132 76566 131160 79591
rect 131120 76560 131172 76566
rect 131120 76502 131172 76508
rect 131028 76492 131080 76498
rect 131028 76434 131080 76440
rect 131040 73982 131068 76434
rect 131120 74044 131172 74050
rect 131120 73986 131172 73992
rect 131028 73976 131080 73982
rect 131028 73918 131080 73924
rect 130844 73908 130896 73914
rect 130844 73850 130896 73856
rect 130568 72752 130620 72758
rect 130568 72694 130620 72700
rect 131132 6914 131160 73986
rect 131224 73953 131252 79716
rect 131304 79620 131356 79626
rect 131304 79562 131356 79568
rect 131210 73944 131266 73953
rect 131210 73879 131266 73888
rect 131316 71330 131344 79562
rect 131408 76673 131436 79716
rect 131500 79716 131574 79744
rect 131638 79744 131666 80036
rect 131730 79966 131758 80036
rect 131718 79960 131770 79966
rect 131822 79937 131850 80036
rect 131718 79902 131770 79908
rect 131808 79928 131864 79937
rect 131808 79863 131864 79872
rect 131914 79812 131942 80036
rect 132006 79966 132034 80036
rect 131994 79960 132046 79966
rect 131994 79902 132046 79908
rect 131914 79784 131988 79812
rect 131638 79716 131712 79744
rect 131394 76664 131450 76673
rect 131394 76599 131450 76608
rect 131500 76514 131528 79716
rect 131578 79656 131634 79665
rect 131578 79591 131634 79600
rect 131408 76486 131528 76514
rect 131304 71324 131356 71330
rect 131304 71266 131356 71272
rect 131408 70394 131436 76486
rect 131592 76430 131620 79591
rect 131684 77858 131712 79716
rect 131856 79688 131908 79694
rect 131856 79630 131908 79636
rect 131672 77852 131724 77858
rect 131672 77794 131724 77800
rect 131670 76664 131726 76673
rect 131670 76599 131726 76608
rect 131764 76628 131816 76634
rect 131580 76424 131632 76430
rect 131580 76366 131632 76372
rect 131580 76288 131632 76294
rect 131580 76230 131632 76236
rect 131488 76016 131540 76022
rect 131488 75958 131540 75964
rect 131316 70366 131436 70394
rect 131316 16574 131344 70366
rect 131316 16546 131436 16574
rect 131132 6886 131344 6914
rect 130384 3596 130436 3602
rect 130384 3538 130436 3544
rect 130212 3454 130608 3482
rect 130580 480 130608 3454
rect 125846 354 125958 480
rect 125612 326 125958 354
rect 125846 -960 125958 326
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131316 354 131344 6886
rect 131408 6390 131436 16546
rect 131500 9110 131528 75958
rect 131592 44878 131620 76230
rect 131580 44872 131632 44878
rect 131580 44814 131632 44820
rect 131488 9104 131540 9110
rect 131488 9046 131540 9052
rect 131684 6458 131712 76599
rect 131764 76570 131816 76576
rect 131776 6526 131804 76570
rect 131868 69834 131896 79630
rect 131960 76294 131988 79784
rect 132098 79744 132126 80036
rect 132052 79716 132126 79744
rect 132052 76634 132080 79716
rect 132190 79676 132218 80036
rect 132282 79966 132310 80036
rect 132374 79971 132402 80036
rect 132270 79960 132322 79966
rect 132270 79902 132322 79908
rect 132360 79962 132416 79971
rect 132360 79897 132416 79906
rect 132466 79812 132494 80036
rect 132420 79784 132494 79812
rect 132316 79756 132368 79762
rect 132316 79698 132368 79704
rect 132144 79648 132218 79676
rect 132040 76628 132092 76634
rect 132040 76570 132092 76576
rect 131948 76288 132000 76294
rect 131948 76230 132000 76236
rect 132144 76022 132172 79648
rect 132224 79552 132276 79558
rect 132224 79494 132276 79500
rect 132132 76016 132184 76022
rect 132132 75958 132184 75964
rect 132236 75410 132264 79494
rect 132224 75404 132276 75410
rect 132224 75346 132276 75352
rect 132328 72554 132356 79698
rect 132420 77382 132448 79784
rect 132558 79744 132586 80036
rect 132650 79801 132678 80036
rect 132742 79937 132770 80036
rect 132728 79928 132784 79937
rect 132728 79863 132784 79872
rect 132834 79812 132862 80036
rect 132926 79966 132954 80036
rect 132914 79960 132966 79966
rect 132914 79902 132966 79908
rect 132512 79716 132586 79744
rect 132636 79792 132692 79801
rect 132636 79727 132692 79736
rect 132788 79784 132862 79812
rect 132512 78130 132540 79716
rect 132788 79506 132816 79784
rect 133018 79744 133046 80036
rect 133110 79812 133138 80036
rect 133202 79966 133230 80036
rect 133190 79960 133242 79966
rect 133190 79902 133242 79908
rect 133110 79784 133184 79812
rect 133018 79716 133092 79744
rect 132868 79688 132920 79694
rect 132868 79630 132920 79636
rect 132604 79478 132816 79506
rect 132500 78124 132552 78130
rect 132500 78066 132552 78072
rect 132408 77376 132460 77382
rect 132408 77318 132460 77324
rect 132408 76696 132460 76702
rect 132408 76638 132460 76644
rect 132316 72548 132368 72554
rect 132316 72490 132368 72496
rect 131856 69828 131908 69834
rect 131856 69770 131908 69776
rect 131764 6520 131816 6526
rect 131764 6462 131816 6468
rect 131672 6452 131724 6458
rect 131672 6394 131724 6400
rect 131396 6384 131448 6390
rect 131396 6326 131448 6332
rect 132420 6118 132448 76638
rect 132604 76498 132632 79478
rect 132776 79416 132828 79422
rect 132776 79358 132828 79364
rect 132684 76628 132736 76634
rect 132684 76570 132736 76576
rect 132592 76492 132644 76498
rect 132592 76434 132644 76440
rect 132592 71732 132644 71738
rect 132592 71674 132644 71680
rect 132604 6914 132632 71674
rect 132696 10334 132724 76570
rect 132788 11830 132816 79358
rect 132880 24274 132908 79630
rect 132960 79620 133012 79626
rect 132960 79562 133012 79568
rect 132868 24268 132920 24274
rect 132868 24210 132920 24216
rect 132972 16574 133000 79562
rect 133064 77926 133092 79716
rect 133052 77920 133104 77926
rect 133052 77862 133104 77868
rect 133052 76900 133104 76906
rect 133052 76842 133104 76848
rect 133064 75818 133092 76842
rect 133052 75812 133104 75818
rect 133052 75754 133104 75760
rect 133156 72622 133184 79784
rect 133294 79744 133322 80036
rect 133248 79716 133322 79744
rect 133386 79744 133414 80036
rect 133478 79937 133506 80036
rect 133464 79928 133520 79937
rect 133464 79863 133520 79872
rect 133570 79778 133598 80036
rect 133662 79971 133690 80036
rect 133648 79962 133704 79971
rect 133648 79897 133704 79906
rect 133754 79898 133782 80036
rect 133742 79892 133794 79898
rect 133742 79834 133794 79840
rect 133570 79750 133736 79778
rect 133386 79716 133460 79744
rect 133248 76634 133276 79716
rect 133328 79552 133380 79558
rect 133328 79494 133380 79500
rect 133340 76838 133368 79494
rect 133328 76832 133380 76838
rect 133328 76774 133380 76780
rect 133432 76634 133460 79716
rect 133602 79656 133658 79665
rect 133512 79620 133564 79626
rect 133602 79591 133658 79600
rect 133512 79562 133564 79568
rect 133524 79286 133552 79562
rect 133512 79280 133564 79286
rect 133512 79222 133564 79228
rect 133236 76628 133288 76634
rect 133236 76570 133288 76576
rect 133420 76628 133472 76634
rect 133420 76570 133472 76576
rect 133144 72616 133196 72622
rect 133144 72558 133196 72564
rect 133616 70394 133644 79591
rect 133708 77722 133736 79750
rect 133846 79744 133874 80036
rect 133938 79966 133966 80036
rect 133926 79960 133978 79966
rect 134030 79937 134058 80036
rect 133926 79902 133978 79908
rect 134016 79928 134072 79937
rect 134016 79863 134072 79872
rect 133972 79824 134024 79830
rect 133972 79766 134024 79772
rect 133846 79716 133920 79744
rect 133788 79620 133840 79626
rect 133788 79562 133840 79568
rect 133696 77716 133748 77722
rect 133696 77658 133748 77664
rect 133800 76770 133828 79562
rect 133892 79422 133920 79716
rect 133880 79416 133932 79422
rect 133880 79358 133932 79364
rect 133880 79280 133932 79286
rect 133880 79222 133932 79228
rect 133892 79082 133920 79222
rect 133880 79076 133932 79082
rect 133880 79018 133932 79024
rect 133788 76764 133840 76770
rect 133788 76706 133840 76712
rect 133696 76628 133748 76634
rect 133696 76570 133748 76576
rect 133708 71398 133736 76570
rect 133984 73154 134012 79766
rect 134122 79744 134150 80036
rect 134214 79898 134242 80036
rect 134202 79892 134254 79898
rect 134202 79834 134254 79840
rect 134306 79744 134334 80036
rect 134076 79716 134150 79744
rect 134260 79716 134334 79744
rect 134076 76673 134104 79716
rect 134260 76809 134288 79716
rect 134398 79676 134426 80036
rect 134490 79744 134518 80036
rect 134582 79812 134610 80036
rect 134674 79966 134702 80036
rect 134766 79971 134794 80036
rect 134662 79960 134714 79966
rect 134662 79902 134714 79908
rect 134752 79962 134808 79971
rect 134858 79966 134886 80036
rect 134752 79897 134808 79906
rect 134846 79960 134898 79966
rect 134846 79902 134898 79908
rect 134708 79824 134760 79830
rect 134582 79784 134656 79812
rect 134490 79716 134564 79744
rect 134398 79648 134472 79676
rect 134246 76800 134302 76809
rect 134246 76735 134302 76744
rect 134062 76664 134118 76673
rect 134062 76599 134118 76608
rect 134064 75880 134116 75886
rect 134064 75822 134116 75828
rect 133892 73126 134012 73154
rect 133696 71392 133748 71398
rect 133696 71334 133748 71340
rect 133064 70366 133644 70394
rect 133064 69902 133092 70366
rect 133052 69896 133104 69902
rect 133052 69838 133104 69844
rect 132972 16546 133092 16574
rect 132776 11824 132828 11830
rect 132776 11766 132828 11772
rect 132684 10328 132736 10334
rect 132684 10270 132736 10276
rect 132604 6886 133000 6914
rect 132408 6112 132460 6118
rect 132408 6054 132460 6060
rect 132972 480 133000 6886
rect 133064 6594 133092 16546
rect 133052 6588 133104 6594
rect 133052 6530 133104 6536
rect 131734 354 131846 480
rect 131316 326 131846 354
rect 131734 -960 131846 326
rect 132930 -960 133042 480
rect 133892 354 133920 73126
rect 134076 10402 134104 75822
rect 134340 75336 134392 75342
rect 134340 75278 134392 75284
rect 134156 75200 134208 75206
rect 134156 75142 134208 75148
rect 134168 20058 134196 75142
rect 134352 71774 134380 75278
rect 134260 71746 134380 71774
rect 134260 68338 134288 71746
rect 134248 68332 134300 68338
rect 134248 68274 134300 68280
rect 134156 20052 134208 20058
rect 134156 19994 134208 20000
rect 134064 10396 134116 10402
rect 134064 10338 134116 10344
rect 134444 5166 134472 79648
rect 134536 72690 134564 79716
rect 134628 75342 134656 79784
rect 134950 79812 134978 80036
rect 134708 79766 134760 79772
rect 134798 79792 134854 79801
rect 134720 75886 134748 79766
rect 134798 79727 134854 79736
rect 134904 79784 134978 79812
rect 135042 79812 135070 80036
rect 135134 79966 135162 80036
rect 135122 79960 135174 79966
rect 135122 79902 135174 79908
rect 135226 79812 135254 80036
rect 135318 79898 135346 80036
rect 135410 79966 135438 80036
rect 135502 79971 135530 80036
rect 135398 79960 135450 79966
rect 135398 79902 135450 79908
rect 135488 79962 135544 79971
rect 135594 79966 135622 80036
rect 135686 79971 135714 80036
rect 135306 79892 135358 79898
rect 135488 79897 135544 79906
rect 135582 79960 135634 79966
rect 135582 79902 135634 79908
rect 135672 79962 135728 79971
rect 135672 79897 135728 79906
rect 135778 79898 135806 80036
rect 135306 79834 135358 79840
rect 135766 79892 135818 79898
rect 135766 79834 135818 79840
rect 135042 79784 135116 79812
rect 134812 79490 134840 79727
rect 134800 79484 134852 79490
rect 134800 79426 134852 79432
rect 134904 78470 134932 79784
rect 134982 79656 135038 79665
rect 134982 79591 135038 79600
rect 134892 78464 134944 78470
rect 134892 78406 134944 78412
rect 134708 75880 134760 75886
rect 134708 75822 134760 75828
rect 134616 75336 134668 75342
rect 134616 75278 134668 75284
rect 134996 74050 135024 79591
rect 134984 74044 135036 74050
rect 134984 73986 135036 73992
rect 135088 73154 135116 79784
rect 135180 79784 135254 79812
rect 135626 79792 135682 79801
rect 135180 75206 135208 79784
rect 135870 79778 135898 80036
rect 135962 79966 135990 80036
rect 135950 79960 136002 79966
rect 135950 79902 136002 79908
rect 136054 79898 136082 80036
rect 136042 79892 136094 79898
rect 136042 79834 136094 79840
rect 135720 79756 135772 79762
rect 135682 79736 135720 79744
rect 135626 79727 135720 79736
rect 135640 79716 135720 79727
rect 135870 79750 135944 79778
rect 135720 79698 135772 79704
rect 135352 79688 135404 79694
rect 135352 79630 135404 79636
rect 135718 79656 135774 79665
rect 135260 79552 135312 79558
rect 135260 79494 135312 79500
rect 135272 78402 135300 79494
rect 135364 78826 135392 79630
rect 135718 79591 135774 79600
rect 135536 79552 135588 79558
rect 135536 79494 135588 79500
rect 135364 78798 135484 78826
rect 135352 78668 135404 78674
rect 135352 78610 135404 78616
rect 135260 78396 135312 78402
rect 135260 78338 135312 78344
rect 135168 75200 135220 75206
rect 135168 75142 135220 75148
rect 134996 73126 135116 73154
rect 134524 72684 134576 72690
rect 134524 72626 134576 72632
rect 134996 71774 135024 73126
rect 134904 71746 135024 71774
rect 134904 71466 134932 71746
rect 135364 71738 135392 78610
rect 135456 77450 135484 78798
rect 135444 77444 135496 77450
rect 135444 77386 135496 77392
rect 135548 76906 135576 79494
rect 135536 76900 135588 76906
rect 135536 76842 135588 76848
rect 135628 76288 135680 76294
rect 135628 76230 135680 76236
rect 135536 75540 135588 75546
rect 135536 75482 135588 75488
rect 135444 75064 135496 75070
rect 135444 75006 135496 75012
rect 135352 71732 135404 71738
rect 135352 71674 135404 71680
rect 134892 71460 134944 71466
rect 134892 71402 134944 71408
rect 134432 5160 134484 5166
rect 134432 5102 134484 5108
rect 135456 3602 135484 75006
rect 135548 3670 135576 75482
rect 135640 4146 135668 76230
rect 135732 23934 135760 79591
rect 135916 78826 135944 79750
rect 136146 79744 136174 80036
rect 136100 79716 136174 79744
rect 135996 79416 136048 79422
rect 135996 79358 136048 79364
rect 135824 78798 135944 78826
rect 135824 78674 135852 78798
rect 135902 78704 135958 78713
rect 135812 78668 135864 78674
rect 135902 78639 135958 78648
rect 135812 78610 135864 78616
rect 135812 76628 135864 76634
rect 135812 76570 135864 76576
rect 135824 25022 135852 76570
rect 135916 76090 135944 78639
rect 135904 76084 135956 76090
rect 135904 76026 135956 76032
rect 136008 71774 136036 79358
rect 135916 71746 136036 71774
rect 135812 25016 135864 25022
rect 135812 24958 135864 24964
rect 135720 23928 135772 23934
rect 135720 23870 135772 23876
rect 135916 6914 135944 71746
rect 136100 70394 136128 79716
rect 136238 79676 136266 80036
rect 136330 79744 136358 80036
rect 136422 79937 136450 80036
rect 136408 79928 136464 79937
rect 136408 79863 136464 79872
rect 136514 79744 136542 80036
rect 136330 79716 136404 79744
rect 136192 79648 136266 79676
rect 136192 75070 136220 79648
rect 136376 77294 136404 79716
rect 136284 77266 136404 77294
rect 136468 79716 136542 79744
rect 136606 79744 136634 80036
rect 136698 79898 136726 80036
rect 136790 79937 136818 80036
rect 136776 79928 136832 79937
rect 136686 79892 136738 79898
rect 136882 79898 136910 80036
rect 136776 79863 136832 79872
rect 136870 79892 136922 79898
rect 136686 79834 136738 79840
rect 136870 79834 136922 79840
rect 136974 79801 137002 80036
rect 136730 79792 136786 79801
rect 136606 79716 136680 79744
rect 136730 79727 136786 79736
rect 136960 79792 137016 79801
rect 136960 79727 137016 79736
rect 137066 79744 137094 80036
rect 137158 79812 137186 80036
rect 137250 79966 137278 80036
rect 137238 79960 137290 79966
rect 137238 79902 137290 79908
rect 137158 79784 137232 79812
rect 136284 75546 136312 77266
rect 136468 76634 136496 79716
rect 136456 76628 136508 76634
rect 136456 76570 136508 76576
rect 136652 76294 136680 79716
rect 136640 76288 136692 76294
rect 136640 76230 136692 76236
rect 136640 76152 136692 76158
rect 136640 76094 136692 76100
rect 136272 75540 136324 75546
rect 136272 75482 136324 75488
rect 136180 75064 136232 75070
rect 136180 75006 136232 75012
rect 136008 70366 136128 70394
rect 136008 16574 136036 70366
rect 136008 16546 136496 16574
rect 135732 6886 135944 6914
rect 135628 4140 135680 4146
rect 135628 4082 135680 4088
rect 135536 3664 135588 3670
rect 135536 3606 135588 3612
rect 135444 3596 135496 3602
rect 135444 3538 135496 3544
rect 135732 3482 135760 6886
rect 135272 3454 135760 3482
rect 135272 480 135300 3454
rect 136468 480 136496 16546
rect 136652 4894 136680 76094
rect 136744 74662 136772 79727
rect 137066 79716 137140 79744
rect 136824 79688 136876 79694
rect 136824 79630 136876 79636
rect 136914 79656 136970 79665
rect 136732 74656 136784 74662
rect 136732 74598 136784 74604
rect 136732 73772 136784 73778
rect 136732 73714 136784 73720
rect 136744 5234 136772 73714
rect 136836 11830 136864 79630
rect 136914 79591 136970 79600
rect 137008 79620 137060 79626
rect 136928 76945 136956 79591
rect 137008 79562 137060 79568
rect 136914 76936 136970 76945
rect 136914 76871 136970 76880
rect 136916 76764 136968 76770
rect 136916 76706 136968 76712
rect 136928 22846 136956 76706
rect 137020 76616 137048 79562
rect 137112 76770 137140 79716
rect 137100 76764 137152 76770
rect 137100 76706 137152 76712
rect 137020 76588 137140 76616
rect 137008 74656 137060 74662
rect 137008 74598 137060 74604
rect 137020 57934 137048 74598
rect 137112 60722 137140 76588
rect 137204 62830 137232 79784
rect 137342 79744 137370 80036
rect 137296 79716 137370 79744
rect 137296 69018 137324 79716
rect 137434 79676 137462 80036
rect 137526 79744 137554 80036
rect 137618 79966 137646 80036
rect 137606 79960 137658 79966
rect 137606 79902 137658 79908
rect 137710 79812 137738 80036
rect 137664 79784 137738 79812
rect 137526 79716 137600 79744
rect 137388 79648 137462 79676
rect 137388 75954 137416 79648
rect 137468 79552 137520 79558
rect 137468 79494 137520 79500
rect 137376 75948 137428 75954
rect 137376 75890 137428 75896
rect 137480 73914 137508 79494
rect 137468 73908 137520 73914
rect 137468 73850 137520 73856
rect 137572 73778 137600 79716
rect 137664 76537 137692 79784
rect 137802 79744 137830 80036
rect 137894 79801 137922 80036
rect 137986 79937 138014 80036
rect 137972 79928 138028 79937
rect 137972 79863 138028 79872
rect 138078 79812 138106 80036
rect 137756 79716 137830 79744
rect 137880 79792 137936 79801
rect 137880 79727 137936 79736
rect 138032 79784 138106 79812
rect 137650 76528 137706 76537
rect 137650 76463 137706 76472
rect 137756 76158 137784 79716
rect 137836 79620 137888 79626
rect 137836 79562 137888 79568
rect 137848 77994 137876 79562
rect 138032 78690 138060 79784
rect 138170 79744 138198 80036
rect 137940 78662 138060 78690
rect 138124 79716 138198 79744
rect 138262 79744 138290 80036
rect 138354 79898 138382 80036
rect 138342 79892 138394 79898
rect 138342 79834 138394 79840
rect 138446 79744 138474 80036
rect 138538 79966 138566 80036
rect 138526 79960 138578 79966
rect 138630 79937 138658 80036
rect 138722 79966 138750 80036
rect 138710 79960 138762 79966
rect 138526 79902 138578 79908
rect 138616 79928 138672 79937
rect 138710 79902 138762 79908
rect 138616 79863 138672 79872
rect 138814 79830 138842 80036
rect 138906 79966 138934 80036
rect 138998 79971 139026 80036
rect 138894 79960 138946 79966
rect 138894 79902 138946 79908
rect 138984 79962 139040 79971
rect 139090 79966 139118 80036
rect 138984 79897 139040 79906
rect 139078 79960 139130 79966
rect 139078 79902 139130 79908
rect 139182 79898 139210 80036
rect 139170 79892 139222 79898
rect 139170 79834 139222 79840
rect 138572 79824 138624 79830
rect 138572 79766 138624 79772
rect 138664 79824 138716 79830
rect 138664 79766 138716 79772
rect 138802 79824 138854 79830
rect 138802 79766 138854 79772
rect 138262 79716 138336 79744
rect 137836 77988 137888 77994
rect 137836 77930 137888 77936
rect 137940 76673 137968 78662
rect 138020 77988 138072 77994
rect 138020 77930 138072 77936
rect 137926 76664 137982 76673
rect 137926 76599 137982 76608
rect 137928 76492 137980 76498
rect 137928 76434 137980 76440
rect 137744 76152 137796 76158
rect 137744 76094 137796 76100
rect 137560 73772 137612 73778
rect 137560 73714 137612 73720
rect 137940 73154 137968 76434
rect 138032 73302 138060 77930
rect 138020 73296 138072 73302
rect 138020 73238 138072 73244
rect 137940 73126 138060 73154
rect 137284 69012 137336 69018
rect 137284 68954 137336 68960
rect 137192 62824 137244 62830
rect 137192 62766 137244 62772
rect 137100 60716 137152 60722
rect 137100 60658 137152 60664
rect 137008 57928 137060 57934
rect 137008 57870 137060 57876
rect 136916 22840 136968 22846
rect 136916 22782 136968 22788
rect 136824 11824 136876 11830
rect 136824 11766 136876 11772
rect 136732 5228 136784 5234
rect 136732 5170 136784 5176
rect 138032 5166 138060 73126
rect 138020 5160 138072 5166
rect 138020 5102 138072 5108
rect 136640 4888 136692 4894
rect 136640 4830 136692 4836
rect 138124 4826 138152 79716
rect 138204 79620 138256 79626
rect 138204 79562 138256 79568
rect 138216 11762 138244 79562
rect 138308 76634 138336 79716
rect 138400 79716 138474 79744
rect 138296 76628 138348 76634
rect 138296 76570 138348 76576
rect 138294 76528 138350 76537
rect 138294 76463 138350 76472
rect 138308 44946 138336 76463
rect 138400 49026 138428 79716
rect 138480 74588 138532 74594
rect 138480 74530 138532 74536
rect 138492 51746 138520 74530
rect 138584 66230 138612 79766
rect 138676 76498 138704 79766
rect 139032 79756 139084 79762
rect 139274 79744 139302 80036
rect 139366 79778 139394 80036
rect 139458 79966 139486 80036
rect 139446 79960 139498 79966
rect 139446 79902 139498 79908
rect 139550 79812 139578 80036
rect 139642 79937 139670 80036
rect 139628 79928 139684 79937
rect 139628 79863 139684 79872
rect 139550 79784 139624 79812
rect 139596 79778 139624 79784
rect 139366 79750 139440 79778
rect 139596 79750 139670 79778
rect 139032 79698 139084 79704
rect 139228 79716 139302 79744
rect 138756 79688 138808 79694
rect 138756 79630 138808 79636
rect 138848 79688 138900 79694
rect 138848 79630 138900 79636
rect 138664 76492 138716 76498
rect 138664 76434 138716 76440
rect 138768 74594 138796 79630
rect 138860 76770 138888 79630
rect 138940 79620 138992 79626
rect 138940 79562 138992 79568
rect 138848 76764 138900 76770
rect 138848 76706 138900 76712
rect 138952 76673 138980 79562
rect 138938 76664 138994 76673
rect 138848 76628 138900 76634
rect 138938 76599 138994 76608
rect 138848 76570 138900 76576
rect 138756 74588 138808 74594
rect 138756 74530 138808 74536
rect 138860 70394 138888 76570
rect 139044 75857 139072 79698
rect 139228 78690 139256 79716
rect 139412 79642 139440 79750
rect 139136 78662 139256 78690
rect 139320 79614 139440 79642
rect 139492 79688 139544 79694
rect 139642 79676 139670 79750
rect 139734 79744 139762 80036
rect 139826 79812 139854 80036
rect 139918 79966 139946 80036
rect 139906 79960 139958 79966
rect 139906 79902 139958 79908
rect 139826 79784 139900 79812
rect 139734 79716 139808 79744
rect 139492 79630 139544 79636
rect 139596 79648 139670 79676
rect 139136 76809 139164 78662
rect 139320 77294 139348 79614
rect 139504 77994 139532 79630
rect 139492 77988 139544 77994
rect 139492 77930 139544 77936
rect 139228 77266 139348 77294
rect 139122 76800 139178 76809
rect 139122 76735 139178 76744
rect 139030 75848 139086 75857
rect 139030 75783 139086 75792
rect 139228 75721 139256 77266
rect 139308 76764 139360 76770
rect 139308 76706 139360 76712
rect 139492 76764 139544 76770
rect 139492 76706 139544 76712
rect 139214 75712 139270 75721
rect 139214 75647 139270 75656
rect 139216 73908 139268 73914
rect 139216 73850 139268 73856
rect 139228 70394 139256 73850
rect 139320 71058 139348 76706
rect 139504 76378 139532 76706
rect 139596 76566 139624 79648
rect 139676 79552 139728 79558
rect 139676 79494 139728 79500
rect 139584 76560 139636 76566
rect 139584 76502 139636 76508
rect 139504 76350 139624 76378
rect 139492 74656 139544 74662
rect 139492 74598 139544 74604
rect 139308 71052 139360 71058
rect 139308 70994 139360 71000
rect 138676 70366 138888 70394
rect 138952 70366 139256 70394
rect 138676 68950 138704 70366
rect 138756 69012 138808 69018
rect 138756 68954 138808 68960
rect 138664 68944 138716 68950
rect 138664 68886 138716 68892
rect 138572 66224 138624 66230
rect 138572 66166 138624 66172
rect 138480 51740 138532 51746
rect 138480 51682 138532 51688
rect 138388 49020 138440 49026
rect 138388 48962 138440 48968
rect 138296 44940 138348 44946
rect 138296 44882 138348 44888
rect 138204 11756 138256 11762
rect 138204 11698 138256 11704
rect 138112 4820 138164 4826
rect 138112 4762 138164 4768
rect 136548 4140 136600 4146
rect 136548 4082 136600 4088
rect 136560 3330 136588 4082
rect 138768 3602 138796 68954
rect 138952 64874 138980 70366
rect 138860 64846 138980 64874
rect 138860 22098 138888 64846
rect 138848 22092 138900 22098
rect 138848 22034 138900 22040
rect 139504 4078 139532 74598
rect 139596 27130 139624 76350
rect 139688 43586 139716 79494
rect 139780 76498 139808 79716
rect 139768 76492 139820 76498
rect 139768 76434 139820 76440
rect 139768 76356 139820 76362
rect 139768 76298 139820 76304
rect 139780 46374 139808 76298
rect 139872 49298 139900 79784
rect 140010 79744 140038 80036
rect 140102 79898 140130 80036
rect 140090 79892 140142 79898
rect 140090 79834 140142 79840
rect 140194 79778 140222 80036
rect 140286 79898 140314 80036
rect 140378 79966 140406 80036
rect 140366 79960 140418 79966
rect 140366 79902 140418 79908
rect 140274 79892 140326 79898
rect 140274 79834 140326 79840
rect 140470 79801 140498 80036
rect 140562 79937 140590 80036
rect 140548 79928 140604 79937
rect 140548 79863 140604 79872
rect 140148 79750 140222 79778
rect 140456 79792 140512 79801
rect 140010 79716 140084 79744
rect 139950 79656 140006 79665
rect 139950 79591 140006 79600
rect 140056 79608 140084 79716
rect 140148 79676 140176 79750
rect 140654 79744 140682 80036
rect 140456 79727 140512 79736
rect 140608 79716 140682 79744
rect 140148 79648 140268 79676
rect 139964 76650 139992 79591
rect 140056 79580 140176 79608
rect 140044 79484 140096 79490
rect 140044 79426 140096 79432
rect 140056 76770 140084 79426
rect 140044 76764 140096 76770
rect 140044 76706 140096 76712
rect 139964 76622 140084 76650
rect 139952 76560 140004 76566
rect 139952 76502 140004 76508
rect 139964 57594 139992 76502
rect 140056 60382 140084 76622
rect 140148 70394 140176 79580
rect 140240 76362 140268 79648
rect 140320 79552 140372 79558
rect 140320 79494 140372 79500
rect 140504 79552 140556 79558
rect 140504 79494 140556 79500
rect 140228 76356 140280 76362
rect 140228 76298 140280 76304
rect 140332 74662 140360 79494
rect 140516 76702 140544 79494
rect 140504 76696 140556 76702
rect 140608 76673 140636 79716
rect 140746 79676 140774 80036
rect 140838 79801 140866 80036
rect 140930 79898 140958 80036
rect 141022 79898 141050 80036
rect 141114 79898 141142 80036
rect 140918 79892 140970 79898
rect 140918 79834 140970 79840
rect 141010 79892 141062 79898
rect 141010 79834 141062 79840
rect 141102 79892 141154 79898
rect 141102 79834 141154 79840
rect 140824 79792 140880 79801
rect 141206 79744 141234 80036
rect 141298 79966 141326 80036
rect 141286 79960 141338 79966
rect 141286 79902 141338 79908
rect 140824 79727 140880 79736
rect 141068 79716 141234 79744
rect 141390 79744 141418 80036
rect 141482 79898 141510 80036
rect 141574 79966 141602 80036
rect 141562 79960 141614 79966
rect 141562 79902 141614 79908
rect 141470 79892 141522 79898
rect 141470 79834 141522 79840
rect 141516 79756 141568 79762
rect 141390 79716 141464 79744
rect 140700 79648 140774 79676
rect 140964 79688 141016 79694
rect 140504 76638 140556 76644
rect 140594 76664 140650 76673
rect 140594 76599 140650 76608
rect 140320 74656 140372 74662
rect 140320 74598 140372 74604
rect 140700 74361 140728 79648
rect 140884 79636 140964 79642
rect 140884 79630 141016 79636
rect 140884 79614 141004 79630
rect 140780 76628 140832 76634
rect 140780 76570 140832 76576
rect 140686 74352 140742 74361
rect 140686 74287 140742 74296
rect 140148 70366 140360 70394
rect 140136 68944 140188 68950
rect 140136 68886 140188 68892
rect 140044 60376 140096 60382
rect 140044 60318 140096 60324
rect 140044 57928 140096 57934
rect 140044 57870 140096 57876
rect 139952 57588 140004 57594
rect 139952 57530 140004 57536
rect 139860 49292 139912 49298
rect 139860 49234 139912 49240
rect 139768 46368 139820 46374
rect 139768 46310 139820 46316
rect 139676 43580 139728 43586
rect 139676 43522 139728 43528
rect 139584 27124 139636 27130
rect 139584 27066 139636 27072
rect 139584 23928 139636 23934
rect 139584 23870 139636 23876
rect 139492 4072 139544 4078
rect 139492 4014 139544 4020
rect 138848 3664 138900 3670
rect 138848 3606 138900 3612
rect 137652 3596 137704 3602
rect 137652 3538 137704 3544
rect 138756 3596 138808 3602
rect 138756 3538 138808 3544
rect 136548 3324 136600 3330
rect 136548 3266 136600 3272
rect 137664 480 137692 3538
rect 138860 480 138888 3606
rect 134126 354 134238 480
rect 133892 326 134238 354
rect 134126 -960 134238 326
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 139596 354 139624 23870
rect 140056 3262 140084 57870
rect 140148 3534 140176 68886
rect 140228 66224 140280 66230
rect 140228 66166 140280 66172
rect 140136 3528 140188 3534
rect 140136 3470 140188 3476
rect 140240 3466 140268 66166
rect 140332 4146 140360 70366
rect 140792 5098 140820 76570
rect 140884 24410 140912 79614
rect 140964 79552 141016 79558
rect 140964 79494 141016 79500
rect 140976 25906 141004 79494
rect 141068 28558 141096 79716
rect 141238 79656 141294 79665
rect 141148 79620 141200 79626
rect 141238 79591 141294 79600
rect 141332 79620 141384 79626
rect 141148 79562 141200 79568
rect 141160 77926 141188 79562
rect 141252 78538 141280 79591
rect 141332 79562 141384 79568
rect 141240 78532 141292 78538
rect 141240 78474 141292 78480
rect 141148 77920 141200 77926
rect 141148 77862 141200 77868
rect 141344 76650 141372 79562
rect 141160 76622 141372 76650
rect 141160 45082 141188 76622
rect 141240 76560 141292 76566
rect 141240 76502 141292 76508
rect 141252 51882 141280 76502
rect 141332 73840 141384 73846
rect 141332 73782 141384 73788
rect 141344 64462 141372 73782
rect 141436 68610 141464 79716
rect 141666 79744 141694 80036
rect 141758 79898 141786 80036
rect 141746 79892 141798 79898
rect 141746 79834 141798 79840
rect 141850 79744 141878 80036
rect 141516 79698 141568 79704
rect 141620 79716 141694 79744
rect 141804 79716 141878 79744
rect 141528 76566 141556 79698
rect 141516 76560 141568 76566
rect 141516 76502 141568 76508
rect 141620 73846 141648 79716
rect 141700 79552 141752 79558
rect 141700 79494 141752 79500
rect 141712 76634 141740 79494
rect 141700 76628 141752 76634
rect 141700 76570 141752 76576
rect 141804 74186 141832 79716
rect 141942 79676 141970 80036
rect 142034 79778 142062 80036
rect 142126 79937 142154 80036
rect 142112 79928 142168 79937
rect 142218 79898 142246 80036
rect 142112 79863 142168 79872
rect 142206 79892 142258 79898
rect 142206 79834 142258 79840
rect 142034 79750 142200 79778
rect 141942 79648 142016 79676
rect 141884 79484 141936 79490
rect 141884 79426 141936 79432
rect 141896 77586 141924 79426
rect 141884 77580 141936 77586
rect 141884 77522 141936 77528
rect 141792 74180 141844 74186
rect 141792 74122 141844 74128
rect 141608 73840 141660 73846
rect 141608 73782 141660 73788
rect 141988 71774 142016 79648
rect 142172 79642 142200 79750
rect 142310 79744 142338 80036
rect 142402 79971 142430 80036
rect 142388 79962 142444 79971
rect 142494 79966 142522 80036
rect 142586 79966 142614 80036
rect 142388 79897 142444 79906
rect 142482 79960 142534 79966
rect 142482 79902 142534 79908
rect 142574 79960 142626 79966
rect 142574 79902 142626 79908
rect 142678 79778 142706 80036
rect 142770 79966 142798 80036
rect 142862 79966 142890 80036
rect 142954 79966 142982 80036
rect 143046 79966 143074 80036
rect 142758 79960 142810 79966
rect 142758 79902 142810 79908
rect 142850 79960 142902 79966
rect 142850 79902 142902 79908
rect 142942 79960 142994 79966
rect 142942 79902 142994 79908
rect 143034 79960 143086 79966
rect 143138 79937 143166 80036
rect 143034 79902 143086 79908
rect 143124 79928 143180 79937
rect 143124 79863 143180 79872
rect 142894 79792 142950 79801
rect 142528 79756 142580 79762
rect 142310 79716 142430 79744
rect 142402 79676 142430 79716
rect 142678 79750 142752 79778
rect 142724 79744 142752 79750
rect 142724 79716 142844 79744
rect 143230 79778 143258 80036
rect 143322 79830 143350 80036
rect 143414 79830 143442 80036
rect 143506 79971 143534 80036
rect 143492 79962 143548 79971
rect 143492 79897 143548 79906
rect 143598 79830 143626 80036
rect 143690 79830 143718 80036
rect 142894 79727 142950 79736
rect 143184 79750 143258 79778
rect 143310 79824 143362 79830
rect 143310 79766 143362 79772
rect 143402 79824 143454 79830
rect 143402 79766 143454 79772
rect 143586 79824 143638 79830
rect 143586 79766 143638 79772
rect 143678 79824 143730 79830
rect 143678 79766 143730 79772
rect 143782 79778 143810 80036
rect 143874 79898 143902 80036
rect 143862 79892 143914 79898
rect 143862 79834 143914 79840
rect 143966 79830 143994 80036
rect 144058 79971 144086 80036
rect 144044 79962 144100 79971
rect 144150 79966 144178 80036
rect 144242 79966 144270 80036
rect 144334 79966 144362 80036
rect 144426 79966 144454 80036
rect 144518 79971 144546 80036
rect 144044 79897 144100 79906
rect 144138 79960 144190 79966
rect 144138 79902 144190 79908
rect 144230 79960 144282 79966
rect 144230 79902 144282 79908
rect 144322 79960 144374 79966
rect 144322 79902 144374 79908
rect 144414 79960 144466 79966
rect 144414 79902 144466 79908
rect 144504 79962 144560 79971
rect 144610 79966 144638 80036
rect 144702 79966 144730 80036
rect 144504 79897 144560 79906
rect 144598 79960 144650 79966
rect 144598 79902 144650 79908
rect 144690 79960 144742 79966
rect 144690 79902 144742 79908
rect 143954 79824 144006 79830
rect 143782 79750 143902 79778
rect 144794 79801 144822 80036
rect 143954 79766 144006 79772
rect 144780 79792 144836 79801
rect 142528 79698 142580 79704
rect 142402 79648 142476 79676
rect 142080 79614 142200 79642
rect 142252 79620 142304 79626
rect 142080 77217 142108 79614
rect 142252 79562 142304 79568
rect 142160 79484 142212 79490
rect 142160 79426 142212 79432
rect 142066 77208 142122 77217
rect 142066 77143 142122 77152
rect 141896 71746 142016 71774
rect 141896 70394 141924 71746
rect 141528 70366 141924 70394
rect 141528 70038 141556 70366
rect 141516 70032 141568 70038
rect 141516 69974 141568 69980
rect 141424 68604 141476 68610
rect 141424 68546 141476 68552
rect 141332 64456 141384 64462
rect 141332 64398 141384 64404
rect 141240 51876 141292 51882
rect 141240 51818 141292 51824
rect 141148 45076 141200 45082
rect 141148 45018 141200 45024
rect 141056 28552 141108 28558
rect 141056 28494 141108 28500
rect 140964 25900 141016 25906
rect 140964 25842 141016 25848
rect 140964 25016 141016 25022
rect 140964 24958 141016 24964
rect 140872 24404 140924 24410
rect 140872 24346 140924 24352
rect 140976 16574 141004 24958
rect 140976 16546 141280 16574
rect 140780 5092 140832 5098
rect 140780 5034 140832 5040
rect 140320 4140 140372 4146
rect 140320 4082 140372 4088
rect 140228 3460 140280 3466
rect 140228 3402 140280 3408
rect 140044 3256 140096 3262
rect 140044 3198 140096 3204
rect 141252 480 141280 16546
rect 142172 7954 142200 79426
rect 142264 78334 142292 79562
rect 142344 79552 142396 79558
rect 142344 79494 142396 79500
rect 142252 78328 142304 78334
rect 142252 78270 142304 78276
rect 142252 76560 142304 76566
rect 142252 76502 142304 76508
rect 142264 32434 142292 76502
rect 142356 42226 142384 79494
rect 142448 47734 142476 79648
rect 142540 75546 142568 79698
rect 142712 79620 142764 79626
rect 142712 79562 142764 79568
rect 142724 76650 142752 79562
rect 142632 76622 142752 76650
rect 142528 75540 142580 75546
rect 142528 75482 142580 75488
rect 142528 75404 142580 75410
rect 142528 75346 142580 75352
rect 142540 61674 142568 75346
rect 142632 64394 142660 76622
rect 142816 76566 142844 79716
rect 142908 76702 142936 79727
rect 143080 79620 143132 79626
rect 143080 79562 143132 79568
rect 142896 76696 142948 76702
rect 142896 76638 142948 76644
rect 142804 76560 142856 76566
rect 142804 76502 142856 76508
rect 142712 75540 142764 75546
rect 142712 75482 142764 75488
rect 142724 65686 142752 75482
rect 143092 75410 143120 79562
rect 143184 76673 143212 79750
rect 143264 79688 143316 79694
rect 143264 79630 143316 79636
rect 143540 79688 143592 79694
rect 143540 79630 143592 79636
rect 143874 79642 143902 79750
rect 144780 79727 144836 79736
rect 144000 79688 144052 79694
rect 143170 76664 143226 76673
rect 143170 76599 143226 76608
rect 143276 76537 143304 79630
rect 143448 79620 143500 79626
rect 143448 79562 143500 79568
rect 143356 79552 143408 79558
rect 143356 79494 143408 79500
rect 143262 76528 143318 76537
rect 143262 76463 143318 76472
rect 143080 75404 143132 75410
rect 143080 75346 143132 75352
rect 143368 74050 143396 79494
rect 143460 76673 143488 79562
rect 143552 77790 143580 79630
rect 143874 79614 143948 79642
rect 144000 79630 144052 79636
rect 144184 79688 144236 79694
rect 144886 79676 144914 80036
rect 144184 79630 144236 79636
rect 144458 79656 144514 79665
rect 143724 79552 143776 79558
rect 143724 79494 143776 79500
rect 143540 77784 143592 77790
rect 143540 77726 143592 77732
rect 143632 77172 143684 77178
rect 143632 77114 143684 77120
rect 143446 76664 143502 76673
rect 143446 76599 143502 76608
rect 143356 74044 143408 74050
rect 143356 73986 143408 73992
rect 142988 73296 143040 73302
rect 142988 73238 143040 73244
rect 142712 65680 142764 65686
rect 142712 65622 142764 65628
rect 142620 64388 142672 64394
rect 142620 64330 142672 64336
rect 142528 61668 142580 61674
rect 142528 61610 142580 61616
rect 142804 60716 142856 60722
rect 142804 60658 142856 60664
rect 142436 47728 142488 47734
rect 142436 47670 142488 47676
rect 142344 42220 142396 42226
rect 142344 42162 142396 42168
rect 142252 32428 142304 32434
rect 142252 32370 142304 32376
rect 142160 7948 142212 7954
rect 142160 7890 142212 7896
rect 142816 3330 142844 60658
rect 143000 3670 143028 73238
rect 143644 18902 143672 77114
rect 143736 20058 143764 79494
rect 143816 79484 143868 79490
rect 143816 79426 143868 79432
rect 143828 76770 143856 79426
rect 143920 77178 143948 79614
rect 143908 77172 143960 77178
rect 143908 77114 143960 77120
rect 144012 76906 144040 79630
rect 144092 79620 144144 79626
rect 144092 79562 144144 79568
rect 144000 76900 144052 76906
rect 144000 76842 144052 76848
rect 144104 76838 144132 79562
rect 144196 77058 144224 79630
rect 144840 79648 144914 79676
rect 144978 79676 145006 80036
rect 145070 79744 145098 80036
rect 145162 79898 145190 80036
rect 145254 79898 145282 80036
rect 145150 79892 145202 79898
rect 145150 79834 145202 79840
rect 145242 79892 145294 79898
rect 145242 79834 145294 79840
rect 145346 79778 145374 80036
rect 145208 79750 145374 79778
rect 145070 79716 145144 79744
rect 144978 79648 145052 79676
rect 144458 79591 144514 79600
rect 144736 79620 144788 79626
rect 144368 79484 144420 79490
rect 144368 79426 144420 79432
rect 144196 77030 144316 77058
rect 144184 76900 144236 76906
rect 144184 76842 144236 76848
rect 143908 76832 143960 76838
rect 143908 76774 143960 76780
rect 144092 76832 144144 76838
rect 144092 76774 144144 76780
rect 143816 76764 143868 76770
rect 143816 76706 143868 76712
rect 143816 76628 143868 76634
rect 143816 76570 143868 76576
rect 143828 28490 143856 76570
rect 143920 46306 143948 76774
rect 144000 76764 144052 76770
rect 144000 76706 144052 76712
rect 144012 50658 144040 76706
rect 144092 74588 144144 74594
rect 144092 74530 144144 74536
rect 144104 62966 144132 74530
rect 144196 65618 144224 76842
rect 144288 68542 144316 77030
rect 144380 74594 144408 79426
rect 144472 76634 144500 79591
rect 144736 79562 144788 79568
rect 144748 76809 144776 79562
rect 144734 76800 144790 76809
rect 144734 76735 144790 76744
rect 144550 76664 144606 76673
rect 144460 76628 144512 76634
rect 144550 76599 144606 76608
rect 144460 76570 144512 76576
rect 144460 75948 144512 75954
rect 144460 75890 144512 75896
rect 144368 74588 144420 74594
rect 144368 74530 144420 74536
rect 144276 68536 144328 68542
rect 144276 68478 144328 68484
rect 144184 65612 144236 65618
rect 144184 65554 144236 65560
rect 144092 62960 144144 62966
rect 144092 62902 144144 62908
rect 144184 62824 144236 62830
rect 144184 62766 144236 62772
rect 144000 50652 144052 50658
rect 144000 50594 144052 50600
rect 143908 46300 143960 46306
rect 143908 46242 143960 46248
rect 143816 28484 143868 28490
rect 143816 28426 143868 28432
rect 143816 22092 143868 22098
rect 143816 22034 143868 22040
rect 143724 20052 143776 20058
rect 143724 19994 143776 20000
rect 143632 18896 143684 18902
rect 143632 18838 143684 18844
rect 143828 6914 143856 22034
rect 143552 6886 143856 6914
rect 142988 3664 143040 3670
rect 142988 3606 143040 3612
rect 142436 3324 142488 3330
rect 142436 3266 142488 3272
rect 142804 3324 142856 3330
rect 142804 3266 142856 3272
rect 142448 480 142476 3266
rect 143552 480 143580 6886
rect 144196 3398 144224 62766
rect 144184 3392 144236 3398
rect 144184 3334 144236 3340
rect 144472 3194 144500 75890
rect 144564 16114 144592 76599
rect 144840 76537 144868 79648
rect 144920 79552 144972 79558
rect 144920 79494 144972 79500
rect 144932 78266 144960 79494
rect 144920 78260 144972 78266
rect 144920 78202 144972 78208
rect 145024 77654 145052 79648
rect 145012 77648 145064 77654
rect 145012 77590 145064 77596
rect 145012 76628 145064 76634
rect 145012 76570 145064 76576
rect 144826 76528 144882 76537
rect 144826 76463 144882 76472
rect 144920 76152 144972 76158
rect 144920 76094 144972 76100
rect 144932 20194 144960 76094
rect 144920 20188 144972 20194
rect 144920 20130 144972 20136
rect 145024 20126 145052 76570
rect 145116 29986 145144 79716
rect 145104 29980 145156 29986
rect 145104 29922 145156 29928
rect 145208 29918 145236 79750
rect 145288 79688 145340 79694
rect 145438 79676 145466 80036
rect 145288 79630 145340 79636
rect 145392 79648 145466 79676
rect 145530 79676 145558 80036
rect 145622 79778 145650 80036
rect 145714 79966 145742 80036
rect 145806 79966 145834 80036
rect 145702 79960 145754 79966
rect 145702 79902 145754 79908
rect 145794 79960 145846 79966
rect 145794 79902 145846 79908
rect 145748 79824 145800 79830
rect 145622 79750 145696 79778
rect 145748 79766 145800 79772
rect 145530 79648 145604 79676
rect 145300 78198 145328 79630
rect 145288 78192 145340 78198
rect 145288 78134 145340 78140
rect 145288 78056 145340 78062
rect 145288 77998 145340 78004
rect 145300 33998 145328 77998
rect 145392 76634 145420 79648
rect 145472 79212 145524 79218
rect 145472 79154 145524 79160
rect 145484 78946 145512 79154
rect 145472 78940 145524 78946
rect 145472 78882 145524 78888
rect 145380 76628 145432 76634
rect 145380 76570 145432 76576
rect 145380 76424 145432 76430
rect 145380 76366 145432 76372
rect 145392 38010 145420 76366
rect 145472 74316 145524 74322
rect 145472 74258 145524 74264
rect 145484 60314 145512 74258
rect 145576 67114 145604 79648
rect 145668 76430 145696 79750
rect 145656 76424 145708 76430
rect 145656 76366 145708 76372
rect 145760 74322 145788 79766
rect 145898 79540 145926 80036
rect 145990 79676 146018 80036
rect 146082 79801 146110 80036
rect 146174 79937 146202 80036
rect 146266 79966 146294 80036
rect 146358 79966 146386 80036
rect 146254 79960 146306 79966
rect 146160 79928 146216 79937
rect 146254 79902 146306 79908
rect 146346 79960 146398 79966
rect 146346 79902 146398 79908
rect 146450 79898 146478 80036
rect 146160 79863 146216 79872
rect 146438 79892 146490 79898
rect 146438 79834 146490 79840
rect 146068 79792 146124 79801
rect 146068 79727 146124 79736
rect 146300 79756 146352 79762
rect 146542 79744 146570 80036
rect 146634 79937 146662 80036
rect 146620 79928 146676 79937
rect 146620 79863 146676 79872
rect 146726 79801 146754 80036
rect 146818 79830 146846 80036
rect 146910 79937 146938 80036
rect 146896 79928 146952 79937
rect 147002 79898 147030 80036
rect 146896 79863 146952 79872
rect 146990 79892 147042 79898
rect 146990 79834 147042 79840
rect 146806 79824 146858 79830
rect 146712 79792 146768 79801
rect 146542 79716 146616 79744
rect 146806 79766 146858 79772
rect 146712 79727 146768 79736
rect 147094 79744 147122 80036
rect 147186 79966 147214 80036
rect 147174 79960 147226 79966
rect 147278 79937 147306 80036
rect 147370 79966 147398 80036
rect 147462 79966 147490 80036
rect 147554 79966 147582 80036
rect 147646 79966 147674 80036
rect 147358 79960 147410 79966
rect 147174 79902 147226 79908
rect 147264 79928 147320 79937
rect 147358 79902 147410 79908
rect 147450 79960 147502 79966
rect 147450 79902 147502 79908
rect 147542 79960 147594 79966
rect 147542 79902 147594 79908
rect 147634 79960 147686 79966
rect 147634 79902 147686 79908
rect 147264 79863 147320 79872
rect 147496 79756 147548 79762
rect 147094 79716 147168 79744
rect 146300 79698 146352 79704
rect 146116 79688 146168 79694
rect 145990 79648 146064 79676
rect 145898 79512 145972 79540
rect 145840 77988 145892 77994
rect 145840 77930 145892 77936
rect 145852 76430 145880 77930
rect 145944 77042 145972 79512
rect 145932 77036 145984 77042
rect 145932 76978 145984 76984
rect 145840 76424 145892 76430
rect 145840 76366 145892 76372
rect 146036 76158 146064 79648
rect 146116 79630 146168 79636
rect 146128 76974 146156 79630
rect 146116 76968 146168 76974
rect 146116 76910 146168 76916
rect 146208 76764 146260 76770
rect 146208 76706 146260 76712
rect 146024 76152 146076 76158
rect 146024 76094 146076 76100
rect 145748 74316 145800 74322
rect 145748 74258 145800 74264
rect 146220 73154 146248 76706
rect 146312 76673 146340 79698
rect 146392 79620 146444 79626
rect 146392 79562 146444 79568
rect 146298 76664 146354 76673
rect 146404 76634 146432 79562
rect 146588 76906 146616 79716
rect 146852 79688 146904 79694
rect 146772 79648 146852 79676
rect 146668 79620 146720 79626
rect 146668 79562 146720 79568
rect 146576 76900 146628 76906
rect 146576 76842 146628 76848
rect 146574 76800 146630 76809
rect 146680 76770 146708 79562
rect 146574 76735 146630 76744
rect 146668 76764 146720 76770
rect 146482 76664 146538 76673
rect 146298 76599 146354 76608
rect 146392 76628 146444 76634
rect 146482 76599 146538 76608
rect 146392 76570 146444 76576
rect 146390 76528 146446 76537
rect 146390 76463 146446 76472
rect 146298 76392 146354 76401
rect 146298 76327 146354 76336
rect 146312 74118 146340 76327
rect 146300 74112 146352 74118
rect 146300 74054 146352 74060
rect 146220 73126 146340 73154
rect 145564 67108 145616 67114
rect 145564 67050 145616 67056
rect 145472 60308 145524 60314
rect 145472 60250 145524 60256
rect 145380 38004 145432 38010
rect 145380 37946 145432 37952
rect 145288 33992 145340 33998
rect 145288 33934 145340 33940
rect 145196 29912 145248 29918
rect 145196 29854 145248 29860
rect 145012 20120 145064 20126
rect 145012 20062 145064 20068
rect 144552 16108 144604 16114
rect 144552 16050 144604 16056
rect 145472 11824 145524 11830
rect 145472 11766 145524 11772
rect 144736 3256 144788 3262
rect 144736 3198 144788 3204
rect 144460 3188 144512 3194
rect 144460 3130 144512 3136
rect 144748 480 144776 3198
rect 140014 354 140126 480
rect 139596 326 140126 354
rect 140014 -960 140126 326
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145484 354 145512 11766
rect 146312 3874 146340 73126
rect 146404 4010 146432 76463
rect 146392 4004 146444 4010
rect 146392 3946 146444 3952
rect 146496 3942 146524 76599
rect 146588 6798 146616 76735
rect 146668 76706 146720 76712
rect 146668 76628 146720 76634
rect 146668 76570 146720 76576
rect 146680 6866 146708 76570
rect 146668 6860 146720 6866
rect 146668 6802 146720 6808
rect 146576 6792 146628 6798
rect 146576 6734 146628 6740
rect 146772 6730 146800 79648
rect 146852 79630 146904 79636
rect 147034 79656 147090 79665
rect 146944 79620 146996 79626
rect 147034 79591 147090 79600
rect 146944 79562 146996 79568
rect 146852 76560 146904 76566
rect 146852 76502 146904 76508
rect 146864 9382 146892 76502
rect 146852 9376 146904 9382
rect 146852 9318 146904 9324
rect 146956 9314 146984 79562
rect 147048 77081 147076 79591
rect 147034 77072 147090 77081
rect 147034 77007 147090 77016
rect 147036 76900 147088 76906
rect 147036 76842 147088 76848
rect 147048 70394 147076 76842
rect 147140 76566 147168 79716
rect 147738 79744 147766 80036
rect 147496 79698 147548 79704
rect 147692 79716 147766 79744
rect 147312 79688 147364 79694
rect 147312 79630 147364 79636
rect 147404 79688 147456 79694
rect 147404 79630 147456 79636
rect 147220 79552 147272 79558
rect 147220 79494 147272 79500
rect 147128 76560 147180 76566
rect 147128 76502 147180 76508
rect 147232 73982 147260 79494
rect 147324 77897 147352 79630
rect 147310 77888 147366 77897
rect 147310 77823 147366 77832
rect 147416 75041 147444 79630
rect 147508 76945 147536 79698
rect 147692 79642 147720 79716
rect 147830 79676 147858 80036
rect 147922 79830 147950 80036
rect 147910 79824 147962 79830
rect 147910 79766 147962 79772
rect 148014 79744 148042 80036
rect 148106 79937 148134 80036
rect 148092 79928 148148 79937
rect 148092 79863 148148 79872
rect 148198 79744 148226 80036
rect 148290 79898 148318 80036
rect 148382 79898 148410 80036
rect 148278 79892 148330 79898
rect 148278 79834 148330 79840
rect 148370 79892 148422 79898
rect 148370 79834 148422 79840
rect 148324 79756 148376 79762
rect 148014 79716 148088 79744
rect 148198 79716 148272 79744
rect 147600 79614 147720 79642
rect 147784 79648 147858 79676
rect 147954 79656 148010 79665
rect 147600 78674 147628 79614
rect 147680 79552 147732 79558
rect 147680 79494 147732 79500
rect 147588 78668 147640 78674
rect 147588 78610 147640 78616
rect 147494 76936 147550 76945
rect 147494 76871 147550 76880
rect 147402 75032 147458 75041
rect 147402 74967 147458 74976
rect 147220 73976 147272 73982
rect 147220 73918 147272 73924
rect 147048 70366 147168 70394
rect 147140 64874 147168 70366
rect 147048 64846 147168 64874
rect 147048 9450 147076 64846
rect 147036 9444 147088 9450
rect 147036 9386 147088 9392
rect 146944 9308 146996 9314
rect 146944 9250 146996 9256
rect 146760 6724 146812 6730
rect 146760 6666 146812 6672
rect 146484 3936 146536 3942
rect 146484 3878 146536 3884
rect 146300 3868 146352 3874
rect 146300 3810 146352 3816
rect 147692 3806 147720 79494
rect 147784 76362 147812 79648
rect 147954 79591 148010 79600
rect 147772 76356 147824 76362
rect 147772 76298 147824 76304
rect 147772 75132 147824 75138
rect 147772 75074 147824 75080
rect 147784 5030 147812 75074
rect 147862 74488 147918 74497
rect 147862 74423 147918 74432
rect 147876 6662 147904 74423
rect 147968 14754 147996 79591
rect 148060 76906 148088 79716
rect 148140 79620 148192 79626
rect 148140 79562 148192 79568
rect 148048 76900 148100 76906
rect 148048 76842 148100 76848
rect 148048 76628 148100 76634
rect 148048 76570 148100 76576
rect 148060 24342 148088 76570
rect 148152 33930 148180 79562
rect 148244 35426 148272 79716
rect 148474 79744 148502 80036
rect 148566 79937 148594 80036
rect 148552 79928 148608 79937
rect 148552 79863 148608 79872
rect 148658 79744 148686 80036
rect 148324 79698 148376 79704
rect 148428 79716 148502 79744
rect 148612 79716 148686 79744
rect 148336 76634 148364 79698
rect 148324 76628 148376 76634
rect 148324 76570 148376 76576
rect 148324 76356 148376 76362
rect 148324 76298 148376 76304
rect 148336 42158 148364 76298
rect 148428 75138 148456 79716
rect 148508 79484 148560 79490
rect 148508 79426 148560 79432
rect 148416 75132 148468 75138
rect 148416 75074 148468 75080
rect 148520 74089 148548 79426
rect 148612 76838 148640 79716
rect 148750 79676 148778 80036
rect 148842 79744 148870 80036
rect 148934 79937 148962 80036
rect 148920 79928 148976 79937
rect 148920 79863 148976 79872
rect 149026 79801 149054 80036
rect 149012 79792 149068 79801
rect 148842 79716 148916 79744
rect 149012 79727 149068 79736
rect 148704 79648 148778 79676
rect 148600 76832 148652 76838
rect 148600 76774 148652 76780
rect 148506 74080 148562 74089
rect 148506 74015 148562 74024
rect 148704 72457 148732 79648
rect 148888 76673 148916 79716
rect 148968 79688 149020 79694
rect 149118 79676 149146 80036
rect 149210 79966 149238 80036
rect 149302 79966 149330 80036
rect 149198 79960 149250 79966
rect 149198 79902 149250 79908
rect 149290 79960 149342 79966
rect 149290 79902 149342 79908
rect 149394 79898 149422 80036
rect 149486 79898 149514 80036
rect 149578 79966 149606 80036
rect 149566 79960 149618 79966
rect 149670 79937 149698 80036
rect 149566 79902 149618 79908
rect 149656 79928 149712 79937
rect 149382 79892 149434 79898
rect 149382 79834 149434 79840
rect 149474 79892 149526 79898
rect 149656 79863 149712 79872
rect 149474 79834 149526 79840
rect 149610 79792 149666 79801
rect 149762 79778 149790 80036
rect 149854 79898 149882 80036
rect 149842 79892 149894 79898
rect 149842 79834 149894 79840
rect 149610 79727 149666 79736
rect 149716 79750 149790 79778
rect 149520 79688 149572 79694
rect 149118 79648 149192 79676
rect 148968 79630 149020 79636
rect 148874 76664 148930 76673
rect 148874 76599 148930 76608
rect 148980 73953 149008 79630
rect 149060 79416 149112 79422
rect 149060 79358 149112 79364
rect 148966 73944 149022 73953
rect 148966 73879 149022 73888
rect 148690 72448 148746 72457
rect 148690 72383 148746 72392
rect 148324 42152 148376 42158
rect 148324 42094 148376 42100
rect 148232 35420 148284 35426
rect 148232 35362 148284 35368
rect 148140 33924 148192 33930
rect 148140 33866 148192 33872
rect 148048 24336 148100 24342
rect 148048 24278 148100 24284
rect 148048 22840 148100 22846
rect 148048 22782 148100 22788
rect 147956 14748 148008 14754
rect 147956 14690 148008 14696
rect 147864 6656 147916 6662
rect 147864 6598 147916 6604
rect 147772 5024 147824 5030
rect 147772 4966 147824 4972
rect 147680 3800 147732 3806
rect 147680 3742 147732 3748
rect 147126 3632 147182 3641
rect 147126 3567 147182 3576
rect 147140 480 147168 3567
rect 145902 354 146014 480
rect 145484 326 146014 354
rect 145902 -960 146014 326
rect 147098 -960 147210 480
rect 148060 354 148088 22782
rect 149072 7886 149100 79358
rect 149164 76770 149192 79648
rect 149520 79630 149572 79636
rect 149244 79620 149296 79626
rect 149244 79562 149296 79568
rect 149256 77110 149284 79562
rect 149428 79552 149480 79558
rect 149428 79494 149480 79500
rect 149244 77104 149296 77110
rect 149244 77046 149296 77052
rect 149152 76764 149204 76770
rect 149152 76706 149204 76712
rect 149336 76696 149388 76702
rect 149336 76638 149388 76644
rect 149244 76560 149296 76566
rect 149244 76502 149296 76508
rect 149152 74452 149204 74458
rect 149152 74394 149204 74400
rect 149164 9246 149192 74394
rect 149256 14686 149284 76502
rect 149348 24274 149376 76638
rect 149440 25838 149468 79494
rect 149532 78402 149560 79630
rect 149520 78396 149572 78402
rect 149520 78338 149572 78344
rect 149520 77104 149572 77110
rect 149520 77046 149572 77052
rect 149532 35358 149560 77046
rect 149624 58818 149652 79727
rect 149716 76566 149744 79750
rect 149946 79744 149974 80036
rect 149900 79716 149974 79744
rect 150038 79744 150066 80036
rect 150130 79937 150158 80036
rect 150116 79928 150172 79937
rect 150116 79863 150172 79872
rect 150222 79744 150250 80036
rect 150314 79801 150342 80036
rect 150038 79716 150112 79744
rect 149796 79688 149848 79694
rect 149796 79630 149848 79636
rect 149704 76560 149756 76566
rect 149704 76502 149756 76508
rect 149808 73154 149836 79630
rect 149900 76702 149928 79716
rect 149980 79620 150032 79626
rect 149980 79562 150032 79568
rect 149888 76696 149940 76702
rect 149888 76638 149940 76644
rect 149716 73126 149836 73154
rect 149992 73154 150020 79562
rect 150084 74458 150112 79716
rect 150176 79716 150250 79744
rect 150300 79792 150356 79801
rect 150300 79727 150356 79736
rect 150176 75177 150204 79716
rect 150406 79676 150434 80036
rect 150498 79744 150526 80036
rect 150590 79903 150618 80036
rect 150576 79894 150632 79903
rect 150682 79898 150710 80036
rect 150576 79829 150632 79838
rect 150670 79892 150722 79898
rect 150670 79834 150722 79840
rect 150774 79744 150802 80036
rect 150866 79898 150894 80036
rect 150854 79892 150906 79898
rect 150854 79834 150906 79840
rect 150958 79744 150986 80036
rect 150498 79716 150710 79744
rect 150774 79716 150848 79744
rect 150360 79648 150434 79676
rect 150682 79676 150710 79716
rect 150530 79656 150586 79665
rect 150256 79620 150308 79626
rect 150256 79562 150308 79568
rect 150268 76702 150296 79562
rect 150256 76696 150308 76702
rect 150256 76638 150308 76644
rect 150162 75168 150218 75177
rect 150162 75103 150218 75112
rect 150072 74452 150124 74458
rect 150072 74394 150124 74400
rect 150360 73817 150388 79648
rect 150682 79648 150756 79676
rect 150530 79591 150586 79600
rect 150440 79552 150492 79558
rect 150440 79494 150492 79500
rect 150346 73808 150402 73817
rect 150346 73743 150402 73752
rect 149992 73126 150112 73154
rect 149716 72758 149744 73126
rect 150084 72826 150112 73126
rect 150072 72820 150124 72826
rect 150072 72762 150124 72768
rect 149704 72752 149756 72758
rect 149704 72694 149756 72700
rect 149612 58812 149664 58818
rect 149612 58754 149664 58760
rect 149520 35352 149572 35358
rect 149520 35294 149572 35300
rect 149428 25832 149480 25838
rect 149428 25774 149480 25780
rect 149336 24268 149388 24274
rect 149336 24210 149388 24216
rect 149244 14680 149296 14686
rect 149244 14622 149296 14628
rect 149152 9240 149204 9246
rect 149152 9182 149204 9188
rect 149060 7880 149112 7886
rect 149060 7822 149112 7828
rect 150452 7818 150480 79494
rect 150544 10470 150572 79591
rect 150624 79552 150676 79558
rect 150624 79494 150676 79500
rect 150636 29850 150664 79494
rect 150728 78062 150756 79648
rect 150820 78198 150848 79716
rect 150912 79716 150986 79744
rect 150808 78192 150860 78198
rect 150808 78134 150860 78140
rect 150716 78056 150768 78062
rect 150716 77998 150768 78004
rect 150912 76362 150940 79716
rect 151050 79676 151078 80036
rect 151142 79966 151170 80036
rect 151130 79960 151182 79966
rect 151130 79902 151182 79908
rect 151234 79898 151262 80036
rect 151326 79898 151354 80036
rect 151222 79892 151274 79898
rect 151222 79834 151274 79840
rect 151314 79892 151366 79898
rect 151314 79834 151366 79840
rect 151268 79756 151320 79762
rect 151004 79648 151078 79676
rect 151188 79716 151268 79744
rect 150900 76356 150952 76362
rect 150900 76298 150952 76304
rect 150716 75336 150768 75342
rect 150716 75278 150768 75284
rect 150728 31142 150756 75278
rect 150808 75268 150860 75274
rect 150808 75210 150860 75216
rect 150820 42090 150848 75210
rect 150900 75200 150952 75206
rect 150900 75142 150952 75148
rect 150912 54806 150940 75142
rect 151004 60246 151032 79648
rect 151188 78656 151216 79716
rect 151418 79744 151446 80036
rect 151510 79966 151538 80036
rect 151602 79966 151630 80036
rect 151498 79960 151550 79966
rect 151498 79902 151550 79908
rect 151590 79960 151642 79966
rect 151694 79937 151722 80036
rect 151590 79902 151642 79908
rect 151680 79928 151736 79937
rect 151680 79863 151736 79872
rect 151544 79824 151596 79830
rect 151544 79766 151596 79772
rect 151418 79716 151492 79744
rect 151268 79698 151320 79704
rect 151360 79620 151412 79626
rect 151360 79562 151412 79568
rect 151268 79484 151320 79490
rect 151268 79426 151320 79432
rect 151096 78628 151216 78656
rect 151096 75342 151124 78628
rect 151176 78192 151228 78198
rect 151176 78134 151228 78140
rect 151084 75336 151136 75342
rect 151084 75278 151136 75284
rect 151188 70394 151216 78134
rect 151280 75274 151308 79426
rect 151268 75268 151320 75274
rect 151268 75210 151320 75216
rect 151372 75206 151400 79562
rect 151464 77450 151492 79716
rect 151556 78713 151584 79766
rect 151636 79756 151688 79762
rect 151786 79744 151814 80036
rect 151878 79830 151906 80036
rect 151970 79966 151998 80036
rect 152062 79971 152090 80036
rect 151958 79960 152010 79966
rect 151958 79902 152010 79908
rect 152048 79962 152104 79971
rect 152048 79897 152104 79906
rect 151866 79824 151918 79830
rect 151866 79766 151918 79772
rect 152002 79792 152058 79801
rect 151636 79698 151688 79704
rect 151740 79716 151814 79744
rect 152002 79727 152058 79736
rect 151542 78704 151598 78713
rect 151542 78639 151598 78648
rect 151648 77625 151676 79698
rect 151740 78849 151768 79716
rect 152016 79694 152044 79727
rect 152004 79688 152056 79694
rect 151910 79656 151966 79665
rect 152154 79676 152182 80036
rect 152246 79898 152274 80036
rect 152234 79892 152286 79898
rect 152234 79834 152286 79840
rect 152338 79778 152366 80036
rect 152430 79971 152458 80036
rect 152416 79962 152472 79971
rect 152522 79966 152550 80036
rect 152416 79897 152472 79906
rect 152510 79960 152562 79966
rect 152510 79902 152562 79908
rect 152614 79898 152642 80036
rect 152706 79966 152734 80036
rect 152694 79960 152746 79966
rect 152694 79902 152746 79908
rect 152602 79892 152654 79898
rect 152602 79834 152654 79840
rect 152338 79762 152412 79778
rect 152338 79756 152424 79762
rect 152338 79750 152372 79756
rect 152372 79698 152424 79704
rect 152648 79756 152700 79762
rect 152648 79698 152700 79704
rect 152004 79630 152056 79636
rect 152108 79648 152182 79676
rect 152280 79688 152332 79694
rect 151910 79591 151912 79600
rect 151964 79591 151966 79600
rect 151912 79562 151964 79568
rect 152108 79506 152136 79648
rect 152556 79688 152608 79694
rect 152462 79656 152518 79665
rect 152280 79630 152332 79636
rect 152016 79478 152136 79506
rect 151912 79348 151964 79354
rect 151912 79290 151964 79296
rect 151726 78840 151782 78849
rect 151726 78775 151782 78784
rect 151634 77616 151690 77625
rect 151634 77551 151690 77560
rect 151726 77480 151782 77489
rect 151452 77444 151504 77450
rect 151726 77415 151782 77424
rect 151452 77386 151504 77392
rect 151452 76356 151504 76362
rect 151452 76298 151504 76304
rect 151360 75200 151412 75206
rect 151360 75142 151412 75148
rect 151464 72690 151492 76298
rect 151452 72684 151504 72690
rect 151452 72626 151504 72632
rect 151740 72622 151768 77415
rect 151820 77308 151872 77314
rect 151820 77250 151872 77256
rect 151728 72616 151780 72622
rect 151728 72558 151780 72564
rect 151096 70366 151216 70394
rect 151096 62898 151124 70366
rect 151084 62892 151136 62898
rect 151084 62834 151136 62840
rect 150992 60240 151044 60246
rect 150992 60182 151044 60188
rect 150900 54800 150952 54806
rect 150900 54742 150952 54748
rect 150808 42084 150860 42090
rect 150808 42026 150860 42032
rect 150716 31136 150768 31142
rect 150716 31078 150768 31084
rect 150624 29844 150676 29850
rect 150624 29786 150676 29792
rect 151832 13258 151860 77250
rect 151924 16046 151952 79290
rect 152016 77858 152044 79478
rect 152096 79416 152148 79422
rect 152096 79358 152148 79364
rect 152004 77852 152056 77858
rect 152004 77794 152056 77800
rect 152004 77240 152056 77246
rect 152004 77182 152056 77188
rect 152016 28422 152044 77182
rect 152108 37942 152136 79358
rect 152188 75132 152240 75138
rect 152188 75074 152240 75080
rect 152200 43518 152228 75074
rect 152292 45014 152320 79630
rect 152384 79614 152462 79642
rect 152384 57526 152412 79614
rect 152556 79630 152608 79636
rect 152462 79591 152518 79600
rect 152464 79416 152516 79422
rect 152464 79358 152516 79364
rect 152476 79150 152504 79358
rect 152464 79144 152516 79150
rect 152464 79086 152516 79092
rect 152568 78826 152596 79630
rect 152476 78798 152596 78826
rect 152476 77246 152504 78798
rect 152556 77852 152608 77858
rect 152556 77794 152608 77800
rect 152464 77240 152516 77246
rect 152464 77182 152516 77188
rect 152464 77104 152516 77110
rect 152464 77046 152516 77052
rect 152476 76702 152504 77046
rect 152464 76696 152516 76702
rect 152464 76638 152516 76644
rect 152464 76560 152516 76566
rect 152464 76502 152516 76508
rect 152476 72486 152504 76502
rect 152464 72480 152516 72486
rect 152464 72422 152516 72428
rect 152568 70394 152596 77794
rect 152660 75138 152688 79698
rect 152798 79676 152826 80036
rect 152890 79801 152918 80036
rect 152982 79830 153010 80036
rect 153074 79971 153102 80036
rect 153060 79962 153116 79971
rect 153060 79897 153116 79906
rect 152970 79824 153022 79830
rect 152876 79792 152932 79801
rect 152970 79766 153022 79772
rect 152876 79727 152932 79736
rect 152752 79648 152826 79676
rect 153166 79676 153194 80036
rect 153258 79971 153286 80036
rect 153244 79962 153300 79971
rect 153350 79966 153378 80036
rect 153442 79971 153470 80036
rect 153244 79897 153300 79906
rect 153338 79960 153390 79966
rect 153338 79902 153390 79908
rect 153428 79962 153484 79971
rect 153534 79966 153562 80036
rect 153428 79897 153484 79906
rect 153522 79960 153574 79966
rect 153522 79902 153574 79908
rect 153626 79778 153654 80036
rect 153718 79966 153746 80036
rect 153706 79960 153758 79966
rect 153706 79902 153758 79908
rect 153810 79778 153838 80036
rect 153902 79898 153930 80036
rect 153890 79892 153942 79898
rect 153890 79834 153942 79840
rect 153580 79750 153654 79778
rect 153764 79750 153838 79778
rect 153166 79648 153240 79676
rect 152752 77314 152780 79648
rect 152832 79552 152884 79558
rect 152832 79494 152884 79500
rect 153016 79552 153068 79558
rect 153016 79494 153068 79500
rect 152844 78010 152872 79494
rect 152924 79484 152976 79490
rect 152924 79426 152976 79432
rect 152936 78946 152964 79426
rect 152924 78940 152976 78946
rect 152924 78882 152976 78888
rect 152844 77982 152964 78010
rect 152832 77920 152884 77926
rect 152832 77862 152884 77868
rect 152740 77308 152792 77314
rect 152740 77250 152792 77256
rect 152740 77172 152792 77178
rect 152740 77114 152792 77120
rect 152752 76634 152780 77114
rect 152740 76628 152792 76634
rect 152740 76570 152792 76576
rect 152844 75546 152872 77862
rect 152936 76566 152964 77982
rect 153028 77353 153056 79494
rect 153108 79348 153160 79354
rect 153108 79290 153160 79296
rect 153120 79014 153148 79290
rect 153108 79008 153160 79014
rect 153108 78950 153160 78956
rect 153212 78470 153240 79648
rect 153476 79620 153528 79626
rect 153476 79562 153528 79568
rect 153292 79552 153344 79558
rect 153292 79494 153344 79500
rect 153200 78464 153252 78470
rect 153200 78406 153252 78412
rect 153198 78024 153254 78033
rect 153198 77959 153254 77968
rect 153014 77344 153070 77353
rect 153014 77279 153070 77288
rect 152924 76560 152976 76566
rect 152924 76502 152976 76508
rect 152832 75540 152884 75546
rect 152832 75482 152884 75488
rect 152648 75132 152700 75138
rect 152648 75074 152700 75080
rect 152476 70366 152596 70394
rect 153212 70394 153240 77959
rect 153304 73914 153332 79494
rect 153384 75948 153436 75954
rect 153384 75890 153436 75896
rect 153292 73908 153344 73914
rect 153292 73850 153344 73856
rect 153212 70366 153332 70394
rect 152476 58750 152504 70366
rect 152464 58744 152516 58750
rect 152464 58686 152516 58692
rect 152372 57520 152424 57526
rect 152372 57462 152424 57468
rect 152280 45008 152332 45014
rect 152280 44950 152332 44956
rect 152188 43512 152240 43518
rect 152188 43454 152240 43460
rect 152462 43480 152518 43489
rect 152462 43415 152518 43424
rect 152096 37936 152148 37942
rect 152096 37878 152148 37884
rect 152004 28416 152056 28422
rect 152004 28358 152056 28364
rect 151912 16040 151964 16046
rect 151912 15982 151964 15988
rect 151820 13252 151872 13258
rect 151820 13194 151872 13200
rect 150532 10464 150584 10470
rect 150532 10406 150584 10412
rect 150440 7812 150492 7818
rect 150440 7754 150492 7760
rect 152476 3602 152504 43415
rect 153304 9178 153332 70366
rect 153396 15978 153424 75890
rect 153488 49230 153516 79562
rect 153580 75954 153608 79750
rect 153660 79688 153712 79694
rect 153660 79630 153712 79636
rect 153568 75948 153620 75954
rect 153568 75890 153620 75896
rect 153672 75478 153700 79630
rect 153660 75472 153712 75478
rect 153660 75414 153712 75420
rect 153568 75132 153620 75138
rect 153568 75074 153620 75080
rect 153580 55962 153608 75074
rect 153764 70394 153792 79750
rect 153994 79744 154022 80036
rect 154086 79778 154114 80036
rect 154178 79898 154206 80036
rect 154166 79892 154218 79898
rect 154166 79834 154218 79840
rect 154086 79750 154160 79778
rect 153948 79716 154022 79744
rect 153844 79688 153896 79694
rect 153844 79630 153896 79636
rect 153856 77976 153884 79630
rect 153948 78169 153976 79716
rect 154028 79620 154080 79626
rect 154028 79562 154080 79568
rect 154040 79082 154068 79562
rect 154028 79076 154080 79082
rect 154028 79018 154080 79024
rect 153934 78160 153990 78169
rect 153934 78095 153990 78104
rect 153856 77948 153976 77976
rect 153844 77444 153896 77450
rect 153844 77386 153896 77392
rect 153672 70366 153792 70394
rect 153856 70394 153884 77386
rect 153948 75018 153976 77948
rect 154132 75138 154160 79750
rect 154270 79744 154298 80036
rect 154362 79937 154390 80036
rect 154348 79928 154404 79937
rect 154348 79863 154404 79872
rect 154454 79812 154482 80036
rect 154224 79716 154298 79744
rect 154408 79784 154482 79812
rect 154546 79801 154574 80036
rect 154532 79792 154588 79801
rect 154224 77994 154252 79716
rect 154304 79620 154356 79626
rect 154304 79562 154356 79568
rect 154212 77988 154264 77994
rect 154212 77930 154264 77936
rect 154316 77246 154344 79562
rect 154408 77897 154436 79784
rect 154532 79727 154588 79736
rect 154638 79744 154666 80036
rect 154730 79898 154758 80036
rect 154718 79892 154770 79898
rect 154718 79834 154770 79840
rect 154822 79812 154850 80036
rect 154914 79966 154942 80036
rect 154902 79960 154954 79966
rect 154902 79902 154954 79908
rect 154822 79784 154896 79812
rect 154638 79716 154712 79744
rect 154684 79665 154712 79716
rect 154486 79656 154542 79665
rect 154670 79656 154726 79665
rect 154486 79591 154542 79600
rect 154580 79620 154632 79626
rect 154394 77888 154450 77897
rect 154394 77823 154450 77832
rect 154500 77704 154528 79591
rect 154868 79608 154896 79784
rect 155006 79744 155034 80036
rect 154670 79591 154726 79600
rect 154580 79562 154632 79568
rect 154776 79580 154896 79608
rect 154960 79716 155034 79744
rect 154592 77790 154620 79562
rect 154672 78804 154724 78810
rect 154672 78746 154724 78752
rect 154580 77784 154632 77790
rect 154580 77726 154632 77732
rect 154408 77676 154528 77704
rect 154304 77240 154356 77246
rect 154304 77182 154356 77188
rect 154408 76702 154436 77676
rect 154486 77616 154542 77625
rect 154486 77551 154542 77560
rect 154396 76696 154448 76702
rect 154396 76638 154448 76644
rect 154120 75132 154172 75138
rect 154120 75074 154172 75080
rect 153948 74990 154252 75018
rect 154224 70394 154252 74990
rect 154500 72554 154528 77551
rect 154580 75336 154632 75342
rect 154580 75278 154632 75284
rect 154488 72548 154540 72554
rect 154488 72490 154540 72496
rect 153856 70366 154160 70394
rect 154224 70366 154436 70394
rect 153672 64326 153700 70366
rect 153660 64320 153712 64326
rect 153660 64262 153712 64268
rect 153568 55956 153620 55962
rect 153568 55898 153620 55904
rect 153476 49224 153528 49230
rect 153476 49166 153528 49172
rect 154132 31210 154160 70366
rect 154120 31204 154172 31210
rect 154120 31146 154172 31152
rect 153384 15972 153436 15978
rect 153384 15914 153436 15920
rect 153292 9172 153344 9178
rect 153292 9114 153344 9120
rect 154212 5228 154264 5234
rect 154212 5170 154264 5176
rect 151820 3596 151872 3602
rect 151820 3538 151872 3544
rect 152464 3596 152516 3602
rect 152464 3538 152516 3544
rect 149520 3392 149572 3398
rect 149520 3334 149572 3340
rect 149532 480 149560 3334
rect 150624 3324 150676 3330
rect 150624 3266 150676 3272
rect 150636 480 150664 3266
rect 151832 480 151860 3538
rect 153016 3392 153068 3398
rect 153016 3334 153068 3340
rect 153028 480 153056 3334
rect 154224 480 154252 5170
rect 154408 4962 154436 70366
rect 154592 7750 154620 75278
rect 154684 10402 154712 78746
rect 154776 78266 154804 79580
rect 154960 79506 154988 79716
rect 155098 79676 155126 80036
rect 154868 79478 154988 79506
rect 155052 79648 155126 79676
rect 155190 79676 155218 80036
rect 155282 79801 155310 80036
rect 155268 79792 155324 79801
rect 155268 79727 155324 79736
rect 155374 79676 155402 80036
rect 155466 79966 155494 80036
rect 155454 79960 155506 79966
rect 155454 79902 155506 79908
rect 155558 79812 155586 80036
rect 155190 79648 155264 79676
rect 154764 78260 154816 78266
rect 154764 78202 154816 78208
rect 154764 77920 154816 77926
rect 154764 77862 154816 77868
rect 154776 14618 154804 77862
rect 154868 28354 154896 79478
rect 154948 79348 155000 79354
rect 154948 79290 155000 79296
rect 154960 78946 154988 79290
rect 154948 78940 155000 78946
rect 154948 78882 155000 78888
rect 155052 78810 155080 79648
rect 155132 79552 155184 79558
rect 155132 79494 155184 79500
rect 155040 78804 155092 78810
rect 155040 78746 155092 78752
rect 155038 78704 155094 78713
rect 155038 78639 155094 78648
rect 155052 75682 155080 78639
rect 155040 75676 155092 75682
rect 155040 75618 155092 75624
rect 154948 75268 155000 75274
rect 154948 75210 155000 75216
rect 154960 54738 154988 75210
rect 155040 75200 155092 75206
rect 155040 75142 155092 75148
rect 155052 58682 155080 75142
rect 155144 64190 155172 79494
rect 155236 75274 155264 79648
rect 155328 79648 155402 79676
rect 155512 79784 155586 79812
rect 155328 78198 155356 79648
rect 155408 79552 155460 79558
rect 155408 79494 155460 79500
rect 155316 78192 155368 78198
rect 155316 78134 155368 78140
rect 155316 75676 155368 75682
rect 155316 75618 155368 75624
rect 155224 75268 155276 75274
rect 155224 75210 155276 75216
rect 155328 71330 155356 75618
rect 155420 75206 155448 79494
rect 155512 75342 155540 79784
rect 155650 79744 155678 80036
rect 155742 79778 155770 80036
rect 155834 79966 155862 80036
rect 155926 79966 155954 80036
rect 155822 79960 155874 79966
rect 155822 79902 155874 79908
rect 155914 79960 155966 79966
rect 155914 79902 155966 79908
rect 155868 79824 155920 79830
rect 155742 79750 155816 79778
rect 156018 79778 156046 80036
rect 155868 79766 155920 79772
rect 155604 79716 155678 79744
rect 155604 77926 155632 79716
rect 155684 79416 155736 79422
rect 155684 79358 155736 79364
rect 155696 79218 155724 79358
rect 155684 79212 155736 79218
rect 155684 79154 155736 79160
rect 155592 77920 155644 77926
rect 155592 77862 155644 77868
rect 155788 77353 155816 79750
rect 155880 78606 155908 79766
rect 155972 79750 156046 79778
rect 155972 78826 156000 79750
rect 156110 79608 156138 80036
rect 156202 79676 156230 80036
rect 156294 79966 156322 80036
rect 156386 79966 156414 80036
rect 156282 79960 156334 79966
rect 156282 79902 156334 79908
rect 156374 79960 156426 79966
rect 156374 79902 156426 79908
rect 156478 79898 156506 80036
rect 156466 79892 156518 79898
rect 156466 79834 156518 79840
rect 156570 79830 156598 80036
rect 156558 79824 156610 79830
rect 156418 79792 156474 79801
rect 156558 79766 156610 79772
rect 156418 79727 156474 79736
rect 156202 79648 156276 79676
rect 156110 79580 156184 79608
rect 155972 78798 156092 78826
rect 155960 78736 156012 78742
rect 155960 78678 156012 78684
rect 155868 78600 155920 78606
rect 155868 78542 155920 78548
rect 155774 77344 155830 77353
rect 155774 77279 155830 77288
rect 155776 77240 155828 77246
rect 155776 77182 155828 77188
rect 155592 75472 155644 75478
rect 155592 75414 155644 75420
rect 155500 75336 155552 75342
rect 155500 75278 155552 75284
rect 155408 75200 155460 75206
rect 155408 75142 155460 75148
rect 155316 71324 155368 71330
rect 155316 71266 155368 71272
rect 155604 70394 155632 75414
rect 155604 70366 155724 70394
rect 155132 64184 155184 64190
rect 155132 64126 155184 64132
rect 155040 58676 155092 58682
rect 155040 58618 155092 58624
rect 154948 54732 155000 54738
rect 154948 54674 155000 54680
rect 154856 28348 154908 28354
rect 154856 28290 154908 28296
rect 154764 14612 154816 14618
rect 154764 14554 154816 14560
rect 155696 13190 155724 70366
rect 155788 65550 155816 77182
rect 155776 65544 155828 65550
rect 155776 65486 155828 65492
rect 155684 13184 155736 13190
rect 155684 13126 155736 13132
rect 154672 10396 154724 10402
rect 154672 10338 154724 10344
rect 154580 7744 154632 7750
rect 154580 7686 154632 7692
rect 155972 6594 156000 78678
rect 156064 75342 156092 78798
rect 156052 75336 156104 75342
rect 156052 75278 156104 75284
rect 156052 75200 156104 75206
rect 156052 75142 156104 75148
rect 156156 75154 156184 79580
rect 156248 78742 156276 79648
rect 156432 79626 156460 79727
rect 156512 79688 156564 79694
rect 156662 79676 156690 80036
rect 156754 79830 156782 80036
rect 156742 79824 156794 79830
rect 156742 79766 156794 79772
rect 156846 79744 156874 80036
rect 156938 79812 156966 80036
rect 157030 79966 157058 80036
rect 157018 79960 157070 79966
rect 157122 79937 157150 80036
rect 157018 79902 157070 79908
rect 157108 79928 157164 79937
rect 157108 79863 157164 79872
rect 157064 79824 157116 79830
rect 156938 79784 157012 79812
rect 156846 79716 156920 79744
rect 156662 79648 156828 79676
rect 156512 79630 156564 79636
rect 156328 79620 156380 79626
rect 156328 79562 156380 79568
rect 156420 79620 156472 79626
rect 156420 79562 156472 79568
rect 156236 78736 156288 78742
rect 156236 78678 156288 78684
rect 156236 78464 156288 78470
rect 156236 78406 156288 78412
rect 156248 76809 156276 78406
rect 156234 76800 156290 76809
rect 156234 76735 156290 76744
rect 156340 75274 156368 79562
rect 156420 79484 156472 79490
rect 156420 79426 156472 79432
rect 156328 75268 156380 75274
rect 156328 75210 156380 75216
rect 156064 11830 156092 75142
rect 156156 75126 156368 75154
rect 156236 75064 156288 75070
rect 156236 75006 156288 75012
rect 156144 74996 156196 75002
rect 156144 74938 156196 74944
rect 156156 25770 156184 74938
rect 156248 26994 156276 75006
rect 156340 29782 156368 75126
rect 156432 54670 156460 79426
rect 156524 77294 156552 79630
rect 156524 77266 156736 77294
rect 156604 75336 156656 75342
rect 156604 75278 156656 75284
rect 156512 75268 156564 75274
rect 156512 75210 156564 75216
rect 156524 57458 156552 75210
rect 156616 61538 156644 75278
rect 156708 67046 156736 77266
rect 156800 75070 156828 79648
rect 156788 75064 156840 75070
rect 156788 75006 156840 75012
rect 156892 75002 156920 79716
rect 156984 79558 157012 79784
rect 157214 79801 157242 80036
rect 157306 79898 157334 80036
rect 157398 79898 157426 80036
rect 157294 79892 157346 79898
rect 157294 79834 157346 79840
rect 157386 79892 157438 79898
rect 157386 79834 157438 79840
rect 157064 79766 157116 79772
rect 157200 79792 157256 79801
rect 156972 79552 157024 79558
rect 156972 79494 157024 79500
rect 156972 79416 157024 79422
rect 156972 79358 157024 79364
rect 156984 75206 157012 79358
rect 157076 77926 157104 79766
rect 157200 79727 157256 79736
rect 157490 79744 157518 80036
rect 157582 79966 157610 80036
rect 157570 79960 157622 79966
rect 157570 79902 157622 79908
rect 157674 79898 157702 80036
rect 157766 79898 157794 80036
rect 157662 79892 157714 79898
rect 157662 79834 157714 79840
rect 157754 79892 157806 79898
rect 157754 79834 157806 79840
rect 157858 79744 157886 80036
rect 157490 79716 157564 79744
rect 157156 79688 157208 79694
rect 157156 79630 157208 79636
rect 157340 79688 157392 79694
rect 157340 79630 157392 79636
rect 157168 78033 157196 79630
rect 157248 79552 157300 79558
rect 157248 79494 157300 79500
rect 157260 78849 157288 79494
rect 157246 78840 157302 78849
rect 157246 78775 157302 78784
rect 157248 78056 157300 78062
rect 157154 78024 157210 78033
rect 157248 77998 157300 78004
rect 157154 77959 157210 77968
rect 157064 77920 157116 77926
rect 157064 77862 157116 77868
rect 156972 75200 157024 75206
rect 156972 75142 157024 75148
rect 156880 74996 156932 75002
rect 156880 74938 156932 74944
rect 157260 70394 157288 77998
rect 157352 75682 157380 79630
rect 157432 79620 157484 79626
rect 157432 79562 157484 79568
rect 157444 77858 157472 79562
rect 157432 77852 157484 77858
rect 157432 77794 157484 77800
rect 157536 75914 157564 79716
rect 157812 79716 157886 79744
rect 157708 79552 157760 79558
rect 157708 79494 157760 79500
rect 157616 79484 157668 79490
rect 157616 79426 157668 79432
rect 157444 75886 157564 75914
rect 157340 75676 157392 75682
rect 157340 75618 157392 75624
rect 157340 75404 157392 75410
rect 157340 75346 157392 75352
rect 157168 70366 157288 70394
rect 157168 68474 157196 70366
rect 157156 68468 157208 68474
rect 157156 68410 157208 68416
rect 156696 67040 156748 67046
rect 156696 66982 156748 66988
rect 156604 61532 156656 61538
rect 156604 61474 156656 61480
rect 156512 57452 156564 57458
rect 156512 57394 156564 57400
rect 156420 54664 156472 54670
rect 156420 54606 156472 54612
rect 156328 29776 156380 29782
rect 156328 29718 156380 29724
rect 156236 26988 156288 26994
rect 156236 26930 156288 26936
rect 156144 25764 156196 25770
rect 156144 25706 156196 25712
rect 157352 19990 157380 75346
rect 157444 22982 157472 75886
rect 157524 75200 157576 75206
rect 157524 75142 157576 75148
rect 157536 24206 157564 75142
rect 157628 25702 157656 79426
rect 157720 78470 157748 79494
rect 157708 78464 157760 78470
rect 157708 78406 157760 78412
rect 157812 77976 157840 79716
rect 157950 79676 157978 80036
rect 157720 77948 157840 77976
rect 157904 79648 157978 79676
rect 157720 75410 157748 77948
rect 157904 77294 157932 79648
rect 158042 79540 158070 80036
rect 158134 79898 158162 80036
rect 158226 79966 158254 80036
rect 158214 79960 158266 79966
rect 158214 79902 158266 79908
rect 158122 79892 158174 79898
rect 158122 79834 158174 79840
rect 158318 79801 158346 80036
rect 158410 79971 158438 80036
rect 158396 79962 158452 79971
rect 158396 79897 158452 79906
rect 158502 79898 158530 80036
rect 158594 79898 158622 80036
rect 158490 79892 158542 79898
rect 158490 79834 158542 79840
rect 158582 79892 158634 79898
rect 158582 79834 158634 79840
rect 158304 79792 158360 79801
rect 158168 79756 158220 79762
rect 158304 79727 158360 79736
rect 158444 79756 158496 79762
rect 158168 79698 158220 79704
rect 158444 79698 158496 79704
rect 157996 79512 158070 79540
rect 157996 78810 158024 79512
rect 157984 78804 158036 78810
rect 157984 78746 158036 78752
rect 157984 78600 158036 78606
rect 157984 78542 158036 78548
rect 157812 77266 157932 77294
rect 157708 75404 157760 75410
rect 157708 75346 157760 75352
rect 157708 75268 157760 75274
rect 157708 75210 157760 75216
rect 157720 53378 157748 75210
rect 157812 55894 157840 77266
rect 157892 75676 157944 75682
rect 157892 75618 157944 75624
rect 157904 71262 157932 75618
rect 157996 73846 158024 78542
rect 158076 78464 158128 78470
rect 158076 78406 158128 78412
rect 157984 73840 158036 73846
rect 157984 73782 158036 73788
rect 157892 71256 157944 71262
rect 157892 71198 157944 71204
rect 158088 70394 158116 78406
rect 158180 75274 158208 79698
rect 158260 79688 158312 79694
rect 158260 79630 158312 79636
rect 158352 79688 158404 79694
rect 158352 79630 158404 79636
rect 158272 78928 158300 79630
rect 158364 79150 158392 79630
rect 158352 79144 158404 79150
rect 158352 79086 158404 79092
rect 158272 78900 158392 78928
rect 158260 78804 158312 78810
rect 158260 78746 158312 78752
rect 158168 75268 158220 75274
rect 158168 75210 158220 75216
rect 158272 75206 158300 78746
rect 158364 77382 158392 78900
rect 158456 78033 158484 79698
rect 158536 79688 158588 79694
rect 158686 79676 158714 80036
rect 158778 79966 158806 80036
rect 158870 79966 158898 80036
rect 158766 79960 158818 79966
rect 158766 79902 158818 79908
rect 158858 79960 158910 79966
rect 158858 79902 158910 79908
rect 158962 79830 158990 80036
rect 159054 79966 159082 80036
rect 159042 79960 159094 79966
rect 159042 79902 159094 79908
rect 158812 79824 158864 79830
rect 158812 79766 158864 79772
rect 158950 79824 159002 79830
rect 159146 79812 159174 80036
rect 159238 79898 159266 80036
rect 159330 79966 159358 80036
rect 159422 79971 159450 80036
rect 159318 79960 159370 79966
rect 159318 79902 159370 79908
rect 159408 79962 159464 79971
rect 159226 79892 159278 79898
rect 159408 79897 159464 79906
rect 159226 79834 159278 79840
rect 159100 79801 159174 79812
rect 158950 79766 159002 79772
rect 159086 79792 159174 79801
rect 158686 79648 158760 79676
rect 158536 79630 158588 79636
rect 158442 78024 158498 78033
rect 158442 77959 158498 77968
rect 158548 77897 158576 79630
rect 158534 77888 158590 77897
rect 158534 77823 158590 77832
rect 158628 77784 158680 77790
rect 158628 77726 158680 77732
rect 158352 77376 158404 77382
rect 158352 77318 158404 77324
rect 158260 75200 158312 75206
rect 158260 75142 158312 75148
rect 158640 70394 158668 77726
rect 158732 77489 158760 79648
rect 158718 77480 158774 77489
rect 158718 77415 158774 77424
rect 158824 77314 158852 79766
rect 159142 79784 159174 79792
rect 159270 79792 159326 79801
rect 159086 79727 159142 79736
rect 159326 79750 159404 79778
rect 159270 79727 159326 79736
rect 158904 79688 158956 79694
rect 158904 79630 158956 79636
rect 158812 77308 158864 77314
rect 158812 77250 158864 77256
rect 157904 70366 158116 70394
rect 158364 70366 158668 70394
rect 157904 61470 157932 70366
rect 158364 64258 158392 70366
rect 158352 64252 158404 64258
rect 158352 64194 158404 64200
rect 157892 61464 157944 61470
rect 157892 61406 157944 61412
rect 157800 55888 157852 55894
rect 157800 55830 157852 55836
rect 157708 53372 157760 53378
rect 157708 53314 157760 53320
rect 158916 33862 158944 79630
rect 159272 79620 159324 79626
rect 159272 79562 159324 79568
rect 159180 79552 159232 79558
rect 159180 79494 159232 79500
rect 158996 79144 159048 79150
rect 159192 79098 159220 79494
rect 158996 79086 159048 79092
rect 159008 78033 159036 79086
rect 159100 79070 159220 79098
rect 158994 78024 159050 78033
rect 158994 77959 159050 77968
rect 158996 77308 159048 77314
rect 158996 77250 159048 77256
rect 159008 46238 159036 77250
rect 159100 57390 159128 79070
rect 159180 79008 159232 79014
rect 159180 78950 159232 78956
rect 159192 78130 159220 78950
rect 159180 78124 159232 78130
rect 159180 78066 159232 78072
rect 159284 77790 159312 79562
rect 159272 77784 159324 77790
rect 159272 77726 159324 77732
rect 159180 77716 159232 77722
rect 159180 77658 159232 77664
rect 159192 77450 159220 77658
rect 159272 77648 159324 77654
rect 159272 77590 159324 77596
rect 159180 77444 159232 77450
rect 159180 77386 159232 77392
rect 159178 77344 159234 77353
rect 159284 77314 159312 77590
rect 159178 77279 159234 77288
rect 159272 77308 159324 77314
rect 159192 61402 159220 77279
rect 159272 77250 159324 77256
rect 159272 76628 159324 76634
rect 159272 76570 159324 76576
rect 159284 69902 159312 76570
rect 159376 69970 159404 79750
rect 159514 79744 159542 80036
rect 159606 79898 159634 80036
rect 159698 79966 159726 80036
rect 159790 79966 159818 80036
rect 159882 79971 159910 80036
rect 159686 79960 159738 79966
rect 159686 79902 159738 79908
rect 159778 79960 159830 79966
rect 159778 79902 159830 79908
rect 159868 79962 159924 79971
rect 159594 79892 159646 79898
rect 159868 79897 159924 79906
rect 159594 79834 159646 79840
rect 159974 79812 160002 80036
rect 160066 79966 160094 80036
rect 160158 79966 160186 80036
rect 160250 79966 160278 80036
rect 160342 79966 160370 80036
rect 160434 79966 160462 80036
rect 160054 79960 160106 79966
rect 160054 79902 160106 79908
rect 160146 79960 160198 79966
rect 160146 79902 160198 79908
rect 160238 79960 160290 79966
rect 160238 79902 160290 79908
rect 160330 79960 160382 79966
rect 160330 79902 160382 79908
rect 160422 79960 160474 79966
rect 160526 79937 160554 80036
rect 160618 79966 160646 80036
rect 160710 79966 160738 80036
rect 160606 79960 160658 79966
rect 160422 79902 160474 79908
rect 160512 79928 160568 79937
rect 160606 79902 160658 79908
rect 160698 79960 160750 79966
rect 160698 79902 160750 79908
rect 160512 79863 160568 79872
rect 160192 79824 160244 79830
rect 159974 79784 160048 79812
rect 159468 79716 159542 79744
rect 159640 79756 159692 79762
rect 159468 76158 159496 79716
rect 159640 79698 159692 79704
rect 159548 79620 159600 79626
rect 159548 79562 159600 79568
rect 159560 76634 159588 79562
rect 159548 76628 159600 76634
rect 159548 76570 159600 76576
rect 159456 76152 159508 76158
rect 159456 76094 159508 76100
rect 159652 75750 159680 79698
rect 159824 79552 159876 79558
rect 159824 79494 159876 79500
rect 159732 79484 159784 79490
rect 159732 79426 159784 79432
rect 159744 79150 159772 79426
rect 159732 79144 159784 79150
rect 159732 79086 159784 79092
rect 159732 78804 159784 78810
rect 159732 78746 159784 78752
rect 159744 78402 159772 78746
rect 159732 78396 159784 78402
rect 159732 78338 159784 78344
rect 159732 78192 159784 78198
rect 159836 78169 159864 79494
rect 159916 79484 159968 79490
rect 159916 79426 159968 79432
rect 159928 78713 159956 79426
rect 159914 78704 159970 78713
rect 159914 78639 159970 78648
rect 159914 78568 159970 78577
rect 159914 78503 159970 78512
rect 159732 78134 159784 78140
rect 159822 78160 159878 78169
rect 159640 75744 159692 75750
rect 159640 75686 159692 75692
rect 159364 69964 159416 69970
rect 159364 69906 159416 69912
rect 159272 69896 159324 69902
rect 159272 69838 159324 69844
rect 159180 61396 159232 61402
rect 159180 61338 159232 61344
rect 159088 57384 159140 57390
rect 159088 57326 159140 57332
rect 159744 49162 159772 78134
rect 159822 78095 159878 78104
rect 159824 76152 159876 76158
rect 159824 76094 159876 76100
rect 159732 49156 159784 49162
rect 159732 49098 159784 49104
rect 158996 46232 159048 46238
rect 158996 46174 159048 46180
rect 158904 33856 158956 33862
rect 158904 33798 158956 33804
rect 157616 25696 157668 25702
rect 157616 25638 157668 25644
rect 157524 24200 157576 24206
rect 157524 24142 157576 24148
rect 157432 22976 157484 22982
rect 157432 22918 157484 22924
rect 157340 19984 157392 19990
rect 157340 19926 157392 19932
rect 156052 11824 156104 11830
rect 156052 11766 156104 11772
rect 155960 6588 156012 6594
rect 155960 6530 156012 6536
rect 158902 6216 158958 6225
rect 158902 6151 158958 6160
rect 154396 4956 154448 4962
rect 154396 4898 154448 4904
rect 157800 4888 157852 4894
rect 157800 4830 157852 4836
rect 155408 3664 155460 3670
rect 155408 3606 155460 3612
rect 155420 480 155448 3606
rect 156602 3496 156658 3505
rect 156602 3431 156658 3440
rect 156616 480 156644 3431
rect 157812 480 157840 4830
rect 158916 480 158944 6151
rect 159836 4894 159864 76094
rect 159928 74534 159956 78503
rect 160020 78305 160048 79784
rect 160192 79766 160244 79772
rect 160284 79824 160336 79830
rect 160606 79824 160658 79830
rect 160284 79766 160336 79772
rect 160374 79792 160430 79801
rect 160006 78296 160062 78305
rect 160006 78231 160062 78240
rect 160204 76786 160232 79766
rect 160296 77246 160324 79766
rect 160802 79812 160830 80036
rect 160756 79801 160830 79812
rect 160742 79792 160830 79801
rect 160658 79772 160692 79778
rect 160606 79766 160692 79772
rect 160618 79750 160692 79766
rect 160374 79727 160430 79736
rect 160284 77240 160336 77246
rect 160284 77182 160336 77188
rect 160204 76758 160324 76786
rect 160192 76628 160244 76634
rect 160192 76570 160244 76576
rect 160098 76528 160154 76537
rect 160098 76463 160154 76472
rect 159928 74506 160048 74534
rect 160020 29714 160048 74506
rect 160008 29708 160060 29714
rect 160008 29650 160060 29656
rect 160112 14550 160140 76463
rect 160204 17338 160232 76570
rect 160296 17406 160324 76758
rect 160388 76634 160416 79727
rect 160468 79688 160520 79694
rect 160468 79630 160520 79636
rect 160480 76634 160508 79630
rect 160560 79620 160612 79626
rect 160560 79562 160612 79568
rect 160376 76628 160428 76634
rect 160376 76570 160428 76576
rect 160468 76628 160520 76634
rect 160468 76570 160520 76576
rect 160376 76356 160428 76362
rect 160376 76298 160428 76304
rect 160388 21486 160416 76298
rect 160468 76220 160520 76226
rect 160468 76162 160520 76168
rect 160480 22914 160508 76162
rect 160572 53310 160600 79562
rect 160664 78577 160692 79750
rect 160798 79784 160830 79792
rect 160894 79744 160922 80036
rect 160986 79830 161014 80036
rect 161078 79898 161106 80036
rect 161170 79966 161198 80036
rect 161158 79960 161210 79966
rect 161262 79937 161290 80036
rect 161158 79902 161210 79908
rect 161248 79928 161304 79937
rect 161066 79892 161118 79898
rect 161354 79898 161382 80036
rect 161248 79863 161304 79872
rect 161342 79892 161394 79898
rect 161066 79834 161118 79840
rect 161342 79834 161394 79840
rect 160974 79824 161026 79830
rect 160974 79766 161026 79772
rect 161204 79824 161256 79830
rect 161204 79766 161256 79772
rect 160742 79727 160798 79736
rect 160848 79716 160922 79744
rect 161112 79756 161164 79762
rect 160650 78568 160706 78577
rect 160650 78503 160706 78512
rect 160848 77330 160876 79716
rect 161112 79698 161164 79704
rect 161020 79688 161072 79694
rect 161020 79630 161072 79636
rect 160928 79620 160980 79626
rect 160928 79562 160980 79568
rect 160756 77302 160876 77330
rect 160652 76628 160704 76634
rect 160652 76570 160704 76576
rect 160664 54602 160692 76570
rect 160756 76362 160784 77302
rect 160836 77240 160888 77246
rect 160836 77182 160888 77188
rect 160744 76356 160796 76362
rect 160744 76298 160796 76304
rect 160744 76152 160796 76158
rect 160744 76094 160796 76100
rect 160756 60178 160784 76094
rect 160848 69834 160876 77182
rect 160940 76158 160968 79562
rect 161032 76226 161060 79630
rect 161124 76537 161152 79698
rect 161110 76528 161166 76537
rect 161110 76463 161166 76472
rect 161020 76220 161072 76226
rect 161020 76162 161072 76168
rect 160928 76152 160980 76158
rect 160928 76094 160980 76100
rect 161216 75449 161244 79766
rect 161446 79676 161474 80036
rect 161538 79744 161566 80036
rect 161630 79898 161658 80036
rect 161618 79892 161670 79898
rect 161618 79834 161670 79840
rect 161722 79744 161750 80036
rect 161538 79716 161612 79744
rect 161446 79648 161520 79676
rect 161388 79552 161440 79558
rect 161388 79494 161440 79500
rect 161296 78260 161348 78266
rect 161296 78202 161348 78208
rect 161202 75440 161258 75449
rect 161202 75375 161258 75384
rect 161308 70394 161336 78202
rect 161400 73154 161428 79494
rect 161492 76362 161520 79648
rect 161584 76786 161612 79716
rect 161676 79716 161750 79744
rect 161814 79744 161842 80036
rect 161906 79898 161934 80036
rect 161998 79937 162026 80036
rect 161984 79928 162040 79937
rect 161894 79892 161946 79898
rect 161984 79863 162040 79872
rect 161894 79834 161946 79840
rect 162090 79778 162118 80036
rect 162182 79898 162210 80036
rect 162170 79892 162222 79898
rect 162170 79834 162222 79840
rect 162274 79830 162302 80036
rect 162262 79824 162314 79830
rect 162090 79750 162164 79778
rect 162262 79766 162314 79772
rect 161814 79716 161888 79744
rect 161676 78470 161704 79716
rect 161664 78464 161716 78470
rect 161664 78406 161716 78412
rect 161584 76758 161796 76786
rect 161572 76628 161624 76634
rect 161572 76570 161624 76576
rect 161480 76356 161532 76362
rect 161480 76298 161532 76304
rect 161400 73126 161520 73154
rect 161124 70366 161336 70394
rect 160836 69828 160888 69834
rect 160836 69770 160888 69776
rect 161124 64874 161152 70366
rect 160940 64846 161152 64874
rect 160744 60172 160796 60178
rect 160744 60114 160796 60120
rect 160652 54596 160704 54602
rect 160652 54538 160704 54544
rect 160560 53304 160612 53310
rect 160560 53246 160612 53252
rect 160940 35290 160968 64846
rect 160928 35284 160980 35290
rect 160928 35226 160980 35232
rect 160468 22908 160520 22914
rect 160468 22850 160520 22856
rect 160376 21480 160428 21486
rect 160376 21422 160428 21428
rect 160284 17400 160336 17406
rect 160284 17342 160336 17348
rect 160192 17332 160244 17338
rect 160192 17274 160244 17280
rect 160100 14544 160152 14550
rect 160100 14486 160152 14492
rect 161492 6322 161520 73126
rect 161584 6390 161612 76570
rect 161664 76560 161716 76566
rect 161664 76502 161716 76508
rect 161572 6384 161624 6390
rect 161572 6326 161624 6332
rect 161480 6316 161532 6322
rect 161480 6258 161532 6264
rect 161676 6254 161704 76502
rect 161768 6526 161796 76758
rect 161756 6520 161808 6526
rect 161756 6462 161808 6468
rect 161860 6458 161888 79716
rect 161940 79688 161992 79694
rect 161940 79630 161992 79636
rect 162032 79688 162084 79694
rect 162136 79676 162164 79750
rect 162366 79676 162394 80036
rect 162458 79812 162486 80036
rect 162550 79966 162578 80036
rect 162538 79960 162590 79966
rect 162642 79937 162670 80036
rect 162538 79902 162590 79908
rect 162628 79928 162684 79937
rect 162734 79898 162762 80036
rect 162628 79863 162684 79872
rect 162722 79892 162774 79898
rect 162722 79834 162774 79840
rect 162584 79824 162636 79830
rect 162458 79784 162532 79812
rect 162136 79648 162256 79676
rect 162032 79630 162084 79636
rect 161952 9110 161980 79630
rect 161940 9104 161992 9110
rect 161940 9046 161992 9052
rect 162044 9042 162072 79630
rect 162124 79416 162176 79422
rect 162124 79358 162176 79364
rect 162136 78402 162164 79358
rect 162124 78396 162176 78402
rect 162124 78338 162176 78344
rect 162228 76634 162256 79648
rect 162320 79648 162394 79676
rect 162216 76628 162268 76634
rect 162216 76570 162268 76576
rect 162320 76566 162348 79648
rect 162308 76560 162360 76566
rect 162122 76528 162178 76537
rect 162504 76537 162532 79784
rect 162584 79766 162636 79772
rect 162308 76502 162360 76508
rect 162490 76528 162546 76537
rect 162122 76463 162178 76472
rect 162490 76463 162546 76472
rect 162136 68406 162164 76463
rect 162596 76401 162624 79766
rect 162676 79756 162728 79762
rect 162676 79698 162728 79704
rect 162688 77897 162716 79698
rect 162826 79676 162854 80036
rect 162918 79801 162946 80036
rect 163010 79937 163038 80036
rect 162996 79928 163052 79937
rect 163102 79898 163130 80036
rect 163194 79898 163222 80036
rect 163286 79966 163314 80036
rect 163274 79960 163326 79966
rect 163274 79902 163326 79908
rect 162996 79863 163052 79872
rect 163090 79892 163142 79898
rect 163090 79834 163142 79840
rect 163182 79892 163234 79898
rect 163182 79834 163234 79840
rect 162904 79792 162960 79801
rect 163378 79778 163406 80036
rect 162904 79727 162960 79736
rect 163044 79756 163096 79762
rect 163044 79698 163096 79704
rect 163136 79756 163188 79762
rect 163332 79750 163406 79778
rect 163188 79716 163268 79744
rect 163136 79698 163188 79704
rect 162780 79648 162854 79676
rect 162952 79688 163004 79694
rect 162780 78266 162808 79648
rect 162952 79630 163004 79636
rect 162860 79484 162912 79490
rect 162860 79426 162912 79432
rect 162768 78260 162820 78266
rect 162768 78202 162820 78208
rect 162768 77988 162820 77994
rect 162768 77930 162820 77936
rect 162674 77888 162730 77897
rect 162674 77823 162730 77832
rect 162582 76392 162638 76401
rect 162582 76327 162638 76336
rect 162124 68400 162176 68406
rect 162124 68342 162176 68348
rect 162780 64874 162808 77930
rect 162320 64846 162808 64874
rect 162320 61606 162348 64846
rect 162308 61600 162360 61606
rect 162308 61542 162360 61548
rect 162032 9036 162084 9042
rect 162032 8978 162084 8984
rect 161848 6452 161900 6458
rect 161848 6394 161900 6400
rect 161664 6248 161716 6254
rect 161664 6190 161716 6196
rect 159824 4888 159876 4894
rect 159824 4830 159876 4836
rect 162872 4826 162900 79426
rect 162964 13122 162992 79630
rect 163056 77246 163084 79698
rect 163136 79076 163188 79082
rect 163136 79018 163188 79024
rect 163148 78849 163176 79018
rect 163134 78840 163190 78849
rect 163134 78775 163190 78784
rect 163240 78305 163268 79716
rect 163226 78296 163282 78305
rect 163226 78231 163282 78240
rect 163044 77240 163096 77246
rect 163044 77182 163096 77188
rect 163044 76628 163096 76634
rect 163044 76570 163096 76576
rect 163056 14482 163084 76570
rect 163136 76016 163188 76022
rect 163136 75958 163188 75964
rect 163148 15910 163176 75958
rect 163228 75064 163280 75070
rect 163228 75006 163280 75012
rect 163240 35222 163268 75006
rect 163332 44878 163360 79750
rect 163470 79676 163498 80036
rect 163562 79830 163590 80036
rect 163550 79824 163602 79830
rect 163550 79766 163602 79772
rect 163654 79778 163682 80036
rect 163746 79898 163774 80036
rect 163838 79898 163866 80036
rect 163930 79966 163958 80036
rect 163918 79960 163970 79966
rect 164022 79937 164050 80036
rect 163918 79902 163970 79908
rect 164008 79928 164064 79937
rect 163734 79892 163786 79898
rect 163734 79834 163786 79840
rect 163826 79892 163878 79898
rect 164008 79863 164064 79872
rect 163826 79834 163878 79840
rect 164114 79801 164142 80036
rect 164206 79937 164234 80036
rect 164192 79928 164248 79937
rect 164192 79863 164248 79872
rect 164100 79792 164156 79801
rect 163654 79750 163820 79778
rect 163424 79648 163498 79676
rect 163424 54534 163452 79648
rect 163504 79552 163556 79558
rect 163504 79494 163556 79500
rect 163688 79552 163740 79558
rect 163688 79494 163740 79500
rect 163516 76634 163544 79494
rect 163596 77240 163648 77246
rect 163596 77182 163648 77188
rect 163504 76628 163556 76634
rect 163504 76570 163556 76576
rect 163502 76528 163558 76537
rect 163502 76463 163558 76472
rect 163516 60110 163544 76463
rect 163608 62830 163636 77182
rect 163700 75070 163728 79494
rect 163792 75342 163820 79750
rect 164298 79744 164326 80036
rect 164100 79727 164156 79736
rect 164252 79716 164326 79744
rect 164148 79688 164200 79694
rect 164148 79630 164200 79636
rect 163872 79620 163924 79626
rect 163872 79562 163924 79568
rect 164056 79620 164108 79626
rect 164056 79562 164108 79568
rect 163884 76022 163912 79562
rect 163964 79416 164016 79422
rect 163964 79358 164016 79364
rect 163976 77246 164004 79358
rect 163964 77240 164016 77246
rect 163964 77182 164016 77188
rect 163872 76016 163924 76022
rect 163872 75958 163924 75964
rect 163780 75336 163832 75342
rect 163780 75278 163832 75284
rect 163688 75064 163740 75070
rect 164068 75041 164096 79562
rect 164160 76294 164188 79630
rect 164252 79422 164280 79716
rect 164390 79676 164418 80036
rect 164482 79744 164510 80036
rect 164574 79966 164602 80036
rect 164562 79960 164614 79966
rect 164562 79902 164614 79908
rect 164666 79812 164694 80036
rect 164620 79784 164694 79812
rect 164482 79716 164556 79744
rect 164344 79648 164418 79676
rect 164240 79416 164292 79422
rect 164240 79358 164292 79364
rect 164240 78804 164292 78810
rect 164240 78746 164292 78752
rect 164148 76288 164200 76294
rect 164148 76230 164200 76236
rect 163688 75006 163740 75012
rect 164054 75032 164110 75041
rect 164054 74967 164110 74976
rect 163596 62824 163648 62830
rect 163596 62766 163648 62772
rect 163504 60104 163556 60110
rect 163504 60046 163556 60052
rect 163412 54528 163464 54534
rect 163412 54470 163464 54476
rect 163320 44872 163372 44878
rect 163320 44814 163372 44820
rect 163228 35216 163280 35222
rect 163228 35158 163280 35164
rect 163136 15904 163188 15910
rect 163136 15846 163188 15852
rect 163044 14476 163096 14482
rect 163044 14418 163096 14424
rect 162952 13116 163004 13122
rect 162952 13058 163004 13064
rect 164252 7614 164280 78746
rect 164344 76566 164372 79648
rect 164424 78124 164476 78130
rect 164424 78066 164476 78072
rect 164332 76560 164384 76566
rect 164332 76502 164384 76508
rect 164436 76378 164464 78066
rect 164344 76350 164464 76378
rect 164344 17270 164372 76350
rect 164424 76288 164476 76294
rect 164424 76230 164476 76236
rect 164436 18834 164464 76230
rect 164528 22846 164556 79716
rect 164620 47666 164648 79784
rect 164758 79744 164786 80036
rect 164850 79830 164878 80036
rect 164838 79824 164890 79830
rect 164838 79766 164890 79772
rect 164712 79716 164786 79744
rect 164942 79744 164970 80036
rect 165034 79898 165062 80036
rect 165022 79892 165074 79898
rect 165022 79834 165074 79840
rect 165126 79744 165154 80036
rect 165218 79966 165246 80036
rect 165206 79960 165258 79966
rect 165310 79937 165338 80036
rect 165206 79902 165258 79908
rect 165296 79928 165352 79937
rect 165296 79863 165352 79872
rect 165252 79824 165304 79830
rect 165252 79766 165304 79772
rect 164942 79716 165016 79744
rect 164712 78810 164740 79716
rect 164882 79656 164938 79665
rect 164792 79620 164844 79626
rect 164882 79591 164938 79600
rect 164792 79562 164844 79568
rect 164700 78804 164752 78810
rect 164700 78746 164752 78752
rect 164700 78600 164752 78606
rect 164700 78542 164752 78548
rect 164712 78198 164740 78542
rect 164700 78192 164752 78198
rect 164700 78134 164752 78140
rect 164804 76650 164832 79562
rect 164896 79490 164924 79591
rect 164884 79484 164936 79490
rect 164884 79426 164936 79432
rect 164884 79348 164936 79354
rect 164884 79290 164936 79296
rect 164896 78810 164924 79290
rect 164884 78804 164936 78810
rect 164884 78746 164936 78752
rect 164882 78432 164938 78441
rect 164882 78367 164938 78376
rect 164896 77790 164924 78367
rect 164988 78130 165016 79716
rect 165080 79716 165154 79744
rect 164976 78124 165028 78130
rect 164976 78066 165028 78072
rect 164974 78024 165030 78033
rect 164974 77959 165030 77968
rect 164884 77784 164936 77790
rect 164884 77726 164936 77732
rect 164988 77625 165016 77959
rect 164974 77616 165030 77625
rect 164884 77580 164936 77586
rect 164974 77551 165030 77560
rect 164884 77522 164936 77528
rect 164896 77314 164924 77522
rect 164884 77308 164936 77314
rect 164884 77250 164936 77256
rect 164882 77208 164938 77217
rect 164882 77143 164938 77152
rect 164712 76622 164832 76650
rect 164712 57322 164740 76622
rect 164792 76560 164844 76566
rect 164792 76502 164844 76508
rect 164804 60042 164832 76502
rect 164896 76265 164924 77143
rect 164882 76256 164938 76265
rect 164882 76191 164938 76200
rect 164884 75744 164936 75750
rect 164884 75686 164936 75692
rect 164896 75410 164924 75686
rect 164884 75404 164936 75410
rect 164884 75346 164936 75352
rect 165080 73154 165108 79716
rect 165158 79520 165214 79529
rect 165158 79455 165214 79464
rect 165172 79286 165200 79455
rect 165160 79280 165212 79286
rect 165160 79222 165212 79228
rect 165160 78736 165212 78742
rect 165160 78678 165212 78684
rect 165172 78402 165200 78678
rect 165160 78396 165212 78402
rect 165160 78338 165212 78344
rect 164896 73126 165108 73154
rect 164896 71126 164924 73126
rect 165264 71194 165292 79766
rect 165402 79744 165430 80036
rect 165494 79801 165522 80036
rect 165356 79716 165430 79744
rect 165480 79792 165536 79801
rect 165480 79727 165536 79736
rect 165586 79744 165614 80036
rect 165678 79898 165706 80036
rect 165770 79937 165798 80036
rect 165756 79928 165812 79937
rect 165666 79892 165718 79898
rect 165756 79863 165812 79872
rect 165666 79834 165718 79840
rect 165862 79744 165890 80036
rect 165954 79966 165982 80036
rect 165942 79960 165994 79966
rect 165942 79902 165994 79908
rect 166046 79744 166074 80036
rect 166138 79898 166166 80036
rect 166126 79892 166178 79898
rect 166126 79834 166178 79840
rect 166230 79744 166258 80036
rect 165586 79716 165660 79744
rect 165356 76537 165384 79716
rect 165528 79620 165580 79626
rect 165528 79562 165580 79568
rect 165540 79354 165568 79562
rect 165528 79348 165580 79354
rect 165528 79290 165580 79296
rect 165436 79280 165488 79286
rect 165436 79222 165488 79228
rect 165448 78946 165476 79222
rect 165436 78940 165488 78946
rect 165436 78882 165488 78888
rect 165528 78940 165580 78946
rect 165528 78882 165580 78888
rect 165434 78704 165490 78713
rect 165434 78639 165490 78648
rect 165448 78198 165476 78639
rect 165540 78334 165568 78882
rect 165528 78328 165580 78334
rect 165528 78270 165580 78276
rect 165436 78192 165488 78198
rect 165436 78134 165488 78140
rect 165342 76528 165398 76537
rect 165342 76463 165398 76472
rect 165632 76401 165660 79716
rect 165816 79716 165890 79744
rect 166000 79716 166074 79744
rect 166184 79716 166258 79744
rect 166322 79744 166350 80036
rect 166414 79966 166442 80036
rect 166402 79960 166454 79966
rect 166402 79902 166454 79908
rect 166506 79812 166534 80036
rect 166460 79784 166534 79812
rect 166322 79716 166396 79744
rect 165712 79620 165764 79626
rect 165712 79562 165764 79568
rect 165618 76392 165674 76401
rect 165618 76327 165674 76336
rect 165724 76242 165752 79562
rect 165816 79218 165844 79716
rect 165894 79656 165950 79665
rect 165894 79591 165950 79600
rect 165804 79212 165856 79218
rect 165804 79154 165856 79160
rect 165804 79076 165856 79082
rect 165804 79018 165856 79024
rect 165816 78334 165844 79018
rect 165804 78328 165856 78334
rect 165804 78270 165856 78276
rect 165804 76628 165856 76634
rect 165804 76570 165856 76576
rect 165632 76214 165752 76242
rect 165252 71188 165304 71194
rect 165252 71130 165304 71136
rect 164884 71120 164936 71126
rect 164884 71062 164936 71068
rect 165068 71052 165120 71058
rect 165068 70994 165120 71000
rect 164792 60036 164844 60042
rect 164792 59978 164844 59984
rect 164700 57316 164752 57322
rect 164700 57258 164752 57264
rect 164608 47660 164660 47666
rect 164608 47602 164660 47608
rect 164516 22840 164568 22846
rect 164516 22782 164568 22788
rect 164424 18828 164476 18834
rect 164424 18770 164476 18776
rect 164332 17264 164384 17270
rect 164332 17206 164384 17212
rect 164240 7608 164292 7614
rect 164240 7550 164292 7556
rect 162492 4820 162544 4826
rect 162492 4762 162544 4768
rect 162860 4820 162912 4826
rect 162860 4762 162912 4768
rect 160100 3596 160152 3602
rect 160100 3538 160152 3544
rect 160112 480 160140 3538
rect 161294 3360 161350 3369
rect 161294 3295 161350 3304
rect 161308 480 161336 3295
rect 162504 480 162532 4762
rect 163688 3528 163740 3534
rect 163688 3470 163740 3476
rect 163700 480 163728 3470
rect 164884 3460 164936 3466
rect 164884 3402 164936 3408
rect 164896 480 164924 3402
rect 165080 3126 165108 70994
rect 165632 8974 165660 76214
rect 165712 76152 165764 76158
rect 165712 76094 165764 76100
rect 165724 26926 165752 76094
rect 165816 50522 165844 76570
rect 165804 50516 165856 50522
rect 165804 50458 165856 50464
rect 165908 49026 165936 79591
rect 166000 50590 166028 79716
rect 166080 79076 166132 79082
rect 166080 79018 166132 79024
rect 166092 77654 166120 79018
rect 166080 77648 166132 77654
rect 166080 77590 166132 77596
rect 166184 71058 166212 79716
rect 166264 79620 166316 79626
rect 166264 79562 166316 79568
rect 166276 76158 166304 79562
rect 166368 76634 166396 79716
rect 166460 76634 166488 79784
rect 166598 79744 166626 80036
rect 166552 79716 166626 79744
rect 166690 79744 166718 80036
rect 166782 79937 166810 80036
rect 166768 79928 166824 79937
rect 166768 79863 166824 79872
rect 166874 79801 166902 80036
rect 166860 79792 166916 79801
rect 166690 79716 166764 79744
rect 166860 79727 166916 79736
rect 166966 79744 166994 80036
rect 167058 79898 167086 80036
rect 167046 79892 167098 79898
rect 167046 79834 167098 79840
rect 167150 79744 167178 80036
rect 166966 79716 167040 79744
rect 166356 76628 166408 76634
rect 166356 76570 166408 76576
rect 166448 76628 166500 76634
rect 166448 76570 166500 76576
rect 166264 76152 166316 76158
rect 166264 76094 166316 76100
rect 166172 71052 166224 71058
rect 166172 70994 166224 71000
rect 166552 70394 166580 79716
rect 166632 79552 166684 79558
rect 166632 79494 166684 79500
rect 166644 77314 166672 79494
rect 166632 77308 166684 77314
rect 166632 77250 166684 77256
rect 166632 76628 166684 76634
rect 166632 76570 166684 76576
rect 166644 72418 166672 76570
rect 166736 76537 166764 79716
rect 166816 79688 166868 79694
rect 166816 79630 166868 79636
rect 166828 77994 166856 79630
rect 166908 79416 166960 79422
rect 166908 79358 166960 79364
rect 166920 78606 166948 79358
rect 166908 78600 166960 78606
rect 166908 78542 166960 78548
rect 166816 77988 166868 77994
rect 166816 77930 166868 77936
rect 166816 77376 166868 77382
rect 166816 77318 166868 77324
rect 166722 76528 166778 76537
rect 166722 76463 166778 76472
rect 166632 72412 166684 72418
rect 166632 72354 166684 72360
rect 166828 70394 166856 77318
rect 167012 76401 167040 79716
rect 167104 79716 167178 79744
rect 167242 79744 167270 80036
rect 167334 79937 167362 80036
rect 167320 79928 167376 79937
rect 167320 79863 167376 79872
rect 167426 79744 167454 80036
rect 167518 79966 167546 80036
rect 167506 79960 167558 79966
rect 167506 79902 167558 79908
rect 167610 79812 167638 80036
rect 167702 79937 167730 80036
rect 167794 79966 167822 80036
rect 167782 79960 167834 79966
rect 167688 79928 167744 79937
rect 167782 79902 167834 79908
rect 167688 79863 167744 79872
rect 167610 79784 167776 79812
rect 167242 79716 167316 79744
rect 167426 79716 167592 79744
rect 166998 76392 167054 76401
rect 166998 76327 167054 76336
rect 167000 76288 167052 76294
rect 167000 76230 167052 76236
rect 166092 70366 166580 70394
rect 166644 70366 166856 70394
rect 167012 70394 167040 76230
rect 167104 75478 167132 79716
rect 167182 79656 167238 79665
rect 167182 79591 167238 79600
rect 167092 75472 167144 75478
rect 167092 75414 167144 75420
rect 167012 70366 167132 70394
rect 166092 51814 166120 70366
rect 166080 51808 166132 51814
rect 166080 51750 166132 51756
rect 166264 51740 166316 51746
rect 166264 51682 166316 51688
rect 165988 50584 166040 50590
rect 165988 50526 166040 50532
rect 165804 49020 165856 49026
rect 165804 48962 165856 48968
rect 165896 49020 165948 49026
rect 165896 48962 165948 48968
rect 165712 26920 165764 26926
rect 165712 26862 165764 26868
rect 165816 16574 165844 48962
rect 165816 16546 166120 16574
rect 165620 8968 165672 8974
rect 165620 8910 165672 8916
rect 165068 3120 165120 3126
rect 165068 3062 165120 3068
rect 166092 480 166120 16546
rect 166276 3398 166304 51682
rect 166644 36582 166672 70366
rect 166632 36576 166684 36582
rect 166632 36518 166684 36524
rect 167104 25566 167132 70366
rect 167196 25634 167224 79591
rect 167288 29646 167316 79716
rect 167368 79620 167420 79626
rect 167368 79562 167420 79568
rect 167380 31074 167408 79562
rect 167460 79348 167512 79354
rect 167460 79290 167512 79296
rect 167472 75614 167500 79290
rect 167460 75608 167512 75614
rect 167460 75550 167512 75556
rect 167460 75472 167512 75478
rect 167460 75414 167512 75420
rect 167472 51746 167500 75414
rect 167564 53242 167592 79716
rect 167642 78568 167698 78577
rect 167642 78503 167698 78512
rect 167656 78470 167684 78503
rect 167644 78464 167696 78470
rect 167644 78406 167696 78412
rect 167644 76628 167696 76634
rect 167644 76570 167696 76576
rect 167656 66910 167684 76570
rect 167748 66978 167776 79784
rect 167886 79744 167914 80036
rect 167840 79716 167914 79744
rect 167840 76634 167868 79716
rect 167978 79676 168006 80036
rect 168070 79801 168098 80036
rect 168056 79792 168112 79801
rect 168056 79727 168112 79736
rect 168162 79744 168190 80036
rect 168254 79937 168282 80036
rect 168346 79966 168374 80036
rect 168334 79960 168386 79966
rect 168240 79928 168296 79937
rect 168334 79902 168386 79908
rect 168438 79898 168466 80036
rect 168240 79863 168296 79872
rect 168426 79892 168478 79898
rect 168426 79834 168478 79840
rect 168288 79824 168340 79830
rect 168530 79778 168558 80036
rect 168288 79766 168340 79772
rect 168162 79716 168236 79744
rect 167932 79648 168006 79676
rect 168102 79656 168158 79665
rect 167828 76628 167880 76634
rect 167828 76570 167880 76576
rect 167826 76392 167882 76401
rect 167826 76327 167828 76336
rect 167880 76327 167882 76336
rect 167828 76298 167880 76304
rect 167932 76294 167960 79648
rect 168102 79591 168158 79600
rect 168012 79212 168064 79218
rect 168012 79154 168064 79160
rect 167920 76288 167972 76294
rect 167920 76230 167972 76236
rect 167828 75608 167880 75614
rect 167828 75550 167880 75556
rect 167840 75274 167868 75550
rect 167828 75268 167880 75274
rect 167828 75210 167880 75216
rect 168024 75206 168052 79154
rect 168012 75200 168064 75206
rect 168012 75142 168064 75148
rect 168116 70394 168144 79591
rect 168208 76537 168236 79716
rect 168194 76528 168250 76537
rect 168194 76463 168250 76472
rect 168300 73154 168328 79766
rect 168380 79756 168432 79762
rect 168380 79698 168432 79704
rect 168484 79750 168558 79778
rect 168392 78062 168420 79698
rect 168380 78056 168432 78062
rect 168380 77998 168432 78004
rect 168380 76560 168432 76566
rect 168380 76502 168432 76508
rect 167932 70366 168144 70394
rect 168208 73126 168328 73154
rect 167932 69766 167960 70366
rect 167920 69760 167972 69766
rect 167920 69702 167972 69708
rect 167736 66972 167788 66978
rect 167736 66914 167788 66920
rect 167644 66904 167696 66910
rect 167644 66846 167696 66852
rect 167552 53236 167604 53242
rect 167552 53178 167604 53184
rect 167460 51740 167512 51746
rect 167460 51682 167512 51688
rect 167368 31068 167420 31074
rect 167368 31010 167420 31016
rect 167276 29640 167328 29646
rect 167276 29582 167328 29588
rect 167184 25628 167236 25634
rect 167184 25570 167236 25576
rect 167092 25560 167144 25566
rect 167092 25502 167144 25508
rect 167184 11756 167236 11762
rect 167184 11698 167236 11704
rect 166264 3392 166316 3398
rect 166264 3334 166316 3340
rect 167196 480 167224 11698
rect 168208 10334 168236 73126
rect 168392 18630 168420 76502
rect 168484 76362 168512 79750
rect 168622 79676 168650 80036
rect 168714 79744 168742 80036
rect 168806 79937 168834 80036
rect 168898 79966 168926 80036
rect 168886 79960 168938 79966
rect 168792 79928 168848 79937
rect 168990 79937 169018 80036
rect 169082 79966 169110 80036
rect 169070 79960 169122 79966
rect 168886 79902 168938 79908
rect 168976 79928 169032 79937
rect 168792 79863 168848 79872
rect 169070 79902 169122 79908
rect 168976 79863 169032 79872
rect 169174 79812 169202 80036
rect 169266 79898 169294 80036
rect 169254 79892 169306 79898
rect 169254 79834 169306 79840
rect 169128 79784 169202 79812
rect 169024 79756 169076 79762
rect 168714 79716 168788 79744
rect 168576 79648 168650 79676
rect 168760 79665 168788 79716
rect 169024 79698 169076 79704
rect 168932 79688 168984 79694
rect 168746 79656 168802 79665
rect 168472 76356 168524 76362
rect 168472 76298 168524 76304
rect 168472 76220 168524 76226
rect 168472 76162 168524 76168
rect 168484 18698 168512 76162
rect 168576 18766 168604 79648
rect 168932 79630 168984 79636
rect 168746 79591 168802 79600
rect 168840 79620 168892 79626
rect 168840 79562 168892 79568
rect 168656 79416 168708 79422
rect 168656 79358 168708 79364
rect 168668 78577 168696 79358
rect 168852 79218 168880 79562
rect 168840 79212 168892 79218
rect 168840 79154 168892 79160
rect 168838 78704 168894 78713
rect 168838 78639 168894 78648
rect 168654 78568 168710 78577
rect 168654 78503 168710 78512
rect 168746 78432 168802 78441
rect 168746 78367 168802 78376
rect 168656 76628 168708 76634
rect 168656 76570 168708 76576
rect 168668 47598 168696 76570
rect 168656 47592 168708 47598
rect 168656 47534 168708 47540
rect 168656 44940 168708 44946
rect 168656 44882 168708 44888
rect 168564 18760 168616 18766
rect 168564 18702 168616 18708
rect 168472 18692 168524 18698
rect 168472 18634 168524 18640
rect 168380 18624 168432 18630
rect 168380 18566 168432 18572
rect 168196 10328 168248 10334
rect 168196 10270 168248 10276
rect 168668 6914 168696 44882
rect 168760 43450 168788 78367
rect 168852 77450 168880 78639
rect 168840 77444 168892 77450
rect 168840 77386 168892 77392
rect 168840 76356 168892 76362
rect 168840 76298 168892 76304
rect 168852 53174 168880 76298
rect 168944 57254 168972 79630
rect 169036 76226 169064 79698
rect 169128 76566 169156 79784
rect 169358 79778 169386 80036
rect 169450 79966 169478 80036
rect 169438 79960 169490 79966
rect 169438 79902 169490 79908
rect 169312 79750 169386 79778
rect 169208 79688 169260 79694
rect 169208 79630 169260 79636
rect 169312 79642 169340 79750
rect 169542 79744 169570 80036
rect 169496 79716 169570 79744
rect 169116 76560 169168 76566
rect 169116 76502 169168 76508
rect 169024 76220 169076 76226
rect 169024 76162 169076 76168
rect 169220 70394 169248 79630
rect 169312 79614 169432 79642
rect 169300 79416 169352 79422
rect 169300 79358 169352 79364
rect 169312 77654 169340 79358
rect 169300 77648 169352 77654
rect 169300 77590 169352 77596
rect 169300 77240 169352 77246
rect 169300 77182 169352 77188
rect 169312 76566 169340 77182
rect 169404 76634 169432 79614
rect 169392 76628 169444 76634
rect 169392 76570 169444 76576
rect 169300 76560 169352 76566
rect 169300 76502 169352 76508
rect 169036 70366 169248 70394
rect 169036 68338 169064 70366
rect 169496 69698 169524 79716
rect 169634 79676 169662 80036
rect 169726 79801 169754 80036
rect 169818 79830 169846 80036
rect 169806 79824 169858 79830
rect 169712 79792 169768 79801
rect 169806 79766 169858 79772
rect 169712 79727 169768 79736
rect 169760 79688 169812 79694
rect 169634 79648 169708 79676
rect 169576 79212 169628 79218
rect 169576 79154 169628 79160
rect 169588 75177 169616 79154
rect 169680 76537 169708 79648
rect 169760 79630 169812 79636
rect 169772 79336 169800 79630
rect 169910 79540 169938 80036
rect 170002 79694 170030 80036
rect 169990 79688 170042 79694
rect 170094 79676 170122 80036
rect 170186 79744 170214 80036
rect 170278 79937 170306 80036
rect 170264 79928 170320 79937
rect 170264 79863 170320 79872
rect 170370 79744 170398 80036
rect 170186 79716 170260 79744
rect 170094 79648 170168 79676
rect 169990 79630 170042 79636
rect 170036 79552 170088 79558
rect 169910 79512 169984 79540
rect 169772 79308 169892 79336
rect 169760 79212 169812 79218
rect 169760 79154 169812 79160
rect 169666 76528 169722 76537
rect 169666 76463 169722 76472
rect 169574 75168 169630 75177
rect 169574 75103 169630 75112
rect 169484 69692 169536 69698
rect 169484 69634 169536 69640
rect 169024 68332 169076 68338
rect 169024 68274 169076 68280
rect 168932 57248 168984 57254
rect 168932 57190 168984 57196
rect 168840 53168 168892 53174
rect 168840 53110 168892 53116
rect 168748 43444 168800 43450
rect 168748 43386 168800 43392
rect 168392 6886 168696 6914
rect 168392 480 168420 6886
rect 169772 6186 169800 79154
rect 169864 77353 169892 79308
rect 169850 77344 169906 77353
rect 169850 77279 169906 77288
rect 169850 75984 169906 75993
rect 169850 75919 169906 75928
rect 169864 11762 169892 75919
rect 169956 75914 169984 79512
rect 170036 79494 170088 79500
rect 170048 78656 170076 79494
rect 170140 79218 170168 79648
rect 170128 79212 170180 79218
rect 170128 79154 170180 79160
rect 170048 78628 170168 78656
rect 169956 75886 170076 75914
rect 169944 75132 169996 75138
rect 169944 75074 169996 75080
rect 169956 33794 169984 75074
rect 170048 50386 170076 75886
rect 170140 53106 170168 78628
rect 170232 75138 170260 79716
rect 170324 79716 170398 79744
rect 170324 79506 170352 79716
rect 170462 79676 170490 80036
rect 170554 79744 170582 80036
rect 170646 79966 170674 80036
rect 170634 79960 170686 79966
rect 170634 79902 170686 79908
rect 170738 79898 170766 80036
rect 170726 79892 170778 79898
rect 170726 79834 170778 79840
rect 170830 79801 170858 80036
rect 170922 79971 170950 80036
rect 170908 79962 170964 79971
rect 170908 79897 170964 79906
rect 171014 79812 171042 80036
rect 171106 79966 171134 80036
rect 171198 79971 171226 80036
rect 171094 79960 171146 79966
rect 171094 79902 171146 79908
rect 171184 79962 171240 79971
rect 171184 79897 171240 79906
rect 170816 79792 170872 79801
rect 170554 79716 170628 79744
rect 171014 79784 171088 79812
rect 170816 79727 170872 79736
rect 170462 79648 170536 79676
rect 170324 79478 170444 79506
rect 170312 79416 170364 79422
rect 170312 79358 170364 79364
rect 170324 78713 170352 79358
rect 170310 78704 170366 78713
rect 170310 78639 170366 78648
rect 170312 77648 170364 77654
rect 170312 77590 170364 77596
rect 170324 76566 170352 77590
rect 170312 76560 170364 76566
rect 170312 76502 170364 76508
rect 170416 75993 170444 79478
rect 170508 77489 170536 79648
rect 170494 77480 170550 77489
rect 170494 77415 170550 77424
rect 170496 77308 170548 77314
rect 170496 77250 170548 77256
rect 170402 75984 170458 75993
rect 170402 75919 170458 75928
rect 170220 75132 170272 75138
rect 170220 75074 170272 75080
rect 170508 70394 170536 77250
rect 170600 76129 170628 79716
rect 170864 79688 170916 79694
rect 170864 79630 170916 79636
rect 170772 79620 170824 79626
rect 170772 79562 170824 79568
rect 170678 78976 170734 78985
rect 170678 78911 170734 78920
rect 170692 78713 170720 78911
rect 170678 78704 170734 78713
rect 170678 78639 170734 78648
rect 170784 78146 170812 79562
rect 170876 78538 170904 79630
rect 170956 79144 171008 79150
rect 170956 79086 171008 79092
rect 170968 78985 170996 79086
rect 170954 78976 171010 78985
rect 170954 78911 171010 78920
rect 170956 78736 171008 78742
rect 170956 78678 171008 78684
rect 170968 78538 170996 78678
rect 170864 78532 170916 78538
rect 170864 78474 170916 78480
rect 170956 78532 171008 78538
rect 170956 78474 171008 78480
rect 170784 78118 170904 78146
rect 170876 78062 170904 78118
rect 170772 78056 170824 78062
rect 170772 77998 170824 78004
rect 170864 78056 170916 78062
rect 170864 77998 170916 78004
rect 170586 76120 170642 76129
rect 170586 76055 170642 76064
rect 170508 70366 170628 70394
rect 170600 64874 170628 70366
rect 170508 64846 170628 64874
rect 170128 53100 170180 53106
rect 170128 53042 170180 53048
rect 170036 50380 170088 50386
rect 170036 50322 170088 50328
rect 169944 33788 169996 33794
rect 169944 33730 169996 33736
rect 170508 21418 170536 64846
rect 170784 50454 170812 77998
rect 170954 77888 171010 77897
rect 170954 77823 171010 77832
rect 170968 75954 170996 77823
rect 170956 75948 171008 75954
rect 170956 75890 171008 75896
rect 171060 73166 171088 79784
rect 171290 79642 171318 80036
rect 171382 79812 171410 80036
rect 171474 79971 171502 80036
rect 171460 79962 171516 79971
rect 171566 79966 171594 80036
rect 171460 79897 171516 79906
rect 171554 79960 171606 79966
rect 171554 79902 171606 79908
rect 171658 79898 171686 80036
rect 171750 79971 171778 80036
rect 171736 79962 171792 79971
rect 171842 79966 171870 80036
rect 171934 79966 171962 80036
rect 172026 79971 172054 80036
rect 171646 79892 171698 79898
rect 171736 79897 171792 79906
rect 171830 79960 171882 79966
rect 171830 79902 171882 79908
rect 171922 79960 171974 79966
rect 171922 79902 171974 79908
rect 172012 79962 172068 79971
rect 172118 79966 172146 80036
rect 172210 79966 172238 80036
rect 172012 79897 172068 79906
rect 172106 79960 172158 79966
rect 172106 79902 172158 79908
rect 172198 79960 172250 79966
rect 172198 79902 172250 79908
rect 171646 79834 171698 79840
rect 172060 79824 172112 79830
rect 171382 79784 171456 79812
rect 171244 79614 171318 79642
rect 171244 78742 171272 79614
rect 171324 79144 171376 79150
rect 171324 79086 171376 79092
rect 171232 78736 171284 78742
rect 171232 78678 171284 78684
rect 171140 78532 171192 78538
rect 171140 78474 171192 78480
rect 171152 75478 171180 78474
rect 171336 78441 171364 79086
rect 171428 78985 171456 79784
rect 172060 79766 172112 79772
rect 172152 79824 172204 79830
rect 172152 79766 172204 79772
rect 171600 79756 171652 79762
rect 171600 79698 171652 79704
rect 171508 79416 171560 79422
rect 171508 79358 171560 79364
rect 171414 78976 171470 78985
rect 171414 78911 171470 78920
rect 171520 78441 171548 79358
rect 171612 79286 171640 79698
rect 171968 79688 172020 79694
rect 171968 79630 172020 79636
rect 171704 79580 171916 79608
rect 171704 79490 171732 79580
rect 171692 79484 171744 79490
rect 171692 79426 171744 79432
rect 171784 79484 171836 79490
rect 171784 79426 171836 79432
rect 171692 79348 171744 79354
rect 171692 79290 171744 79296
rect 171600 79280 171652 79286
rect 171600 79222 171652 79228
rect 171704 79218 171732 79290
rect 171692 79212 171744 79218
rect 171692 79154 171744 79160
rect 171796 78713 171824 79426
rect 171888 79218 171916 79580
rect 171876 79212 171928 79218
rect 171876 79154 171928 79160
rect 171874 78840 171930 78849
rect 171874 78775 171930 78784
rect 171782 78704 171838 78713
rect 171782 78639 171838 78648
rect 171692 78600 171744 78606
rect 171692 78542 171744 78548
rect 171888 78554 171916 78775
rect 171980 78674 172008 79630
rect 171968 78668 172020 78674
rect 171968 78610 172020 78616
rect 171322 78432 171378 78441
rect 171322 78367 171378 78376
rect 171506 78432 171562 78441
rect 171506 78367 171562 78376
rect 171598 78296 171654 78305
rect 171598 78231 171654 78240
rect 171230 78160 171286 78169
rect 171230 78095 171286 78104
rect 171508 78124 171560 78130
rect 171244 77897 171272 78095
rect 171508 78066 171560 78072
rect 171324 77920 171376 77926
rect 171230 77888 171286 77897
rect 171324 77862 171376 77868
rect 171230 77823 171286 77832
rect 171230 77752 171286 77761
rect 171230 77687 171286 77696
rect 171140 75472 171192 75478
rect 171140 75414 171192 75420
rect 171244 74526 171272 77687
rect 171232 74520 171284 74526
rect 171232 74462 171284 74468
rect 171048 73160 171100 73166
rect 171048 73102 171100 73108
rect 171336 70394 171364 77862
rect 171520 76362 171548 78066
rect 171612 77897 171640 78231
rect 171704 78130 171732 78542
rect 171888 78526 172008 78554
rect 171692 78124 171744 78130
rect 171692 78066 171744 78072
rect 171980 77994 172008 78526
rect 172072 78305 172100 79766
rect 172058 78296 172114 78305
rect 172058 78231 172114 78240
rect 171876 77988 171928 77994
rect 171876 77930 171928 77936
rect 171968 77988 172020 77994
rect 171968 77930 172020 77936
rect 171598 77888 171654 77897
rect 171598 77823 171654 77832
rect 171784 77852 171836 77858
rect 171784 77794 171836 77800
rect 171692 77716 171744 77722
rect 171692 77658 171744 77664
rect 171600 77444 171652 77450
rect 171600 77386 171652 77392
rect 171508 76356 171560 76362
rect 171508 76298 171560 76304
rect 171612 76242 171640 77386
rect 171520 76214 171640 76242
rect 171336 70366 171456 70394
rect 170772 50448 170824 50454
rect 170772 50390 170824 50396
rect 171428 28286 171456 70366
rect 171416 28280 171468 28286
rect 171416 28222 171468 28228
rect 171520 27062 171548 76214
rect 171704 74610 171732 77658
rect 171796 77450 171824 77794
rect 171784 77444 171836 77450
rect 171784 77386 171836 77392
rect 171784 76628 171836 76634
rect 171784 76570 171836 76576
rect 171612 74582 171732 74610
rect 171612 49094 171640 74582
rect 171692 74520 171744 74526
rect 171692 74462 171744 74468
rect 171600 49088 171652 49094
rect 171600 49030 171652 49036
rect 171704 44946 171732 74462
rect 171692 44940 171744 44946
rect 171692 44882 171744 44888
rect 171508 27056 171560 27062
rect 171508 26998 171560 27004
rect 170496 21412 170548 21418
rect 170496 21354 170548 21360
rect 169852 11756 169904 11762
rect 169852 11698 169904 11704
rect 169760 6180 169812 6186
rect 169760 6122 169812 6128
rect 169576 5160 169628 5166
rect 169576 5102 169628 5108
rect 169588 480 169616 5102
rect 171796 3670 171824 76570
rect 171784 3664 171836 3670
rect 171784 3606 171836 3612
rect 170772 3392 170824 3398
rect 170772 3334 170824 3340
rect 170784 480 170812 3334
rect 171888 3262 171916 77930
rect 172164 77790 172192 79766
rect 172302 79744 172330 80036
rect 172394 79971 172422 80036
rect 172380 79962 172436 79971
rect 172380 79897 172436 79906
rect 172486 79744 172514 80036
rect 172578 79966 172606 80036
rect 172566 79960 172618 79966
rect 172566 79902 172618 79908
rect 172670 79812 172698 80036
rect 172624 79784 172698 79812
rect 172302 79716 172376 79744
rect 172486 79716 172560 79744
rect 172152 77784 172204 77790
rect 172152 77726 172204 77732
rect 172242 77752 172298 77761
rect 172242 77687 172298 77696
rect 172058 77616 172114 77625
rect 172058 77551 172114 77560
rect 171966 75848 172022 75857
rect 171966 75783 172022 75792
rect 171980 3534 172008 75783
rect 172072 23050 172100 77551
rect 172150 77208 172206 77217
rect 172150 77143 172206 77152
rect 172164 76634 172192 77143
rect 172152 76628 172204 76634
rect 172152 76570 172204 76576
rect 172150 75032 172206 75041
rect 172150 74967 172206 74976
rect 172060 23044 172112 23050
rect 172060 22986 172112 22992
rect 172164 3602 172192 74967
rect 172256 7682 172284 77687
rect 172348 77246 172376 79716
rect 172426 78976 172482 78985
rect 172426 78911 172482 78920
rect 172440 78742 172468 78911
rect 172532 78849 172560 79716
rect 172624 79626 172652 79784
rect 172762 79744 172790 80036
rect 172716 79716 172790 79744
rect 172854 79744 172882 80036
rect 172946 79898 172974 80036
rect 172934 79892 172986 79898
rect 172934 79834 172986 79840
rect 173038 79778 173066 80036
rect 172992 79750 173066 79778
rect 173130 79778 173158 80036
rect 173222 79971 173250 80036
rect 173208 79962 173264 79971
rect 173208 79897 173264 79906
rect 173314 79898 173342 80036
rect 173302 79892 173354 79898
rect 173302 79834 173354 79840
rect 173130 79750 173204 79778
rect 172854 79716 172928 79744
rect 172612 79620 172664 79626
rect 172612 79562 172664 79568
rect 172716 79472 172744 79716
rect 172624 79444 172744 79472
rect 172518 78840 172574 78849
rect 172518 78775 172574 78784
rect 172624 78742 172652 79444
rect 172428 78736 172480 78742
rect 172428 78678 172480 78684
rect 172612 78736 172664 78742
rect 172612 78678 172664 78684
rect 172900 78538 172928 79716
rect 172992 79393 173020 79750
rect 173072 79688 173124 79694
rect 173072 79630 173124 79636
rect 172978 79384 173034 79393
rect 172978 79319 173034 79328
rect 173084 79257 173112 79630
rect 173176 79490 173204 79750
rect 173256 79756 173308 79762
rect 173406 79744 173434 80036
rect 173498 79812 173526 80036
rect 173590 79937 173618 80036
rect 173682 79966 173710 80036
rect 173670 79960 173722 79966
rect 173576 79928 173632 79937
rect 173670 79902 173722 79908
rect 173576 79863 173632 79872
rect 173624 79824 173676 79830
rect 173498 79784 173572 79812
rect 173256 79698 173308 79704
rect 173360 79716 173434 79744
rect 173268 79529 173296 79698
rect 173360 79665 173388 79716
rect 173346 79656 173402 79665
rect 173346 79591 173402 79600
rect 173254 79520 173310 79529
rect 173164 79484 173216 79490
rect 173254 79455 173310 79464
rect 173164 79426 173216 79432
rect 173348 79416 173400 79422
rect 173346 79384 173348 79393
rect 173400 79384 173402 79393
rect 173346 79319 173402 79328
rect 173070 79248 173126 79257
rect 173070 79183 173126 79192
rect 173544 78606 173572 79784
rect 173774 79812 173802 80036
rect 173624 79766 173676 79772
rect 173728 79784 173802 79812
rect 173636 79529 173664 79766
rect 173622 79520 173678 79529
rect 173728 79490 173756 79784
rect 173866 79744 173894 80036
rect 173958 79898 173986 80036
rect 174050 79937 174078 80036
rect 174036 79928 174092 79937
rect 173946 79892 173998 79898
rect 174036 79863 174092 79872
rect 173946 79834 173998 79840
rect 174142 79830 174170 80036
rect 174130 79824 174182 79830
rect 174130 79766 174182 79772
rect 173820 79716 173894 79744
rect 173992 79756 174044 79762
rect 173622 79455 173678 79464
rect 173716 79484 173768 79490
rect 173716 79426 173768 79432
rect 173820 79354 173848 79716
rect 173992 79698 174044 79704
rect 173898 79656 173954 79665
rect 173898 79591 173954 79600
rect 173808 79348 173860 79354
rect 173808 79290 173860 79296
rect 173912 78810 173940 79591
rect 173900 78804 173952 78810
rect 173900 78746 173952 78752
rect 173532 78600 173584 78606
rect 173532 78542 173584 78548
rect 172888 78532 172940 78538
rect 172888 78474 172940 78480
rect 174004 77518 174032 79698
rect 174084 79688 174136 79694
rect 174234 79642 174262 80036
rect 174326 79914 174354 80036
rect 174326 79886 174400 79914
rect 174084 79630 174136 79636
rect 174096 77994 174124 79630
rect 174188 79614 174262 79642
rect 174084 77988 174136 77994
rect 174084 77930 174136 77936
rect 173992 77512 174044 77518
rect 173992 77454 174044 77460
rect 172336 77240 172388 77246
rect 172336 77182 172388 77188
rect 173162 76392 173218 76401
rect 173162 76327 173218 76336
rect 172518 67008 172574 67017
rect 172518 66943 172574 66952
rect 172532 16574 172560 66943
rect 172532 16546 172744 16574
rect 172244 7676 172296 7682
rect 172244 7618 172296 7624
rect 172152 3596 172204 3602
rect 172152 3538 172204 3544
rect 171968 3528 172020 3534
rect 171968 3470 172020 3476
rect 171876 3256 171928 3262
rect 171876 3198 171928 3204
rect 171968 3120 172020 3126
rect 171968 3062 172020 3068
rect 171980 480 172008 3062
rect 148294 354 148406 480
rect 148060 326 148406 354
rect 148294 -960 148406 326
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 172716 354 172744 16546
rect 173176 3738 173204 76327
rect 173348 75948 173400 75954
rect 173348 75890 173400 75896
rect 173256 72412 173308 72418
rect 173256 72354 173308 72360
rect 173164 3732 173216 3738
rect 173164 3674 173216 3680
rect 173268 3466 173296 72354
rect 173360 33114 173388 75890
rect 174188 70394 174216 79614
rect 174372 70394 174400 79886
rect 174464 77586 174492 80174
rect 174544 79688 174596 79694
rect 174544 79630 174596 79636
rect 174556 79393 174584 79630
rect 174648 79490 174676 80582
rect 175740 80572 175792 80578
rect 175740 80514 175792 80520
rect 175752 80170 175780 80514
rect 175924 80504 175976 80510
rect 175924 80446 175976 80452
rect 175740 80164 175792 80170
rect 175740 80106 175792 80112
rect 175832 80164 175884 80170
rect 175832 80106 175884 80112
rect 175096 80096 175148 80102
rect 175096 80038 175148 80044
rect 175108 79490 175136 80038
rect 174636 79484 174688 79490
rect 174636 79426 174688 79432
rect 175096 79484 175148 79490
rect 175096 79426 175148 79432
rect 174542 79384 174598 79393
rect 174542 79319 174598 79328
rect 175844 79218 175872 80106
rect 175936 80102 175964 80446
rect 178052 80209 178080 80582
rect 178038 80200 178094 80209
rect 178038 80135 178094 80144
rect 175924 80096 175976 80102
rect 175924 80038 175976 80044
rect 177396 79552 177448 79558
rect 177394 79520 177396 79529
rect 177448 79520 177450 79529
rect 177394 79455 177450 79464
rect 175832 79212 175884 79218
rect 175832 79154 175884 79160
rect 178604 78985 178632 80650
rect 179512 79620 179564 79626
rect 179512 79562 179564 79568
rect 179524 78985 179552 79562
rect 178590 78976 178646 78985
rect 178590 78911 178646 78920
rect 179510 78976 179566 78985
rect 179510 78911 179566 78920
rect 174542 78432 174598 78441
rect 174542 78367 174598 78376
rect 174556 78062 174584 78367
rect 179142 78160 179198 78169
rect 179142 78095 179198 78104
rect 174544 78056 174596 78062
rect 174544 77998 174596 78004
rect 179156 77654 179184 78095
rect 179144 77648 179196 77654
rect 179144 77590 179196 77596
rect 174452 77580 174504 77586
rect 174452 77522 174504 77528
rect 178040 76424 178092 76430
rect 178040 76366 178092 76372
rect 175922 76256 175978 76265
rect 175922 76191 175978 76200
rect 174542 74352 174598 74361
rect 174542 74287 174598 74296
rect 174004 70366 174216 70394
rect 174280 70366 174400 70394
rect 174004 45558 174032 70366
rect 174280 64874 174308 70366
rect 174096 64846 174308 64874
rect 173992 45552 174044 45558
rect 173992 45494 174044 45500
rect 173348 33108 173400 33114
rect 173348 33050 173400 33056
rect 174096 23118 174124 64846
rect 174084 23112 174136 23118
rect 174084 23054 174136 23060
rect 174268 3528 174320 3534
rect 174268 3470 174320 3476
rect 173256 3460 173308 3466
rect 173256 3402 173308 3408
rect 174280 480 174308 3470
rect 174556 3330 174584 74287
rect 175278 69592 175334 69601
rect 175278 69527 175334 69536
rect 175292 16574 175320 69527
rect 175292 16546 175504 16574
rect 174544 3324 174596 3330
rect 174544 3266 174596 3272
rect 175476 480 175504 16546
rect 175936 3398 175964 76191
rect 176658 75712 176714 75721
rect 176658 75647 176714 75656
rect 176672 3534 176700 75647
rect 178052 16574 178080 76366
rect 179420 57588 179472 57594
rect 179420 57530 179472 57536
rect 179432 16574 179460 57530
rect 179892 24138 179920 130455
rect 180076 80345 180104 271866
rect 180156 229152 180208 229158
rect 180156 229094 180208 229100
rect 180168 202162 180196 229094
rect 180156 202156 180208 202162
rect 180156 202098 180208 202104
rect 180156 111852 180208 111858
rect 180156 111794 180208 111800
rect 180168 80442 180196 111794
rect 180156 80436 180208 80442
rect 180156 80378 180208 80384
rect 180062 80336 180118 80345
rect 180062 80271 180118 80280
rect 180812 78538 180840 700266
rect 182364 536852 182416 536858
rect 182364 536794 182416 536800
rect 180892 514820 180944 514826
rect 180892 514762 180944 514768
rect 180904 117473 180932 514762
rect 182272 484424 182324 484430
rect 182272 484366 182324 484372
rect 180984 357468 181036 357474
rect 180984 357410 181036 357416
rect 180996 121553 181024 357410
rect 182180 233844 182232 233850
rect 182180 233786 182232 233792
rect 182192 224262 182220 233786
rect 182180 224256 182232 224262
rect 182180 224198 182232 224204
rect 181076 196716 181128 196722
rect 181076 196658 181128 196664
rect 180982 121544 181038 121553
rect 180982 121479 181038 121488
rect 180890 117464 180946 117473
rect 180890 117399 180946 117408
rect 181088 109313 181116 196658
rect 181260 151088 181312 151094
rect 181260 151030 181312 151036
rect 181168 149116 181220 149122
rect 181168 149058 181220 149064
rect 181180 126993 181208 149058
rect 181166 126984 181222 126993
rect 181166 126919 181222 126928
rect 181272 114753 181300 151030
rect 181352 148368 181404 148374
rect 181352 148310 181404 148316
rect 181258 114744 181314 114753
rect 181258 114679 181314 114688
rect 181364 113393 181392 148310
rect 181444 140208 181496 140214
rect 181444 140150 181496 140156
rect 181456 120193 181484 140150
rect 182180 139392 182232 139398
rect 182180 139334 182232 139340
rect 181534 129704 181590 129713
rect 181534 129639 181590 129648
rect 181442 120184 181498 120193
rect 181442 120119 181498 120128
rect 181350 113384 181406 113393
rect 181350 113319 181406 113328
rect 181074 109304 181130 109313
rect 181074 109239 181130 109248
rect 180800 78532 180852 78538
rect 180800 78474 180852 78480
rect 180800 60376 180852 60382
rect 180800 60318 180852 60324
rect 179880 24132 179932 24138
rect 179880 24074 179932 24080
rect 180812 16574 180840 60318
rect 181548 59362 181576 129639
rect 182192 124273 182220 139334
rect 182178 124264 182234 124273
rect 182178 124199 182234 124208
rect 182180 99340 182232 99346
rect 182180 99282 182232 99288
rect 182192 98433 182220 99282
rect 182178 98424 182234 98433
rect 182178 98359 182234 98368
rect 182180 97436 182232 97442
rect 182180 97378 182232 97384
rect 182192 97073 182220 97378
rect 182178 97064 182234 97073
rect 182178 96999 182234 97008
rect 182284 78674 182312 484366
rect 182272 78668 182324 78674
rect 182272 78610 182324 78616
rect 182376 78305 182404 536794
rect 182560 233850 182588 700334
rect 185584 700324 185636 700330
rect 185584 700266 185636 700272
rect 184204 683188 184256 683194
rect 184204 683130 184256 683136
rect 182824 418192 182876 418198
rect 182824 418134 182876 418140
rect 182548 233844 182600 233850
rect 182548 233786 182600 233792
rect 182836 231606 182864 418134
rect 182824 231600 182876 231606
rect 182824 231542 182876 231548
rect 182560 229158 182588 230588
rect 182824 230376 182876 230382
rect 182824 230318 182876 230324
rect 182548 229152 182600 229158
rect 182548 229094 182600 229100
rect 182548 224256 182600 224262
rect 182548 224198 182600 224204
rect 182456 139324 182508 139330
rect 182456 139266 182508 139272
rect 182468 122913 182496 139266
rect 182454 122904 182510 122913
rect 182454 122839 182510 122848
rect 182560 110673 182588 224198
rect 182546 110664 182602 110673
rect 182546 110599 182602 110608
rect 182640 101312 182692 101318
rect 182640 101254 182692 101260
rect 182652 101153 182680 101254
rect 182638 101144 182694 101153
rect 182638 101079 182694 101088
rect 182456 100496 182508 100502
rect 182456 100438 182508 100444
rect 182468 99793 182496 100438
rect 182454 99784 182510 99793
rect 182454 99719 182510 99728
rect 182836 92993 182864 230318
rect 182916 151836 182968 151842
rect 182916 151778 182968 151784
rect 182822 92984 182878 92993
rect 182822 92919 182878 92928
rect 182822 80744 182878 80753
rect 182822 80679 182878 80688
rect 182362 78296 182418 78305
rect 182362 78231 182418 78240
rect 182180 76492 182232 76498
rect 182180 76434 182232 76440
rect 181536 59356 181588 59362
rect 181536 59298 181588 59304
rect 178052 16546 178632 16574
rect 179432 16546 180288 16574
rect 180812 16546 181024 16574
rect 176750 3904 176806 3913
rect 176750 3839 176806 3848
rect 176660 3528 176712 3534
rect 176660 3470 176712 3476
rect 175924 3392 175976 3398
rect 175924 3334 175976 3340
rect 176764 1986 176792 3839
rect 177856 3528 177908 3534
rect 177856 3470 177908 3476
rect 177948 3528 178000 3534
rect 177948 3470 178000 3476
rect 176672 1958 176792 1986
rect 176672 480 176700 1958
rect 177868 480 177896 3470
rect 177960 3262 177988 3470
rect 177948 3256 178000 3262
rect 177948 3198 178000 3204
rect 173134 354 173246 480
rect 172716 326 173246 354
rect 173134 -960 173246 326
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 178604 354 178632 16546
rect 180260 480 180288 16546
rect 179022 354 179134 480
rect 178604 326 179134 354
rect 179022 -960 179134 326
rect 180218 -960 180330 480
rect 180996 354 181024 16546
rect 181414 354 181526 480
rect 180996 326 181526 354
rect 182192 354 182220 76434
rect 182836 24138 182864 80679
rect 182928 79150 182956 151778
rect 183284 108996 183336 109002
rect 183284 108938 183336 108944
rect 183296 107953 183324 108938
rect 183282 107944 183338 107953
rect 183282 107879 183338 107888
rect 183284 107636 183336 107642
rect 183284 107578 183336 107584
rect 183296 106593 183324 107578
rect 183282 106584 183338 106593
rect 183282 106519 183338 106528
rect 183284 106276 183336 106282
rect 183284 106218 183336 106224
rect 183296 105233 183324 106218
rect 183282 105224 183338 105233
rect 183282 105159 183338 105168
rect 183284 104644 183336 104650
rect 183284 104586 183336 104592
rect 183296 103873 183324 104586
rect 183282 103864 183338 103873
rect 183282 103799 183338 103808
rect 183468 102944 183520 102950
rect 183468 102886 183520 102892
rect 183480 102513 183508 102886
rect 183466 102504 183522 102513
rect 183466 102439 183522 102448
rect 184216 100502 184244 683130
rect 184296 630692 184348 630698
rect 184296 630634 184348 630640
rect 184204 100496 184256 100502
rect 184204 100438 184256 100444
rect 184308 99346 184336 630634
rect 184388 576904 184440 576910
rect 184388 576846 184440 576852
rect 184296 99340 184348 99346
rect 184296 99282 184348 99288
rect 184400 97442 184428 576846
rect 185596 101318 185624 700266
rect 188356 102950 188384 700334
rect 189736 104650 189764 700402
rect 192496 106282 192524 700470
rect 193876 107642 193904 700538
rect 193956 138032 194008 138038
rect 193956 137974 194008 137980
rect 193864 107636 193916 107642
rect 193864 107578 193916 107584
rect 192484 106276 192536 106282
rect 192484 106218 192536 106224
rect 189724 104644 189776 104650
rect 189724 104586 189776 104592
rect 188344 102944 188396 102950
rect 188344 102886 188396 102892
rect 185584 101312 185636 101318
rect 185584 101254 185636 101260
rect 192484 99408 192536 99414
rect 192484 99350 192536 99356
rect 184388 97436 184440 97442
rect 184388 97378 184440 97384
rect 183192 96620 183244 96626
rect 183192 96562 183244 96568
rect 183204 95713 183232 96562
rect 183190 95704 183246 95713
rect 183190 95639 183246 95648
rect 183468 95192 183520 95198
rect 183468 95134 183520 95140
rect 183480 94353 183508 95134
rect 183466 94344 183522 94353
rect 183466 94279 183522 94288
rect 183376 93152 183428 93158
rect 183376 93094 183428 93100
rect 183388 91633 183416 93094
rect 183468 91792 183520 91798
rect 183468 91734 183520 91740
rect 183374 91624 183430 91633
rect 183374 91559 183430 91568
rect 183376 90364 183428 90370
rect 183376 90306 183428 90312
rect 183388 88913 183416 90306
rect 183480 90273 183508 91734
rect 183466 90264 183522 90273
rect 183466 90199 183522 90208
rect 183468 89004 183520 89010
rect 183468 88946 183520 88952
rect 183374 88904 183430 88913
rect 183374 88839 183430 88848
rect 183376 87644 183428 87650
rect 183376 87586 183428 87592
rect 183388 86193 183416 87586
rect 183480 87553 183508 88946
rect 183466 87544 183522 87553
rect 183466 87479 183522 87488
rect 183374 86184 183430 86193
rect 183374 86119 183430 86128
rect 183468 85536 183520 85542
rect 183468 85478 183520 85484
rect 183480 84833 183508 85478
rect 183466 84824 183522 84833
rect 183466 84759 183522 84768
rect 192496 84182 192524 99350
rect 193968 85542 193996 137974
rect 196636 109002 196664 700606
rect 196624 108996 196676 109002
rect 196624 108938 196676 108944
rect 193956 85536 194008 85542
rect 193956 85478 194008 85484
rect 183468 84176 183520 84182
rect 183468 84118 183520 84124
rect 192484 84176 192536 84182
rect 192484 84118 192536 84124
rect 183480 83473 183508 84118
rect 183466 83464 183522 83473
rect 183466 83399 183522 83408
rect 183006 82104 183062 82113
rect 183006 82039 183062 82048
rect 182916 79144 182968 79150
rect 182916 79086 182968 79092
rect 183020 60722 183048 82039
rect 200120 79076 200172 79082
rect 200120 79018 200172 79024
rect 195980 76356 196032 76362
rect 195980 76298 196032 76304
rect 193218 66872 193274 66881
rect 193218 66807 193274 66816
rect 183008 60716 183060 60722
rect 183008 60658 183060 60664
rect 183560 49292 183612 49298
rect 183560 49234 183612 49240
rect 182824 24132 182876 24138
rect 182824 24074 182876 24080
rect 183572 16574 183600 49234
rect 191838 47832 191894 47841
rect 191838 47767 191894 47776
rect 187700 46368 187752 46374
rect 187700 46310 187752 46316
rect 185032 43580 185084 43586
rect 185032 43522 185084 43528
rect 183572 16546 183784 16574
rect 183756 480 183784 16546
rect 185044 6914 185072 43522
rect 186320 27124 186372 27130
rect 186320 27066 186372 27072
rect 186332 16574 186360 27066
rect 187712 16574 187740 46310
rect 191852 16574 191880 47767
rect 186332 16546 186912 16574
rect 187712 16546 188568 16574
rect 191852 16546 192064 16574
rect 184952 6886 185072 6914
rect 184952 480 184980 6886
rect 186136 4140 186188 4146
rect 186136 4082 186188 4088
rect 186148 480 186176 4082
rect 182518 354 182630 480
rect 182192 326 182630 354
rect 181414 -960 181526 326
rect 182518 -960 182630 326
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 186884 354 186912 16546
rect 188540 480 188568 16546
rect 190828 6112 190880 6118
rect 190828 6054 190880 6060
rect 189724 4072 189776 4078
rect 189724 4014 189776 4020
rect 189736 480 189764 4014
rect 190840 480 190868 6054
rect 192036 480 192064 16546
rect 193232 480 193260 66807
rect 193310 27024 193366 27033
rect 193310 26959 193366 26968
rect 193324 16574 193352 26959
rect 195992 16574 196020 76298
rect 197360 75540 197412 75546
rect 197360 75482 197412 75488
rect 197372 16574 197400 75482
rect 198740 24404 198792 24410
rect 198740 24346 198792 24352
rect 193324 16546 194456 16574
rect 195992 16546 196848 16574
rect 197372 16546 197952 16574
rect 194428 480 194456 16546
rect 195612 3324 195664 3330
rect 195612 3266 195664 3272
rect 195624 480 195652 3266
rect 196820 480 196848 16546
rect 197924 480 197952 16546
rect 187302 354 187414 480
rect 186884 326 187414 354
rect 187302 -960 187414 326
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 198752 354 198780 24346
rect 200132 16574 200160 79018
rect 201512 78810 201540 702986
rect 218992 700670 219020 703520
rect 218980 700664 219032 700670
rect 218980 700606 219032 700612
rect 214564 524476 214616 524482
rect 214564 524418 214616 524424
rect 211804 470620 211856 470626
rect 211804 470562 211856 470568
rect 207664 229832 207716 229838
rect 207664 229774 207716 229780
rect 207676 203590 207704 229774
rect 207664 203584 207716 203590
rect 207664 203526 207716 203532
rect 211816 95198 211844 470562
rect 212552 229838 212580 230588
rect 212540 229832 212592 229838
rect 212540 229774 212592 229780
rect 214576 96626 214604 524418
rect 224224 364404 224276 364410
rect 224224 364346 224276 364352
rect 221464 311908 221516 311914
rect 221464 311850 221516 311856
rect 220084 258120 220136 258126
rect 220084 258062 220136 258068
rect 217324 218068 217376 218074
rect 217324 218010 217376 218016
rect 215944 178084 215996 178090
rect 215944 178026 215996 178032
rect 214564 96620 214616 96626
rect 214564 96562 214616 96568
rect 211804 95192 211856 95198
rect 211804 95134 211856 95140
rect 215956 87650 215984 178026
rect 217336 89010 217364 218010
rect 220096 90370 220124 258062
rect 221476 91798 221504 311850
rect 224236 93158 224264 364346
rect 234632 147014 234660 703582
rect 235000 703474 235028 703582
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299492 703582 299980 703610
rect 235184 703474 235212 703520
rect 235000 703446 235212 703474
rect 267660 697610 267688 703520
rect 283852 700602 283880 703520
rect 283840 700596 283892 700602
rect 283840 700538 283892 700544
rect 266360 697604 266412 697610
rect 266360 697546 266412 697552
rect 267648 697604 267700 697610
rect 267648 697546 267700 697552
rect 242912 204950 242940 230588
rect 242900 204944 242952 204950
rect 242900 204886 242952 204892
rect 234620 147008 234672 147014
rect 234620 146950 234672 146956
rect 224224 93152 224276 93158
rect 224224 93094 224276 93100
rect 221464 91792 221516 91798
rect 221464 91734 221516 91740
rect 220084 90364 220136 90370
rect 220084 90306 220136 90312
rect 217324 89004 217376 89010
rect 217324 88946 217376 88952
rect 215944 87644 215996 87650
rect 215944 87586 215996 87592
rect 231860 80300 231912 80306
rect 231860 80242 231912 80248
rect 213920 78940 213972 78946
rect 213920 78882 213972 78888
rect 201500 78804 201552 78810
rect 201500 78746 201552 78752
rect 209780 74180 209832 74186
rect 209780 74122 209832 74128
rect 202880 68604 202932 68610
rect 202880 68546 202932 68552
rect 201500 28552 201552 28558
rect 201500 28494 201552 28500
rect 200132 16546 200344 16574
rect 200316 480 200344 16546
rect 201512 480 201540 28494
rect 201592 25900 201644 25906
rect 201592 25842 201644 25848
rect 201604 16574 201632 25842
rect 202892 16574 202920 68546
rect 207020 64456 207072 64462
rect 207020 64398 207072 64404
rect 204260 51876 204312 51882
rect 204260 51818 204312 51824
rect 204272 16574 204300 51818
rect 201604 16546 202736 16574
rect 202892 16546 203472 16574
rect 204272 16546 205128 16574
rect 202708 480 202736 16546
rect 199078 354 199190 480
rect 198752 326 199190 354
rect 199078 -960 199190 326
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203444 354 203472 16546
rect 205100 480 205128 16546
rect 206192 5092 206244 5098
rect 206192 5034 206244 5040
rect 206204 480 206232 5034
rect 203862 354 203974 480
rect 203444 326 203974 354
rect 203862 -960 203974 326
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207032 354 207060 64398
rect 208400 45076 208452 45082
rect 208400 45018 208452 45024
rect 208412 16574 208440 45018
rect 208412 16546 208624 16574
rect 208596 480 208624 16546
rect 209792 480 209820 74122
rect 209872 70032 209924 70038
rect 209872 69974 209924 69980
rect 209884 16574 209912 69974
rect 212538 17368 212594 17377
rect 212538 17303 212594 17312
rect 212552 16574 212580 17303
rect 213932 16574 213960 78882
rect 226340 77172 226392 77178
rect 226340 77114 226392 77120
rect 216680 74112 216732 74118
rect 216680 74054 216732 74060
rect 215300 47728 215352 47734
rect 215300 47670 215352 47676
rect 209884 16546 211016 16574
rect 212552 16546 213408 16574
rect 213932 16546 214512 16574
rect 210988 480 211016 16546
rect 212172 3392 212224 3398
rect 212172 3334 212224 3340
rect 212184 480 212212 3334
rect 213380 480 213408 16546
rect 214484 480 214512 16546
rect 207358 354 207470 480
rect 207032 326 207470 354
rect 207358 -960 207470 326
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215312 354 215340 47670
rect 216692 16574 216720 74054
rect 223580 74044 223632 74050
rect 223580 73986 223632 73992
rect 218060 65680 218112 65686
rect 218060 65622 218112 65628
rect 216692 16546 216904 16574
rect 216876 480 216904 16546
rect 218072 480 218100 65622
rect 220820 64388 220872 64394
rect 220820 64330 220872 64336
rect 218152 42220 218204 42226
rect 218152 42162 218204 42168
rect 218164 16574 218192 42162
rect 219440 32428 219492 32434
rect 219440 32370 219492 32376
rect 219452 16574 219480 32370
rect 220832 16574 220860 64330
rect 218164 16546 219296 16574
rect 219452 16546 220032 16574
rect 220832 16546 221136 16574
rect 219268 480 219296 16546
rect 215638 354 215750 480
rect 215312 326 215750 354
rect 215638 -960 215750 326
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220004 354 220032 16546
rect 220422 354 220534 480
rect 220004 326 220534 354
rect 221108 354 221136 16546
rect 222752 7948 222804 7954
rect 222752 7890 222804 7896
rect 222764 480 222792 7890
rect 221526 354 221638 480
rect 221108 326 221638 354
rect 220422 -960 220534 326
rect 221526 -960 221638 326
rect 222722 -960 222834 480
rect 223592 354 223620 73986
rect 224960 61668 225012 61674
rect 224960 61610 225012 61616
rect 224972 16574 225000 61610
rect 224972 16546 225184 16574
rect 225156 480 225184 16546
rect 226352 480 226380 77114
rect 230478 74216 230534 74225
rect 230478 74151 230534 74160
rect 227718 61432 227774 61441
rect 227718 61367 227774 61376
rect 226430 32736 226486 32745
rect 226430 32671 226486 32680
rect 226444 16574 226472 32671
rect 227732 16574 227760 61367
rect 230492 16574 230520 74151
rect 226444 16546 227576 16574
rect 227732 16546 228312 16574
rect 230492 16546 231072 16574
rect 227548 480 227576 16546
rect 223918 354 224030 480
rect 223592 326 224030 354
rect 223918 -960 224030 326
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228284 354 228312 16546
rect 229374 13288 229430 13297
rect 229374 13223 229430 13232
rect 228702 354 228814 480
rect 228284 326 228814 354
rect 229388 354 229416 13223
rect 231044 480 231072 16546
rect 229806 354 229918 480
rect 229388 326 229918 354
rect 228702 -960 228814 326
rect 229806 -960 229918 326
rect 231002 -960 231114 480
rect 231872 354 231900 80242
rect 249800 80232 249852 80238
rect 249800 80174 249852 80180
rect 242164 78464 242216 78470
rect 242164 78406 242216 78412
rect 240140 77104 240192 77110
rect 240140 77046 240192 77052
rect 238760 68536 238812 68542
rect 238760 68478 238812 68484
rect 234620 65612 234672 65618
rect 234620 65554 234672 65560
rect 233240 50652 233292 50658
rect 233240 50594 233292 50600
rect 233252 16574 233280 50594
rect 233252 16546 233464 16574
rect 233436 480 233464 16546
rect 234632 11694 234660 65554
rect 236000 46300 236052 46306
rect 236000 46242 236052 46248
rect 234712 18896 234764 18902
rect 234712 18838 234764 18844
rect 234620 11688 234672 11694
rect 234620 11630 234672 11636
rect 234724 6914 234752 18838
rect 236012 16574 236040 46242
rect 238772 16574 238800 68478
rect 236012 16546 236592 16574
rect 238772 16546 239352 16574
rect 235816 11688 235868 11694
rect 235816 11630 235868 11636
rect 234632 6886 234752 6914
rect 234632 480 234660 6886
rect 235828 480 235856 11630
rect 232198 354 232310 480
rect 231872 326 232310 354
rect 232198 -960 232310 326
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236564 354 236592 16546
rect 237656 16108 237708 16114
rect 237656 16050 237708 16056
rect 236982 354 237094 480
rect 236564 326 237094 354
rect 237668 354 237696 16050
rect 239324 480 239352 16546
rect 238086 354 238198 480
rect 237668 326 238198 354
rect 236982 -960 237094 326
rect 238086 -960 238198 326
rect 239282 -960 239394 480
rect 240152 354 240180 77046
rect 242176 20058 242204 78406
rect 247038 77072 247094 77081
rect 247038 77007 247094 77016
rect 244278 74080 244334 74089
rect 244278 74015 244334 74024
rect 242900 62960 242952 62966
rect 242900 62902 242952 62908
rect 241520 20052 241572 20058
rect 241520 19994 241572 20000
rect 242164 20052 242216 20058
rect 242164 19994 242216 20000
rect 241532 16574 241560 19994
rect 241532 16546 241744 16574
rect 241716 480 241744 16546
rect 242912 480 242940 62902
rect 242992 28484 243044 28490
rect 242992 28426 243044 28432
rect 243004 16574 243032 28426
rect 244292 16574 244320 74015
rect 245658 64288 245714 64297
rect 245658 64223 245714 64232
rect 245672 16574 245700 64223
rect 247052 16574 247080 77007
rect 248418 20088 248474 20097
rect 248418 20023 248474 20032
rect 243004 16546 244136 16574
rect 244292 16546 245240 16574
rect 245672 16546 245976 16574
rect 247052 16546 247632 16574
rect 244108 480 244136 16546
rect 245212 480 245240 16546
rect 240478 354 240590 480
rect 240152 326 240590 354
rect 240478 -960 240590 326
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 245948 354 245976 16546
rect 247604 480 247632 16546
rect 246366 354 246478 480
rect 245948 326 246478 354
rect 246366 -960 246478 326
rect 247562 -960 247674 480
rect 248432 354 248460 20023
rect 249812 16574 249840 80174
rect 252560 79008 252612 79014
rect 266372 78985 266400 697546
rect 272536 228410 272564 230588
rect 272524 228404 272576 228410
rect 272524 228346 272576 228352
rect 299492 145586 299520 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429212 703582 429700 703610
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 332520 703050 332548 703520
rect 331220 703044 331272 703050
rect 331220 702986 331272 702992
rect 332508 703044 332560 703050
rect 332508 702986 332560 702992
rect 302252 230574 302542 230602
rect 302252 196654 302280 230574
rect 302240 196648 302292 196654
rect 302240 196590 302292 196596
rect 299480 145580 299532 145586
rect 299480 145522 299532 145528
rect 284300 80164 284352 80170
rect 284300 80106 284352 80112
rect 252560 78950 252612 78956
rect 266358 78976 266414 78985
rect 251180 73976 251232 73982
rect 251180 73918 251232 73924
rect 249812 16546 250024 16574
rect 249996 480 250024 16546
rect 251192 4078 251220 73918
rect 251272 29980 251324 29986
rect 251272 29922 251324 29928
rect 251180 4072 251232 4078
rect 251180 4014 251232 4020
rect 251284 3482 251312 29922
rect 252572 16574 252600 78950
rect 266358 78911 266414 78920
rect 255962 78024 256018 78033
rect 255962 77959 256018 77968
rect 253940 29912 253992 29918
rect 253940 29854 253992 29860
rect 253952 16574 253980 29854
rect 255976 20126 256004 77959
rect 260840 77036 260892 77042
rect 260840 76978 260892 76984
rect 256700 67108 256752 67114
rect 256700 67050 256752 67056
rect 255320 20120 255372 20126
rect 255320 20062 255372 20068
rect 255964 20120 256016 20126
rect 255964 20062 256016 20068
rect 255332 16574 255360 20062
rect 252572 16546 253520 16574
rect 253952 16546 254256 16574
rect 255332 16546 255912 16574
rect 252376 4072 252428 4078
rect 252376 4014 252428 4020
rect 251192 3454 251312 3482
rect 251192 480 251220 3454
rect 252388 480 252416 4014
rect 253492 480 253520 16546
rect 248758 354 248870 480
rect 248432 326 248870 354
rect 248758 -960 248870 326
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254228 354 254256 16546
rect 255884 480 255912 16546
rect 254646 354 254758 480
rect 254228 326 254758 354
rect 254646 -960 254758 326
rect 255842 -960 255954 480
rect 256712 354 256740 67050
rect 259460 60308 259512 60314
rect 259460 60250 259512 60256
rect 258080 38004 258132 38010
rect 258080 37946 258132 37952
rect 258092 16574 258120 37946
rect 258092 16546 258304 16574
rect 258276 480 258304 16546
rect 259472 11694 259500 60250
rect 259552 33992 259604 33998
rect 259552 33934 259604 33940
rect 259460 11688 259512 11694
rect 259460 11630 259512 11636
rect 259564 6914 259592 33934
rect 260852 16574 260880 76978
rect 267740 76968 267792 76974
rect 267740 76910 267792 76916
rect 282918 76936 282974 76945
rect 263598 62928 263654 62937
rect 263598 62863 263654 62872
rect 262220 20188 262272 20194
rect 262220 20130 262272 20136
rect 262232 16574 262260 20130
rect 263612 16574 263640 62863
rect 266358 52048 266414 52057
rect 266358 51983 266414 51992
rect 264978 39264 265034 39273
rect 264978 39199 265034 39208
rect 260852 16546 261800 16574
rect 262232 16546 262536 16574
rect 263612 16546 264192 16574
rect 260656 11688 260708 11694
rect 260656 11630 260708 11636
rect 259472 6886 259592 6914
rect 259472 480 259500 6886
rect 260668 480 260696 11630
rect 261772 480 261800 16546
rect 257038 354 257150 480
rect 256712 326 257150 354
rect 257038 -960 257150 326
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262508 354 262536 16546
rect 264164 480 264192 16546
rect 262926 354 263038 480
rect 262508 326 263038 354
rect 262926 -960 263038 326
rect 264122 -960 264234 480
rect 264992 354 265020 39199
rect 266372 16574 266400 51983
rect 266372 16546 266584 16574
rect 266556 480 266584 16546
rect 267752 480 267780 76910
rect 282918 76871 282974 76880
rect 282932 16574 282960 76871
rect 282932 16546 283144 16574
rect 279514 9616 279570 9625
rect 279514 9551 279570 9560
rect 270040 9444 270092 9450
rect 270040 9386 270092 9392
rect 268844 6860 268896 6866
rect 268844 6802 268896 6808
rect 268856 480 268884 6802
rect 270052 480 270080 9386
rect 277124 9376 277176 9382
rect 277124 9318 277176 9324
rect 276020 9308 276072 9314
rect 276020 9250 276072 9256
rect 272432 6792 272484 6798
rect 272432 6734 272484 6740
rect 271236 4004 271288 4010
rect 271236 3946 271288 3952
rect 271248 480 271276 3946
rect 272444 480 272472 6734
rect 273628 6724 273680 6730
rect 273628 6666 273680 6672
rect 273640 480 273668 6666
rect 274824 3936 274876 3942
rect 274824 3878 274876 3884
rect 274836 480 274864 3878
rect 276032 480 276060 9250
rect 277136 480 277164 9318
rect 278320 3868 278372 3874
rect 278320 3810 278372 3816
rect 278332 480 278360 3810
rect 279528 480 279556 9551
rect 280710 9480 280766 9489
rect 280710 9415 280766 9424
rect 280724 480 280752 9415
rect 281906 3768 281962 3777
rect 281906 3703 281962 3712
rect 281920 480 281948 3703
rect 283116 480 283144 16546
rect 284312 3874 284340 80106
rect 331232 79558 331260 702986
rect 348804 700534 348832 703520
rect 364996 702434 365024 703520
rect 364352 702406 365024 702434
rect 348792 700528 348844 700534
rect 348792 700470 348844 700476
rect 332612 198014 332640 230588
rect 362972 199442 363000 230588
rect 362960 199436 363012 199442
rect 362960 199378 363012 199384
rect 332600 198008 332652 198014
rect 332600 197950 332652 197956
rect 364352 140146 364380 702406
rect 392504 229770 392532 230588
rect 392492 229764 392544 229770
rect 392492 229706 392544 229712
rect 364340 140140 364392 140146
rect 364340 140082 364392 140088
rect 374000 79688 374052 79694
rect 374000 79630 374052 79636
rect 331220 79552 331272 79558
rect 331220 79494 331272 79500
rect 306380 78872 306432 78878
rect 306380 78814 306432 78820
rect 288440 76900 288492 76906
rect 288440 76842 288492 76848
rect 284390 73944 284446 73953
rect 284390 73879 284446 73888
rect 284300 3868 284352 3874
rect 284300 3810 284352 3816
rect 284404 3482 284432 73879
rect 285680 42152 285732 42158
rect 285680 42094 285732 42100
rect 285692 16574 285720 42094
rect 287060 33924 287112 33930
rect 287060 33866 287112 33872
rect 287072 16574 287100 33866
rect 288452 16574 288480 76842
rect 296720 76832 296772 76838
rect 296720 76774 296772 76780
rect 291200 35420 291252 35426
rect 291200 35362 291252 35368
rect 291212 16574 291240 35362
rect 292672 24336 292724 24342
rect 292672 24278 292724 24284
rect 292684 16574 292712 24278
rect 296732 16574 296760 76774
rect 302240 76764 302292 76770
rect 302240 76706 302292 76712
rect 298098 72448 298154 72457
rect 298098 72383 298154 72392
rect 285692 16546 286640 16574
rect 287072 16546 287376 16574
rect 288452 16546 289032 16574
rect 291212 16546 291424 16574
rect 292684 16546 293264 16574
rect 296732 16546 297312 16574
rect 285036 3868 285088 3874
rect 285036 3810 285088 3816
rect 284312 3454 284432 3482
rect 284312 480 284340 3454
rect 265318 354 265430 480
rect 264992 326 265430 354
rect 265318 -960 265430 326
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285048 354 285076 3810
rect 286612 480 286640 16546
rect 285374 354 285486 480
rect 285048 326 285486 354
rect 285374 -960 285486 326
rect 286570 -960 286682 480
rect 287348 354 287376 16546
rect 289004 480 289032 16546
rect 289820 14748 289872 14754
rect 289820 14690 289872 14696
rect 287766 354 287878 480
rect 287348 326 287878 354
rect 287766 -960 287878 326
rect 288962 -960 289074 480
rect 289832 354 289860 14690
rect 291396 480 291424 16546
rect 292580 3800 292632 3806
rect 292580 3742 292632 3748
rect 292592 480 292620 3742
rect 290158 354 290270 480
rect 289832 326 290270 354
rect 290158 -960 290270 326
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293236 354 293264 16546
rect 296076 6656 296128 6662
rect 296076 6598 296128 6604
rect 294880 5024 294932 5030
rect 294880 4966 294932 4972
rect 294892 480 294920 4966
rect 296088 480 296116 6598
rect 297284 480 297312 16546
rect 293654 354 293766 480
rect 293236 326 293766 354
rect 293654 -960 293766 326
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298112 354 298140 72383
rect 300858 17232 300914 17241
rect 300858 17167 300914 17176
rect 300872 16574 300900 17167
rect 302252 16574 302280 76706
rect 305000 35352 305052 35358
rect 305000 35294 305052 35300
rect 303620 25832 303672 25838
rect 303620 25774 303672 25780
rect 303632 16574 303660 25774
rect 305012 16574 305040 35294
rect 300872 16546 301544 16574
rect 302252 16546 303200 16574
rect 303632 16546 303936 16574
rect 305012 16546 305592 16574
rect 299662 6624 299718 6633
rect 299662 6559 299718 6568
rect 299676 480 299704 6559
rect 300766 6488 300822 6497
rect 300766 6423 300822 6432
rect 300780 480 300808 6423
rect 298438 354 298550 480
rect 298112 326 298550 354
rect 298438 -960 298550 326
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301516 354 301544 16546
rect 303172 480 303200 16546
rect 301934 354 302046 480
rect 301516 326 302046 354
rect 301934 -960 302046 326
rect 303130 -960 303242 480
rect 303908 354 303936 16546
rect 305564 480 305592 16546
rect 304326 354 304438 480
rect 303908 326 304438 354
rect 304326 -960 304438 326
rect 305522 -960 305634 480
rect 306392 354 306420 78814
rect 315304 78396 315356 78402
rect 315304 78338 315356 78344
rect 307760 72820 307812 72826
rect 307760 72762 307812 72768
rect 307772 3398 307800 72762
rect 311900 72752 311952 72758
rect 311900 72694 311952 72700
rect 309140 58812 309192 58818
rect 309140 58754 309192 58760
rect 309152 16574 309180 58754
rect 311912 16574 311940 72694
rect 313280 24268 313332 24274
rect 313280 24210 313332 24216
rect 313292 16574 313320 24210
rect 309152 16546 309824 16574
rect 311912 16546 312216 16574
rect 313292 16546 313872 16574
rect 307944 7880 307996 7886
rect 307944 7822 307996 7828
rect 307760 3392 307812 3398
rect 307760 3334 307812 3340
rect 307956 480 307984 7822
rect 309048 3392 309100 3398
rect 309048 3334 309100 3340
rect 309060 480 309088 3334
rect 306718 354 306830 480
rect 306392 326 306830 354
rect 306718 -960 306830 326
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 309796 354 309824 16546
rect 311440 14680 311492 14686
rect 311440 14622 311492 14628
rect 311452 480 311480 14622
rect 310214 354 310326 480
rect 309796 326 310326 354
rect 310214 -960 310326 326
rect 311410 -960 311522 480
rect 312188 354 312216 16546
rect 313844 480 313872 16546
rect 315316 9246 315344 78338
rect 354678 76800 354734 76809
rect 354678 76735 354734 76744
rect 347780 73908 347832 73914
rect 347780 73850 347832 73856
rect 318798 73808 318854 73817
rect 318798 73743 318854 73752
rect 316038 55992 316094 56001
rect 316038 55927 316094 55936
rect 315028 9240 315080 9246
rect 315028 9182 315080 9188
rect 315304 9240 315356 9246
rect 315304 9182 315356 9188
rect 315040 480 315068 9182
rect 316052 3398 316080 55927
rect 316130 42120 316186 42129
rect 316130 42055 316186 42064
rect 316144 16574 316172 42055
rect 317418 26888 317474 26897
rect 317418 26823 317474 26832
rect 317432 16574 317460 26823
rect 318812 16574 318840 73743
rect 325700 72684 325752 72690
rect 325700 72626 325752 72632
rect 320180 68468 320232 68474
rect 320180 68410 320232 68416
rect 320192 16574 320220 68410
rect 324320 62892 324372 62898
rect 324320 62834 324372 62840
rect 316144 16546 316264 16574
rect 317432 16546 318104 16574
rect 318812 16546 319760 16574
rect 320192 16546 320496 16574
rect 316040 3392 316092 3398
rect 316040 3334 316092 3340
rect 316236 480 316264 16546
rect 317328 3392 317380 3398
rect 317328 3334 317380 3340
rect 317340 480 317368 3334
rect 312606 354 312718 480
rect 312188 326 312718 354
rect 312606 -960 312718 326
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 354 318104 16546
rect 319732 480 319760 16546
rect 318494 354 318606 480
rect 318076 326 318606 354
rect 318494 -960 318606 326
rect 319690 -960 319802 480
rect 320468 354 320496 16546
rect 322112 10464 322164 10470
rect 322112 10406 322164 10412
rect 322124 480 322152 10406
rect 323308 7812 323360 7818
rect 323308 7754 323360 7760
rect 323320 480 323348 7754
rect 324332 3210 324360 62834
rect 324412 29844 324464 29850
rect 324412 29786 324464 29792
rect 324424 3398 324452 29786
rect 325712 16574 325740 72626
rect 332600 72616 332652 72622
rect 332600 72558 332652 72564
rect 327080 60240 327132 60246
rect 327080 60182 327132 60188
rect 327092 16574 327120 60182
rect 331220 54800 331272 54806
rect 331220 54742 331272 54748
rect 328460 42084 328512 42090
rect 328460 42026 328512 42032
rect 328472 16574 328500 42026
rect 329840 31136 329892 31142
rect 329840 31078 329892 31084
rect 329852 16574 329880 31078
rect 325712 16546 326384 16574
rect 327092 16546 328040 16574
rect 328472 16546 328776 16574
rect 329852 16546 330432 16574
rect 324412 3392 324464 3398
rect 324412 3334 324464 3340
rect 325608 3392 325660 3398
rect 325608 3334 325660 3340
rect 324332 3182 324452 3210
rect 324424 480 324452 3182
rect 325620 480 325648 3334
rect 320886 354 320998 480
rect 320468 326 320998 354
rect 320886 -960 320998 326
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326356 354 326384 16546
rect 328012 480 328040 16546
rect 326774 354 326886 480
rect 326356 326 326886 354
rect 326774 -960 326886 326
rect 327970 -960 328082 480
rect 328748 354 328776 16546
rect 330404 480 330432 16546
rect 329166 354 329278 480
rect 328748 326 329278 354
rect 329166 -960 329278 326
rect 330362 -960 330474 480
rect 331232 354 331260 54742
rect 332612 3398 332640 72558
rect 340880 72548 340932 72554
rect 340880 72490 340932 72496
rect 333978 51912 334034 51921
rect 333978 51847 334034 51856
rect 332692 31204 332744 31210
rect 332692 31146 332744 31152
rect 332600 3392 332652 3398
rect 332600 3334 332652 3340
rect 332704 480 332732 31146
rect 333992 16574 334020 51847
rect 339500 45008 339552 45014
rect 339500 44950 339552 44956
rect 338120 37936 338172 37942
rect 338120 37878 338172 37884
rect 336738 35320 336794 35329
rect 336738 35255 336794 35264
rect 336752 16574 336780 35255
rect 338132 16574 338160 37878
rect 333992 16546 334664 16574
rect 336752 16546 337056 16574
rect 338132 16546 338712 16574
rect 333888 3392 333940 3398
rect 333888 3334 333940 3340
rect 333900 480 333928 3334
rect 331558 354 331670 480
rect 331232 326 331670 354
rect 331558 -960 331670 326
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 354 334664 16546
rect 336278 11792 336334 11801
rect 336278 11727 336334 11736
rect 336292 480 336320 11727
rect 335054 354 335166 480
rect 334636 326 335166 354
rect 335054 -960 335166 326
rect 336250 -960 336362 480
rect 337028 354 337056 16546
rect 338684 480 338712 16546
rect 337446 354 337558 480
rect 337028 326 337558 354
rect 337446 -960 337558 326
rect 338642 -960 338754 480
rect 339512 354 339540 44950
rect 340892 3210 340920 72490
rect 343640 72480 343692 72486
rect 343640 72422 343692 72428
rect 340972 58744 341024 58750
rect 340972 58686 341024 58692
rect 340984 3398 341012 58686
rect 343652 16574 343680 72422
rect 345020 57520 345072 57526
rect 345020 57462 345072 57468
rect 345032 16574 345060 57462
rect 346400 28416 346452 28422
rect 346400 28358 346452 28364
rect 346412 16574 346440 28358
rect 347792 16574 347820 73850
rect 353298 68368 353354 68377
rect 353298 68303 353354 68312
rect 351918 47696 351974 47705
rect 351918 47631 351974 47640
rect 349160 43512 349212 43518
rect 349160 43454 349212 43460
rect 343652 16546 344600 16574
rect 345032 16546 345336 16574
rect 346412 16546 346992 16574
rect 347792 16546 348096 16574
rect 342904 16040 342956 16046
rect 342904 15982 342956 15988
rect 340972 3392 341024 3398
rect 340972 3334 341024 3340
rect 342168 3392 342220 3398
rect 342168 3334 342220 3340
rect 340892 3182 341012 3210
rect 340984 480 341012 3182
rect 342180 480 342208 3334
rect 339838 354 339950 480
rect 339512 326 339950 354
rect 339838 -960 339950 326
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342916 354 342944 15982
rect 344572 480 344600 16546
rect 343334 354 343446 480
rect 342916 326 343446 354
rect 343334 -960 343446 326
rect 344530 -960 344642 480
rect 345308 354 345336 16546
rect 346964 480 346992 16546
rect 348068 480 348096 16546
rect 349172 3210 349200 43454
rect 350538 35184 350594 35193
rect 350538 35119 350594 35128
rect 350552 16574 350580 35119
rect 351932 16574 351960 47631
rect 353312 16574 353340 68303
rect 354692 16574 354720 76735
rect 356060 76696 356112 76702
rect 356060 76638 356112 76644
rect 356072 16574 356100 76638
rect 358820 75472 358872 75478
rect 358820 75414 358872 75420
rect 357440 49224 357492 49230
rect 357440 49166 357492 49172
rect 357452 16574 357480 49166
rect 358832 16574 358860 75414
rect 367100 65544 367152 65550
rect 367100 65486 367152 65492
rect 362960 64320 363012 64326
rect 362960 64262 363012 64268
rect 362972 16574 363000 64262
rect 365720 55956 365772 55962
rect 365720 55898 365772 55904
rect 350552 16546 351224 16574
rect 351932 16546 352880 16574
rect 353312 16546 353616 16574
rect 354692 16546 355272 16574
rect 356072 16546 356376 16574
rect 357452 16546 357572 16574
rect 358832 16546 359504 16574
rect 362972 16546 363552 16574
rect 349252 13252 349304 13258
rect 349252 13194 349304 13200
rect 349264 3398 349292 13194
rect 349252 3392 349304 3398
rect 349252 3334 349304 3340
rect 350448 3392 350500 3398
rect 350448 3334 350500 3340
rect 349172 3182 349292 3210
rect 349264 480 349292 3182
rect 350460 480 350488 3334
rect 345726 354 345838 480
rect 345308 326 345838 354
rect 345726 -960 345838 326
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351196 354 351224 16546
rect 352852 480 352880 16546
rect 351614 354 351726 480
rect 351196 326 351726 354
rect 351614 -960 351726 326
rect 352810 -960 352922 480
rect 353588 354 353616 16546
rect 355244 480 355272 16546
rect 356348 480 356376 16546
rect 357544 480 357572 16546
rect 358728 9172 358780 9178
rect 358728 9114 358780 9120
rect 358740 480 358768 9114
rect 354006 354 354118 480
rect 353588 326 354118 354
rect 354006 -960 354118 326
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359476 354 359504 16546
rect 361120 15972 361172 15978
rect 361120 15914 361172 15920
rect 361132 480 361160 15914
rect 361856 13184 361908 13190
rect 361856 13126 361908 13132
rect 359894 354 360006 480
rect 359476 326 360006 354
rect 359894 -960 360006 326
rect 361090 -960 361202 480
rect 361868 354 361896 13126
rect 363524 480 363552 16546
rect 364616 4956 364668 4962
rect 364616 4898 364668 4904
rect 364628 480 364656 4898
rect 365732 3398 365760 55898
rect 367112 16574 367140 65486
rect 368480 61600 368532 61606
rect 368480 61542 368532 61548
rect 368492 16574 368520 61542
rect 369858 51776 369914 51785
rect 369858 51711 369914 51720
rect 369872 16574 369900 51711
rect 372618 21584 372674 21593
rect 372618 21519 372674 21528
rect 372632 16574 372660 21519
rect 367112 16546 367784 16574
rect 368492 16546 369440 16574
rect 369872 16546 370176 16574
rect 372632 16546 372936 16574
rect 365810 15872 365866 15881
rect 365810 15807 365866 15816
rect 365720 3392 365772 3398
rect 365720 3334 365772 3340
rect 365824 480 365852 15807
rect 367008 3392 367060 3398
rect 367008 3334 367060 3340
rect 367020 480 367048 3334
rect 362286 354 362398 480
rect 361868 326 362398 354
rect 362286 -960 362398 326
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 367756 354 367784 16546
rect 369412 480 369440 16546
rect 368174 354 368286 480
rect 367756 326 368286 354
rect 368174 -960 368286 326
rect 369370 -960 369482 480
rect 370148 354 370176 16546
rect 371238 13152 371294 13161
rect 371238 13087 371294 13096
rect 370566 354 370678 480
rect 370148 326 370678 354
rect 371252 354 371280 13087
rect 372908 480 372936 16546
rect 374012 1170 374040 79630
rect 397472 78849 397500 703520
rect 413664 700466 413692 703520
rect 413652 700460 413704 700466
rect 413652 700402 413704 700408
rect 429212 144226 429240 703582
rect 429672 703474 429700 703582
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494072 703582 494652 703610
rect 429856 703474 429884 703520
rect 429672 703446 429884 703474
rect 429200 144220 429252 144226
rect 429200 144162 429252 144168
rect 426440 80096 426492 80102
rect 426440 80038 426492 80044
rect 397458 78840 397514 78849
rect 397458 78775 397514 78784
rect 389178 76664 389234 76673
rect 389178 76599 389234 76608
rect 382280 71324 382332 71330
rect 382280 71266 382332 71272
rect 374092 64252 374144 64258
rect 374092 64194 374144 64200
rect 374104 3398 374132 64194
rect 376760 64184 376812 64190
rect 376760 64126 376812 64132
rect 375380 35284 375432 35290
rect 375380 35226 375432 35232
rect 375392 16574 375420 35226
rect 376772 16574 376800 64126
rect 380900 54732 380952 54738
rect 380900 54674 380952 54680
rect 378140 28348 378192 28354
rect 378140 28290 378192 28296
rect 378152 16574 378180 28290
rect 380912 16574 380940 54674
rect 375392 16546 376064 16574
rect 376772 16546 377720 16574
rect 378152 16546 378456 16574
rect 380912 16546 381216 16574
rect 374092 3392 374144 3398
rect 374092 3334 374144 3340
rect 375288 3392 375340 3398
rect 375288 3334 375340 3340
rect 374012 1142 374132 1170
rect 374104 480 374132 1142
rect 375300 480 375328 3334
rect 371670 354 371782 480
rect 371252 326 371782 354
rect 370566 -960 370678 326
rect 371670 -960 371782 326
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376036 354 376064 16546
rect 377692 480 377720 16546
rect 376454 354 376566 480
rect 376036 326 376566 354
rect 376454 -960 376566 326
rect 377650 -960 377762 480
rect 378428 354 378456 16546
rect 379520 10396 379572 10402
rect 379520 10338 379572 10344
rect 378846 354 378958 480
rect 378428 326 378958 354
rect 379532 354 379560 10338
rect 381188 480 381216 16546
rect 382292 3210 382320 71266
rect 383660 58676 383712 58682
rect 383660 58618 383712 58624
rect 382372 49156 382424 49162
rect 382372 49098 382424 49104
rect 382384 3398 382412 49098
rect 383672 16574 383700 58618
rect 387798 55856 387854 55865
rect 387798 55791 387854 55800
rect 383672 16546 384344 16574
rect 382372 3392 382424 3398
rect 382372 3334 382424 3340
rect 383568 3392 383620 3398
rect 383568 3334 383620 3340
rect 382292 3182 382412 3210
rect 382384 480 382412 3182
rect 383580 480 383608 3334
rect 379950 354 380062 480
rect 379532 326 380062 354
rect 378846 -960 378958 326
rect 379950 -960 380062 326
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384316 354 384344 16546
rect 386696 14612 386748 14618
rect 386696 14554 386748 14560
rect 385960 7744 386012 7750
rect 385960 7686 386012 7692
rect 385972 480 386000 7686
rect 384734 354 384846 480
rect 384316 326 384846 354
rect 384734 -960 384846 326
rect 385930 -960 386042 480
rect 386708 354 386736 14554
rect 387126 354 387238 480
rect 386708 326 387238 354
rect 387812 354 387840 55791
rect 389192 16574 389220 76599
rect 402978 75576 403034 75585
rect 402978 75511 403034 75520
rect 390560 73840 390612 73846
rect 390560 73782 390612 73788
rect 389192 16546 389496 16574
rect 389468 480 389496 16546
rect 390572 3210 390600 73782
rect 396080 67040 396132 67046
rect 396080 66982 396132 66988
rect 390652 61532 390704 61538
rect 390652 61474 390704 61480
rect 390664 3398 390692 61474
rect 394700 57452 394752 57458
rect 394700 57394 394752 57400
rect 391940 29776 391992 29782
rect 391940 29718 391992 29724
rect 391952 16574 391980 29718
rect 394712 16574 394740 57394
rect 391952 16546 392624 16574
rect 394712 16546 395384 16574
rect 390652 3392 390704 3398
rect 390652 3334 390704 3340
rect 391848 3392 391900 3398
rect 391848 3334 391900 3340
rect 390572 3182 390692 3210
rect 390664 480 390692 3182
rect 391860 480 391888 3334
rect 388230 354 388342 480
rect 387812 326 388342 354
rect 387126 -960 387238 326
rect 388230 -960 388342 326
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392596 354 392624 16546
rect 394240 6588 394292 6594
rect 394240 6530 394292 6536
rect 394252 480 394280 6530
rect 395356 480 395384 16546
rect 393014 354 393126 480
rect 392596 326 393126 354
rect 393014 -960 393126 326
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396092 354 396120 66982
rect 398840 54664 398892 54670
rect 398840 54606 398892 54612
rect 397460 28280 397512 28286
rect 397460 28222 397512 28228
rect 397472 16574 397500 28222
rect 397472 16546 397776 16574
rect 397748 480 397776 16546
rect 398852 3210 398880 54606
rect 398932 26988 398984 26994
rect 398932 26930 398984 26936
rect 398944 3398 398972 26930
rect 401600 25764 401652 25770
rect 401600 25706 401652 25712
rect 401612 16574 401640 25706
rect 402992 16574 403020 75511
rect 408500 71256 408552 71262
rect 408500 71198 408552 71204
rect 405738 47560 405794 47569
rect 405738 47495 405794 47504
rect 404360 23044 404412 23050
rect 404360 22986 404412 22992
rect 401612 16546 402560 16574
rect 402992 16546 403664 16574
rect 400864 11824 400916 11830
rect 400864 11766 400916 11772
rect 398932 3392 398984 3398
rect 398932 3334 398984 3340
rect 400128 3392 400180 3398
rect 400128 3334 400180 3340
rect 398852 3182 398972 3210
rect 398944 480 398972 3182
rect 400140 480 400168 3334
rect 396510 354 396622 480
rect 396092 326 396622 354
rect 396510 -960 396622 326
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 400876 354 400904 11766
rect 402532 480 402560 16546
rect 403636 480 403664 16546
rect 401294 354 401406 480
rect 400876 326 401406 354
rect 401294 -960 401406 326
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404372 354 404400 22986
rect 405752 16574 405780 47495
rect 407118 18592 407174 18601
rect 407118 18527 407174 18536
rect 405752 16546 406056 16574
rect 406028 480 406056 16546
rect 407132 3398 407160 18527
rect 408512 16574 408540 71198
rect 412640 61464 412692 61470
rect 412640 61406 412692 61412
rect 411260 27056 411312 27062
rect 411260 26998 411312 27004
rect 409880 22976 409932 22982
rect 409880 22918 409932 22924
rect 409892 16574 409920 22918
rect 411272 16574 411300 26998
rect 408512 16546 409184 16574
rect 409892 16546 410840 16574
rect 411272 16546 411944 16574
rect 407210 9344 407266 9353
rect 407210 9279 407266 9288
rect 407120 3392 407172 3398
rect 407120 3334 407172 3340
rect 407224 480 407252 9279
rect 408408 3392 408460 3398
rect 408408 3334 408460 3340
rect 408420 480 408448 3334
rect 404790 354 404902 480
rect 404372 326 404902 354
rect 404790 -960 404902 326
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409156 354 409184 16546
rect 410812 480 410840 16546
rect 411916 480 411944 16546
rect 409574 354 409686 480
rect 409156 326 409686 354
rect 409574 -960 409686 326
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 412652 354 412680 61406
rect 415400 55888 415452 55894
rect 415400 55830 415452 55836
rect 414020 25696 414072 25702
rect 414020 25638 414072 25644
rect 414032 16574 414060 25638
rect 414032 16546 414336 16574
rect 414308 480 414336 16546
rect 415412 3398 415440 55830
rect 419540 53372 419592 53378
rect 419540 53314 419592 53320
rect 418160 36576 418212 36582
rect 418160 36518 418212 36524
rect 416780 24200 416832 24206
rect 416780 24142 416832 24148
rect 415492 19984 415544 19990
rect 415492 19926 415544 19932
rect 415400 3392 415452 3398
rect 415400 3334 415452 3340
rect 415504 480 415532 19926
rect 416792 16574 416820 24142
rect 418172 16574 418200 36518
rect 419552 16574 419580 53314
rect 423678 48920 423734 48929
rect 423678 48855 423734 48864
rect 422298 19952 422354 19961
rect 422298 19887 422354 19896
rect 422312 16574 422340 19887
rect 416792 16546 417464 16574
rect 418172 16546 418568 16574
rect 419552 16546 420224 16574
rect 422312 16546 422616 16574
rect 416688 3392 416740 3398
rect 416688 3334 416740 3340
rect 416700 480 416728 3334
rect 413070 354 413182 480
rect 412652 326 413182 354
rect 413070 -960 413182 326
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417436 354 417464 16546
rect 417854 354 417966 480
rect 417436 326 417966 354
rect 418540 354 418568 16546
rect 420196 480 420224 16546
rect 420918 10296 420974 10305
rect 420918 10231 420974 10240
rect 418958 354 419070 480
rect 418540 326 419070 354
rect 417854 -960 417966 326
rect 418958 -960 419070 326
rect 420154 -960 420266 480
rect 420932 354 420960 10231
rect 422588 480 422616 16546
rect 423692 3210 423720 48855
rect 425060 44940 425112 44946
rect 425060 44882 425112 44888
rect 425072 16574 425100 44882
rect 426452 16574 426480 80038
rect 462332 78713 462360 703520
rect 478524 700398 478552 703520
rect 478512 700392 478564 700398
rect 478512 700334 478564 700340
rect 494072 141438 494100 703582
rect 494624 703474 494652 703582
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 494808 703474 494836 703520
rect 494624 703446 494836 703474
rect 494060 141432 494112 141438
rect 494060 141374 494112 141380
rect 462318 78704 462374 78713
rect 462318 78639 462374 78648
rect 430580 78328 430632 78334
rect 430580 78270 430632 78276
rect 427820 46232 427872 46238
rect 427820 46174 427872 46180
rect 427832 16574 427860 46174
rect 429200 33856 429252 33862
rect 429200 33798 429252 33804
rect 425072 16546 425744 16574
rect 426452 16546 426848 16574
rect 427832 16546 428504 16574
rect 423770 11656 423826 11665
rect 423770 11591 423826 11600
rect 423784 3398 423812 11591
rect 423772 3392 423824 3398
rect 423772 3334 423824 3340
rect 424968 3392 425020 3398
rect 424968 3334 425020 3340
rect 423692 3182 423812 3210
rect 423784 480 423812 3182
rect 424980 480 425008 3334
rect 421350 354 421462 480
rect 420932 326 421462 354
rect 421350 -960 421462 326
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 425716 354 425744 16546
rect 426134 354 426246 480
rect 425716 326 426246 354
rect 426820 354 426848 16546
rect 428476 480 428504 16546
rect 427238 354 427350 480
rect 426820 326 427350 354
rect 426134 -960 426246 326
rect 427238 -960 427350 326
rect 428434 -960 428546 480
rect 429212 354 429240 33798
rect 430592 16574 430620 78270
rect 436744 78260 436796 78266
rect 436744 78202 436796 78208
rect 431960 69964 432012 69970
rect 431960 69906 432012 69912
rect 430592 16546 430896 16574
rect 430868 480 430896 16546
rect 431972 1170 432000 69906
rect 433340 57384 433392 57390
rect 433340 57326 433392 57332
rect 432052 49088 432104 49094
rect 432052 49030 432104 49036
rect 432064 3398 432092 49030
rect 433352 16574 433380 57326
rect 434720 29708 434772 29714
rect 434720 29650 434772 29656
rect 434732 16574 434760 29650
rect 433352 16546 434024 16574
rect 434732 16546 435128 16574
rect 432052 3392 432104 3398
rect 432052 3334 432104 3340
rect 433248 3392 433300 3398
rect 433248 3334 433300 3340
rect 431972 1142 432092 1170
rect 432064 480 432092 1142
rect 433260 480 433288 3334
rect 429630 354 429742 480
rect 429212 326 429742 354
rect 429630 -960 429742 326
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 433996 354 434024 16546
rect 434414 354 434526 480
rect 433996 326 434526 354
rect 435100 354 435128 16546
rect 436756 5030 436784 78202
rect 480260 78192 480312 78198
rect 480260 78134 480312 78140
rect 459558 75440 459614 75449
rect 438860 75404 438912 75410
rect 459558 75375 459614 75384
rect 438860 75346 438912 75352
rect 437480 69896 437532 69902
rect 437480 69838 437532 69844
rect 436744 5024 436796 5030
rect 436744 4966 436796 4972
rect 436744 4888 436796 4894
rect 436744 4830 436796 4836
rect 436756 480 436784 4830
rect 435518 354 435630 480
rect 435100 326 435630 354
rect 434414 -960 434526 326
rect 435518 -960 435630 326
rect 436714 -960 436826 480
rect 437492 354 437520 69838
rect 438872 16574 438900 75346
rect 447140 69828 447192 69834
rect 447140 69770 447192 69776
rect 440240 61396 440292 61402
rect 440240 61338 440292 61344
rect 438872 16546 439176 16574
rect 439148 480 439176 16546
rect 440252 3398 440280 61338
rect 444380 60172 444432 60178
rect 444380 60114 444432 60120
rect 441618 31104 441674 31113
rect 441618 31039 441674 31048
rect 441632 16574 441660 31039
rect 442998 21448 443054 21457
rect 442998 21383 443054 21392
rect 443012 16574 443040 21383
rect 444392 16574 444420 60114
rect 445760 17400 445812 17406
rect 445760 17342 445812 17348
rect 441632 16546 442672 16574
rect 443012 16546 443408 16574
rect 444392 16546 445064 16574
rect 440332 7676 440384 7682
rect 440332 7618 440384 7624
rect 440240 3392 440292 3398
rect 440240 3334 440292 3340
rect 440344 480 440372 7618
rect 441528 3392 441580 3398
rect 441528 3334 441580 3340
rect 441540 480 441568 3334
rect 442644 480 442672 16546
rect 437910 354 438022 480
rect 437492 326 438022 354
rect 437910 -960 438022 326
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443380 354 443408 16546
rect 445036 480 445064 16546
rect 443798 354 443910 480
rect 443380 326 443910 354
rect 443798 -960 443910 326
rect 444994 -960 445106 480
rect 445772 354 445800 17342
rect 447152 16574 447180 69770
rect 448520 54596 448572 54602
rect 448520 54538 448572 54544
rect 447152 16546 447456 16574
rect 447428 480 447456 16546
rect 448532 3210 448560 54538
rect 451280 53304 451332 53310
rect 451280 53246 451332 53252
rect 449900 20052 449952 20058
rect 449900 19994 449952 20000
rect 448612 17332 448664 17338
rect 448612 17274 448664 17280
rect 448624 3398 448652 17274
rect 449912 16574 449940 19994
rect 451292 16574 451320 53246
rect 456798 30968 456854 30977
rect 456798 30903 456854 30912
rect 455420 22908 455472 22914
rect 455420 22850 455472 22856
rect 454040 21480 454092 21486
rect 454040 21422 454092 21428
rect 449912 16546 450952 16574
rect 451292 16546 451688 16574
rect 448612 3392 448664 3398
rect 448612 3334 448664 3340
rect 449808 3392 449860 3398
rect 449808 3334 449860 3340
rect 448532 3182 448652 3210
rect 448624 480 448652 3182
rect 449820 480 449848 3334
rect 450924 480 450952 16546
rect 446190 354 446302 480
rect 445772 326 446302 354
rect 446190 -960 446302 326
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 451660 354 451688 16546
rect 453304 14544 453356 14550
rect 453304 14486 453356 14492
rect 453316 480 453344 14486
rect 452078 354 452190 480
rect 451660 326 452190 354
rect 452078 -960 452190 326
rect 453274 -960 453386 480
rect 454052 354 454080 21422
rect 455432 16574 455460 22850
rect 455432 16546 455736 16574
rect 455708 480 455736 16546
rect 456812 3210 456840 30903
rect 456892 20120 456944 20126
rect 456892 20062 456944 20068
rect 456904 3398 456932 20062
rect 459572 16574 459600 75375
rect 467840 68400 467892 68406
rect 467840 68342 467892 68348
rect 467852 16574 467880 68342
rect 480272 16574 480300 78134
rect 498200 78124 498252 78130
rect 498200 78066 498252 78072
rect 483018 77888 483074 77897
rect 483018 77823 483074 77832
rect 481640 62824 481692 62830
rect 481640 62766 481692 62772
rect 459572 16546 459968 16574
rect 467852 16546 468248 16574
rect 480272 16546 480576 16574
rect 459190 9208 459246 9217
rect 459190 9143 459246 9152
rect 456892 3392 456944 3398
rect 456892 3334 456944 3340
rect 458088 3392 458140 3398
rect 458088 3334 458140 3340
rect 456812 3182 456932 3210
rect 456904 480 456932 3182
rect 458100 480 458128 3334
rect 459204 480 459232 9143
rect 454470 354 454582 480
rect 454052 326 454582 354
rect 454470 -960 454582 326
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459940 354 459968 16546
rect 465172 9240 465224 9246
rect 465172 9182 465224 9188
rect 463976 9104 464028 9110
rect 463976 9046 464028 9052
rect 462780 6520 462832 6526
rect 462780 6462 462832 6468
rect 462226 4856 462282 4865
rect 462226 4791 462282 4800
rect 461584 3800 461636 3806
rect 461584 3742 461636 3748
rect 461596 480 461624 3742
rect 462240 3738 462268 4791
rect 462228 3732 462280 3738
rect 462228 3674 462280 3680
rect 462792 480 462820 6462
rect 463988 480 464016 9046
rect 465184 480 465212 9182
rect 467472 9036 467524 9042
rect 467472 8978 467524 8984
rect 466276 6452 466328 6458
rect 466276 6394 466328 6400
rect 466288 480 466316 6394
rect 467484 480 467512 8978
rect 460358 354 460470 480
rect 459940 326 460470 354
rect 460358 -960 460470 326
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468220 354 468248 16546
rect 474554 9072 474610 9081
rect 474554 9007 474610 9016
rect 469864 6384 469916 6390
rect 469864 6326 469916 6332
rect 469876 480 469904 6326
rect 471060 6316 471112 6322
rect 471060 6258 471112 6264
rect 471072 480 471100 6258
rect 473452 6248 473504 6254
rect 473452 6190 473504 6196
rect 472256 3664 472308 3670
rect 472256 3606 472308 3612
rect 472268 480 472296 3606
rect 473464 480 473492 6190
rect 474568 480 474596 9007
rect 478142 8936 478198 8945
rect 478142 8871 478198 8880
rect 476946 6352 477002 6361
rect 476946 6287 477002 6296
rect 475752 3596 475804 3602
rect 475752 3538 475804 3544
rect 475764 480 475792 3538
rect 476960 480 476988 6287
rect 478156 480 478184 8871
rect 479340 4888 479392 4894
rect 479340 4830 479392 4836
rect 479352 480 479380 4830
rect 480548 480 480576 16546
rect 481652 3602 481680 62766
rect 481732 60104 481784 60110
rect 481732 60046 481784 60052
rect 481640 3596 481692 3602
rect 481640 3538 481692 3544
rect 481744 480 481772 60046
rect 483032 16574 483060 77823
rect 489920 75336 489972 75342
rect 489920 75278 489972 75284
rect 496818 75304 496874 75313
rect 487160 54528 487212 54534
rect 487160 54470 487212 54476
rect 485780 44872 485832 44878
rect 485780 44814 485832 44820
rect 485792 16574 485820 44814
rect 483032 16546 484072 16574
rect 485792 16546 486464 16574
rect 482468 3596 482520 3602
rect 482468 3538 482520 3544
rect 468638 354 468750 480
rect 468220 326 468750 354
rect 468638 -960 468750 326
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482480 354 482508 3538
rect 484044 480 484072 16546
rect 484768 13116 484820 13122
rect 484768 13058 484820 13064
rect 482806 354 482918 480
rect 482480 326 482918 354
rect 482806 -960 482918 326
rect 484002 -960 484114 480
rect 484780 354 484808 13058
rect 486436 480 486464 16546
rect 485198 354 485310 480
rect 484780 326 485310 354
rect 485198 -960 485310 326
rect 486394 -960 486506 480
rect 487172 354 487200 54470
rect 488816 14476 488868 14482
rect 488816 14418 488868 14424
rect 488828 480 488856 14418
rect 489932 480 489960 75278
rect 496818 75239 496874 75248
rect 494058 53136 494114 53145
rect 494058 53071 494114 53080
rect 490012 35216 490064 35222
rect 490012 35158 490064 35164
rect 490024 16574 490052 35158
rect 494072 16574 494100 53071
rect 495438 43480 495494 43489
rect 495438 43415 495494 43424
rect 490024 16546 490696 16574
rect 494072 16546 494744 16574
rect 487590 354 487702 480
rect 487172 326 487702 354
rect 487590 -960 487702 326
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 490668 354 490696 16546
rect 492312 15904 492364 15910
rect 492312 15846 492364 15852
rect 492324 480 492352 15846
rect 493508 4820 493560 4826
rect 493508 4762 493560 4768
rect 493520 480 493548 4762
rect 494716 480 494744 16546
rect 491086 354 491198 480
rect 490668 326 491198 354
rect 491086 -960 491198 326
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495452 354 495480 43415
rect 496832 16574 496860 75239
rect 496832 16546 497136 16574
rect 497108 480 497136 16546
rect 498212 480 498240 78066
rect 527192 77246 527220 703520
rect 543476 700330 543504 703520
rect 559668 702434 559696 703520
rect 558932 702406 559696 702434
rect 543464 700324 543516 700330
rect 543464 700266 543516 700272
rect 558932 140078 558960 702406
rect 580262 697232 580318 697241
rect 580262 697167 580318 697176
rect 579618 683904 579674 683913
rect 579618 683839 579674 683848
rect 579632 683194 579660 683839
rect 579620 683188 579672 683194
rect 579620 683130 579672 683136
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 579986 617536 580042 617545
rect 579986 617471 580042 617480
rect 580000 616894 580028 617471
rect 579988 616888 580040 616894
rect 579988 616830 580040 616836
rect 579986 577688 580042 577697
rect 579986 577623 580042 577632
rect 580000 576910 580028 577623
rect 579988 576904 580040 576910
rect 579988 576846 580040 576852
rect 580170 564360 580226 564369
rect 580170 564295 580226 564304
rect 580184 563106 580212 564295
rect 580172 563100 580224 563106
rect 580172 563042 580224 563048
rect 579618 537840 579674 537849
rect 579618 537775 579674 537784
rect 579632 536858 579660 537775
rect 579620 536852 579672 536858
rect 579620 536794 579672 536800
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 579618 511320 579674 511329
rect 579618 511255 579674 511264
rect 579632 510678 579660 511255
rect 579620 510672 579672 510678
rect 579620 510614 579672 510620
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 579986 471472 580042 471481
rect 579986 471407 580042 471416
rect 580000 470626 580028 471407
rect 579988 470620 580040 470626
rect 579988 470562 580040 470568
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580184 456822 580212 458079
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 579710 418296 579766 418305
rect 579710 418231 579766 418240
rect 579724 418198 579752 418231
rect 579712 418192 579764 418198
rect 579712 418134 579764 418140
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580184 404394 580212 404903
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 580184 364410 580212 365055
rect 580172 364404 580224 364410
rect 580172 364346 580224 364352
rect 580172 351960 580224 351966
rect 580170 351928 580172 351937
rect 580224 351928 580226 351937
rect 580170 351863 580226 351872
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 580184 311914 580212 312015
rect 580172 311908 580224 311914
rect 580172 311850 580224 311856
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 580184 298178 580212 298687
rect 580172 298172 580224 298178
rect 580172 298114 580224 298120
rect 579618 272232 579674 272241
rect 579618 272167 579674 272176
rect 579632 271930 579660 272167
rect 579620 271924 579672 271930
rect 579620 271866 579672 271872
rect 580170 258904 580226 258913
rect 580170 258839 580226 258848
rect 580184 258126 580212 258839
rect 580172 258120 580224 258126
rect 580172 258062 580224 258068
rect 579618 245576 579674 245585
rect 579618 245511 579674 245520
rect 579632 244322 579660 245511
rect 579620 244316 579672 244322
rect 579620 244258 579672 244264
rect 579986 219056 580042 219065
rect 579986 218991 580042 219000
rect 580000 218074 580028 218991
rect 579988 218068 580040 218074
rect 579988 218010 580040 218016
rect 580170 205728 580226 205737
rect 580170 205663 580172 205672
rect 580224 205663 580226 205672
rect 580172 205634 580224 205640
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580184 178090 580212 179143
rect 580172 178084 580224 178090
rect 580172 178026 580224 178032
rect 579802 165880 579858 165889
rect 579802 165815 579858 165824
rect 579816 165646 579844 165815
rect 579804 165640 579856 165646
rect 579804 165582 579856 165588
rect 579986 152688 580042 152697
rect 579986 152623 580042 152632
rect 580000 151842 580028 152623
rect 579988 151836 580040 151842
rect 579988 151778 580040 151784
rect 558920 140072 558972 140078
rect 558920 140014 558972 140020
rect 580170 139360 580226 139369
rect 580170 139295 580226 139304
rect 580184 138038 580212 139295
rect 580172 138032 580224 138038
rect 580172 137974 580224 137980
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 580078 112840 580134 112849
rect 580078 112775 580134 112784
rect 580092 111858 580120 112775
rect 580080 111852 580132 111858
rect 580080 111794 580132 111800
rect 580078 99512 580134 99521
rect 580078 99447 580134 99456
rect 580092 99414 580120 99447
rect 580080 99408 580132 99414
rect 580080 99350 580132 99356
rect 580080 89412 580132 89418
rect 580080 89354 580132 89360
rect 574744 78056 574796 78062
rect 574744 77998 574796 78004
rect 527180 77240 527232 77246
rect 527180 77182 527232 77188
rect 557540 76628 557592 76634
rect 557540 76570 557592 76576
rect 506480 75268 506532 75274
rect 506480 75210 506532 75216
rect 500960 71188 501012 71194
rect 500960 71130 501012 71136
rect 498292 60036 498344 60042
rect 498292 59978 498344 59984
rect 498304 16574 498332 59978
rect 499580 22840 499632 22846
rect 499580 22782 499632 22788
rect 499592 16574 499620 22782
rect 500972 16574 501000 71130
rect 505100 57316 505152 57322
rect 505100 57258 505152 57264
rect 502340 47660 502392 47666
rect 502340 47602 502392 47608
rect 502352 16574 502380 47602
rect 505112 16574 505140 57258
rect 498304 16546 498976 16574
rect 499592 16546 500632 16574
rect 500972 16546 501368 16574
rect 502352 16546 503024 16574
rect 505112 16546 505416 16574
rect 495870 354 495982 480
rect 495452 326 495982 354
rect 495870 -960 495982 326
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 498948 354 498976 16546
rect 500604 480 500632 16546
rect 499366 354 499478 480
rect 498948 326 499478 354
rect 499366 -960 499478 326
rect 500562 -960 500674 480
rect 501340 354 501368 16546
rect 502996 480 503024 16546
rect 504180 7608 504232 7614
rect 504180 7550 504232 7556
rect 504192 480 504220 7550
rect 505388 480 505416 16546
rect 506492 3602 506520 75210
rect 517520 75200 517572 75206
rect 517520 75142 517572 75148
rect 549258 75168 549314 75177
rect 507860 71120 507912 71126
rect 507860 71062 507912 71068
rect 506572 17264 506624 17270
rect 506572 17206 506624 17212
rect 506480 3596 506532 3602
rect 506480 3538 506532 3544
rect 506584 3482 506612 17206
rect 507872 16574 507900 71062
rect 511998 64152 512054 64161
rect 511998 64087 512054 64096
rect 509240 18828 509292 18834
rect 509240 18770 509292 18776
rect 509252 16574 509280 18770
rect 507872 16546 508912 16574
rect 509252 16546 509648 16574
rect 507308 3596 507360 3602
rect 507308 3538 507360 3544
rect 506492 3454 506612 3482
rect 506492 480 506520 3454
rect 501758 354 501870 480
rect 501340 326 501870 354
rect 501758 -960 501870 326
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507320 354 507348 3538
rect 508884 480 508912 16546
rect 507646 354 507758 480
rect 507320 326 507758 354
rect 507646 -960 507758 326
rect 508842 -960 508954 480
rect 509620 354 509648 16546
rect 511262 14512 511318 14521
rect 511262 14447 511318 14456
rect 511276 480 511304 14447
rect 510038 354 510150 480
rect 509620 326 510150 354
rect 510038 -960 510150 326
rect 511234 -960 511346 480
rect 512012 354 512040 64087
rect 514758 50280 514814 50289
rect 514758 50215 514814 50224
rect 513378 21312 513434 21321
rect 513378 21247 513434 21256
rect 512430 354 512542 480
rect 512012 326 512542 354
rect 513392 354 513420 21247
rect 514772 480 514800 50215
rect 516140 49020 516192 49026
rect 516140 48962 516192 48968
rect 514852 21412 514904 21418
rect 514852 21354 514904 21360
rect 514864 16574 514892 21354
rect 516152 16574 516180 48962
rect 517532 16574 517560 75142
rect 549258 75103 549314 75112
rect 523040 71052 523092 71058
rect 523040 70994 523092 71000
rect 520280 50584 520332 50590
rect 520280 50526 520332 50532
rect 514864 16546 515536 16574
rect 516152 16546 517192 16574
rect 517532 16546 517928 16574
rect 513534 354 513646 480
rect 513392 326 513646 354
rect 512430 -960 512542 326
rect 513534 -960 513646 326
rect 514730 -960 514842 480
rect 515508 354 515536 16546
rect 517164 480 517192 16546
rect 515926 354 516038 480
rect 515508 326 516038 354
rect 515926 -960 516038 326
rect 517122 -960 517234 480
rect 517900 354 517928 16546
rect 519544 3528 519596 3534
rect 519544 3470 519596 3476
rect 519556 480 519584 3470
rect 518318 354 518430 480
rect 517900 326 518430 354
rect 518318 -960 518430 326
rect 519514 -960 519626 480
rect 520292 354 520320 50526
rect 521844 8968 521896 8974
rect 521844 8910 521896 8916
rect 521856 480 521884 8910
rect 523052 480 523080 70994
rect 536840 69760 536892 69766
rect 536840 69702 536892 69708
rect 529938 68232 529994 68241
rect 529938 68167 529994 68176
rect 527180 51808 527232 51814
rect 527180 51750 527232 51756
rect 523132 50516 523184 50522
rect 523132 50458 523184 50464
rect 523144 16574 523172 50458
rect 524420 26920 524472 26926
rect 524420 26862 524472 26868
rect 524432 16574 524460 26862
rect 527192 16574 527220 51750
rect 523144 16546 523816 16574
rect 524432 16546 525472 16574
rect 527192 16546 527864 16574
rect 520710 354 520822 480
rect 520292 326 520822 354
rect 520710 -960 520822 326
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 523788 354 523816 16546
rect 525444 480 525472 16546
rect 526628 3460 526680 3466
rect 526628 3402 526680 3408
rect 526640 480 526668 3402
rect 527836 480 527864 16546
rect 528558 13016 528614 13025
rect 528558 12951 528614 12960
rect 524206 354 524318 480
rect 523788 326 524318 354
rect 524206 -960 524318 326
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528572 354 528600 12951
rect 528990 354 529102 480
rect 528572 326 529102 354
rect 529952 354 529980 68167
rect 534080 51740 534132 51746
rect 534080 51682 534132 51688
rect 531318 28248 531374 28257
rect 531318 28183 531374 28192
rect 531332 3534 531360 28183
rect 531410 24168 531466 24177
rect 531410 24103 531466 24112
rect 531320 3528 531372 3534
rect 531320 3470 531372 3476
rect 531424 3346 531452 24103
rect 534092 16574 534120 51682
rect 535460 29640 535512 29646
rect 535460 29582 535512 29588
rect 535472 16574 535500 29582
rect 536852 16574 536880 69702
rect 539600 66972 539652 66978
rect 539600 66914 539652 66920
rect 538220 53236 538272 53242
rect 538220 53178 538272 53184
rect 534092 16546 534488 16574
rect 535472 16546 536144 16574
rect 536852 16546 537248 16574
rect 533710 3632 533766 3641
rect 533710 3567 533766 3576
rect 532148 3528 532200 3534
rect 532148 3470 532200 3476
rect 531332 3318 531452 3346
rect 531332 480 531360 3318
rect 530094 354 530206 480
rect 529952 326 530206 354
rect 528990 -960 529102 326
rect 530094 -960 530206 326
rect 531290 -960 531402 480
rect 532160 354 532188 3470
rect 533724 480 533752 3567
rect 532486 354 532598 480
rect 532160 326 532598 354
rect 532486 -960 532598 326
rect 533682 -960 533794 480
rect 534460 354 534488 16546
rect 536116 480 536144 16546
rect 537220 480 537248 16546
rect 534878 354 534990 480
rect 534460 326 534990 354
rect 534878 -960 534990 326
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538232 354 538260 53178
rect 539612 3534 539640 66914
rect 543740 66904 543792 66910
rect 543740 66846 543792 66852
rect 542360 31068 542412 31074
rect 542360 31010 542412 31016
rect 540980 25628 541032 25634
rect 540980 25570 541032 25576
rect 540992 16574 541020 25570
rect 542372 16574 542400 31010
rect 543752 16574 543780 66846
rect 547878 46200 547934 46209
rect 547878 46135 547934 46144
rect 546498 32600 546554 32609
rect 546498 32535 546554 32544
rect 545120 25560 545172 25566
rect 545120 25502 545172 25508
rect 545132 16574 545160 25502
rect 540992 16546 542032 16574
rect 542372 16546 542768 16574
rect 543752 16546 544424 16574
rect 545132 16546 545528 16574
rect 539692 10328 539744 10334
rect 539692 10270 539744 10276
rect 539600 3528 539652 3534
rect 539600 3470 539652 3476
rect 539704 3346 539732 10270
rect 540428 3528 540480 3534
rect 540428 3470 540480 3476
rect 539612 3318 539732 3346
rect 539612 480 539640 3318
rect 538374 354 538486 480
rect 538232 326 538486 354
rect 538374 -960 538486 326
rect 539570 -960 539682 480
rect 540440 354 540468 3470
rect 542004 480 542032 16546
rect 540766 354 540878 480
rect 540440 326 540878 354
rect 540766 -960 540878 326
rect 541962 -960 542074 480
rect 542740 354 542768 16546
rect 544396 480 544424 16546
rect 545500 480 545528 16546
rect 543158 354 543270 480
rect 542740 326 543270 354
rect 543158 -960 543270 326
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546512 354 546540 32535
rect 547892 480 547920 46135
rect 549272 16574 549300 75103
rect 552020 53168 552072 53174
rect 552020 53110 552072 53116
rect 550640 50448 550692 50454
rect 550640 50390 550692 50396
rect 550652 16574 550680 50390
rect 552032 16574 552060 53110
rect 556160 43444 556212 43450
rect 556160 43386 556212 43392
rect 553400 18760 553452 18766
rect 553400 18702 553452 18708
rect 553412 16574 553440 18702
rect 549272 16546 550312 16574
rect 550652 16546 551048 16574
rect 552032 16546 552704 16574
rect 553412 16546 553808 16574
rect 549074 6216 549130 6225
rect 549074 6151 549130 6160
rect 549088 480 549116 6151
rect 550284 480 550312 16546
rect 546654 354 546766 480
rect 546512 326 546766 354
rect 546654 -960 546766 326
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551020 354 551048 16546
rect 552676 480 552704 16546
rect 553780 480 553808 16546
rect 554962 3496 555018 3505
rect 554962 3431 555018 3440
rect 554976 480 555004 3431
rect 556172 480 556200 43386
rect 556252 18692 556304 18698
rect 556252 18634 556304 18640
rect 556264 16574 556292 18634
rect 557552 16574 557580 76570
rect 558920 76560 558972 76566
rect 558920 76502 558972 76508
rect 565818 76528 565874 76537
rect 558932 16574 558960 76502
rect 565818 76463 565874 76472
rect 564440 69692 564492 69698
rect 564440 69634 564492 69640
rect 561680 68332 561732 68338
rect 561680 68274 561732 68280
rect 560300 18624 560352 18630
rect 560300 18566 560352 18572
rect 560312 16574 560340 18566
rect 561692 16574 561720 68274
rect 563060 47592 563112 47598
rect 563060 47534 563112 47540
rect 556264 16546 556936 16574
rect 557552 16546 558592 16574
rect 558932 16546 559328 16574
rect 560312 16546 560432 16574
rect 561692 16546 562088 16574
rect 551438 354 551550 480
rect 551020 326 551550 354
rect 551438 -960 551550 326
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 556908 354 556936 16546
rect 558564 480 558592 16546
rect 557326 354 557438 480
rect 556908 326 557438 354
rect 557326 -960 557438 326
rect 558522 -960 558634 480
rect 559300 354 559328 16546
rect 559718 354 559830 480
rect 559300 326 559830 354
rect 560404 354 560432 16546
rect 562060 480 562088 16546
rect 560822 354 560934 480
rect 560404 326 560934 354
rect 559718 -960 559830 326
rect 560822 -960 560934 326
rect 562018 -960 562130 480
rect 563072 354 563100 47534
rect 564452 3534 564480 69634
rect 564532 57248 564584 57254
rect 564532 57190 564584 57196
rect 564440 3528 564492 3534
rect 564440 3470 564492 3476
rect 564544 3346 564572 57190
rect 565832 16574 565860 76463
rect 571340 53100 571392 53106
rect 571340 53042 571392 53048
rect 569960 50380 570012 50386
rect 569960 50322 570012 50328
rect 567198 32464 567254 32473
rect 567198 32399 567254 32408
rect 567212 16574 567240 32399
rect 569972 16574 570000 50322
rect 565832 16546 566872 16574
rect 567212 16546 567608 16574
rect 569972 16546 570368 16574
rect 565268 3528 565320 3534
rect 565268 3470 565320 3476
rect 564452 3318 564572 3346
rect 564452 480 564480 3318
rect 563214 354 563326 480
rect 563072 326 563326 354
rect 563214 -960 563326 326
rect 564410 -960 564522 480
rect 565280 354 565308 3470
rect 566844 480 566872 16546
rect 565606 354 565718 480
rect 565280 326 565718 354
rect 565606 -960 565718 326
rect 566802 -960 566914 480
rect 567580 354 567608 16546
rect 569130 3360 569186 3369
rect 569130 3295 569186 3304
rect 569144 480 569172 3295
rect 570340 480 570368 16546
rect 567998 354 568110 480
rect 567580 326 568110 354
rect 567998 -960 568110 326
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571352 354 571380 53042
rect 572720 33788 572772 33794
rect 572720 33730 572772 33736
rect 572732 16574 572760 33730
rect 572732 16546 573496 16574
rect 572720 6180 572772 6186
rect 572720 6122 572772 6128
rect 572732 480 572760 6122
rect 571494 354 571606 480
rect 571352 326 571606 354
rect 571494 -960 571606 326
rect 572690 -960 572802 480
rect 573468 354 573496 16546
rect 574652 11756 574704 11762
rect 574652 11698 574704 11704
rect 574664 3482 574692 11698
rect 574756 3602 574784 77998
rect 580092 77654 580120 89354
rect 580184 80617 580212 125967
rect 580170 80608 580226 80617
rect 580170 80543 580226 80552
rect 580276 79490 580304 697167
rect 580630 670712 580686 670721
rect 580630 670647 580686 670656
rect 580354 644056 580410 644065
rect 580354 643991 580410 644000
rect 580368 80578 580396 643991
rect 580446 591016 580502 591025
rect 580446 590951 580502 590960
rect 580460 80646 580488 590951
rect 580538 431624 580594 431633
rect 580538 431559 580594 431568
rect 580552 89418 580580 431559
rect 580644 429894 580672 670647
rect 580632 429888 580684 429894
rect 580632 429830 580684 429836
rect 580630 378448 580686 378457
rect 580630 378383 580686 378392
rect 580540 89412 580592 89418
rect 580540 89354 580592 89360
rect 580540 89276 580592 89282
rect 580540 89218 580592 89224
rect 580448 80640 580500 80646
rect 580448 80582 580500 80588
rect 580356 80572 580408 80578
rect 580356 80514 580408 80520
rect 580264 79484 580316 79490
rect 580264 79426 580316 79432
rect 580552 79354 580580 89218
rect 580644 79422 580672 378383
rect 580722 325272 580778 325281
rect 580722 325207 580778 325216
rect 580736 89282 580764 325207
rect 580814 232384 580870 232393
rect 580814 232319 580870 232328
rect 580724 89276 580776 89282
rect 580724 89218 580776 89224
rect 580828 89162 580856 232319
rect 580906 192536 580962 192545
rect 580906 192471 580962 192480
rect 580736 89134 580856 89162
rect 580736 80481 580764 89134
rect 580920 89026 580948 192471
rect 580828 88998 580948 89026
rect 580828 80714 580856 88998
rect 580906 86184 580962 86193
rect 580906 86119 580962 86128
rect 580920 80782 580948 86119
rect 580908 80776 580960 80782
rect 580908 80718 580960 80724
rect 580816 80708 580868 80714
rect 580816 80650 580868 80656
rect 580722 80472 580778 80481
rect 580722 80407 580778 80416
rect 580632 79416 580684 79422
rect 580632 79358 580684 79364
rect 580540 79348 580592 79354
rect 580540 79290 580592 79296
rect 581092 77988 581144 77994
rect 581092 77930 581144 77936
rect 580080 77648 580132 77654
rect 580080 77590 580132 77596
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 575478 62792 575534 62801
rect 575478 62727 575534 62736
rect 575492 16574 575520 62727
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 578238 58576 578294 58585
rect 578238 58511 578294 58520
rect 578252 16574 578280 58511
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 580170 33144 580226 33153
rect 580170 33079 580172 33088
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 579620 24132 579672 24138
rect 579620 24074 579672 24080
rect 579632 19825 579660 24074
rect 580264 22772 580316 22778
rect 580264 22714 580316 22720
rect 579618 19816 579674 19825
rect 579618 19751 579674 19760
rect 575492 16546 575888 16574
rect 578252 16546 578648 16574
rect 574744 3596 574796 3602
rect 574744 3538 574796 3544
rect 574664 3454 575152 3482
rect 575124 480 575152 3454
rect 573886 354 573998 480
rect 573468 326 573998 354
rect 573886 -960 573998 326
rect 575082 -960 575194 480
rect 575860 354 575888 16546
rect 577412 3732 577464 3738
rect 577412 3674 577464 3680
rect 577424 480 577452 3674
rect 578620 480 578648 16546
rect 580276 6633 580304 22714
rect 581104 16574 581132 77930
rect 582378 22672 582434 22681
rect 582378 22607 582434 22616
rect 582392 16574 582420 22607
rect 581104 16546 581776 16574
rect 582392 16546 583432 16574
rect 580262 6624 580318 6633
rect 580262 6559 580318 6568
rect 581000 3460 581052 3466
rect 581000 3402 581052 3408
rect 581012 480 581040 3402
rect 576278 354 576390 480
rect 575860 326 576390 354
rect 576278 -960 576390 326
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 581748 354 581776 16546
rect 583404 480 583432 16546
rect 582166 354 582278 480
rect 581748 326 582278 354
rect 582166 -960 582278 326
rect 583362 -960 583474 480
<< via2 >>
rect 2778 684256 2834 684312
rect 3514 671200 3570 671256
rect 3422 658144 3478 658200
rect 3330 632068 3332 632088
rect 3332 632068 3384 632088
rect 3384 632068 3386 632088
rect 3330 632032 3386 632068
rect 3146 579944 3202 580000
rect 3146 553832 3202 553888
rect 3330 527876 3386 527912
rect 3330 527856 3332 527876
rect 3332 527856 3384 527876
rect 3384 527856 3386 527876
rect 3330 514820 3386 514856
rect 3330 514800 3332 514820
rect 3332 514800 3384 514820
rect 3384 514800 3386 514820
rect 2778 501744 2834 501800
rect 3054 462576 3110 462632
rect 2962 449520 3018 449576
rect 3330 423544 3386 423600
rect 3330 397468 3332 397488
rect 3332 397468 3384 397488
rect 3384 397468 3386 397488
rect 3330 397432 3386 397468
rect 3330 371320 3386 371376
rect 3330 358400 3386 358456
rect 3330 345344 3386 345400
rect 3146 319232 3202 319288
rect 3330 306176 3386 306232
rect 3330 293120 3386 293176
rect 3238 267144 3294 267200
rect 2962 254088 3018 254144
rect 2870 227976 2926 228032
rect 3330 214920 3386 214976
rect 3330 201864 3386 201920
rect 3330 188808 3386 188864
rect 3330 175888 3386 175944
rect 3330 162868 3332 162888
rect 3332 162868 3384 162888
rect 3384 162868 3386 162888
rect 3330 162832 3386 162868
rect 2870 136720 2926 136776
rect 3330 110608 3386 110664
rect 3698 619112 3754 619168
rect 3606 606056 3662 606112
rect 3514 149776 3570 149832
rect 3514 97552 3570 97608
rect 3514 84632 3570 84688
rect 3422 78920 3478 78976
rect 3790 566888 3846 566944
rect 3882 475632 3938 475688
rect 3882 410488 3938 410544
rect 3974 241032 4030 241088
rect 4894 79192 4950 79248
rect 3606 79056 3662 79112
rect 1398 72392 1454 72448
rect 3422 71612 3424 71632
rect 3424 71612 3476 71632
rect 3476 71612 3478 71632
rect 3422 71576 3478 71612
rect 3054 58520 3110 58576
rect 3422 45500 3424 45520
rect 3424 45500 3476 45520
rect 3476 45500 3478 45520
rect 3422 45464 3478 45500
rect 3146 32408 3202 32464
rect 3330 19352 3386 19408
rect 3422 6432 3478 6488
rect 4066 4800 4122 4856
rect 117318 137536 117374 137592
rect 117318 136040 117374 136096
rect 117318 134544 117374 134600
rect 117410 133048 117466 133104
rect 117318 131552 117374 131608
rect 117318 130056 117374 130112
rect 117318 128560 117374 128616
rect 117318 127064 117374 127120
rect 117318 125568 117374 125624
rect 117318 124108 117320 124128
rect 117320 124108 117372 124128
rect 117372 124108 117374 124128
rect 117318 124072 117374 124108
rect 117318 122576 117374 122632
rect 117318 121080 117374 121136
rect 117318 119584 117374 119640
rect 117318 118088 117374 118144
rect 117318 116592 117374 116648
rect 117318 115096 117374 115152
rect 118054 113600 118110 113656
rect 118238 92656 118294 92712
rect 118146 91160 118202 91216
rect 118330 89664 118386 89720
rect 118882 107616 118938 107672
rect 119066 112104 119122 112160
rect 119158 110608 119214 110664
rect 119250 109112 119306 109168
rect 118974 106120 119030 106176
rect 118790 104624 118846 104680
rect 118698 103128 118754 103184
rect 118606 95648 118662 95704
rect 118514 94152 118570 94208
rect 118422 88168 118478 88224
rect 118422 86672 118478 86728
rect 118330 82184 118386 82240
rect 115202 79328 115258 79384
rect 10322 77832 10378 77888
rect 37278 76608 37334 76664
rect 20718 76472 20774 76528
rect 19338 25472 19394 25528
rect 22098 68176 22154 68232
rect 35898 73752 35954 73808
rect 40038 72528 40094 72584
rect 41878 7520 41934 7576
rect 55218 69536 55274 69592
rect 57978 68312 58034 68368
rect 57242 8880 57298 8936
rect 59634 9016 59690 9072
rect 75918 75112 75974 75168
rect 71778 73888 71834 73944
rect 73158 65456 73214 65512
rect 74538 44784 74594 44840
rect 91098 69672 91154 69728
rect 92754 9152 92810 9208
rect 109314 7656 109370 7712
rect 111798 76744 111854 76800
rect 110510 10240 110566 10296
rect 118606 85176 118662 85232
rect 118514 83680 118570 83736
rect 118422 80552 118478 80608
rect 120722 102040 120778 102096
rect 120814 100680 120870 100736
rect 120906 98640 120962 98696
rect 120998 97144 121054 97200
rect 143538 200640 143594 200696
rect 139398 195900 139454 195936
rect 139398 195880 139400 195900
rect 139400 195880 139452 195900
rect 139452 195880 139454 195900
rect 142342 195880 142398 195936
rect 153198 196152 153254 196208
rect 138110 195744 138166 195800
rect 140778 195744 140834 195800
rect 146206 195744 146262 195800
rect 148782 194656 148838 194712
rect 153474 195916 153476 195936
rect 153476 195916 153528 195936
rect 153528 195916 153530 195936
rect 153474 195880 153530 195916
rect 153934 195880 153990 195936
rect 157246 195880 157302 195936
rect 157154 195472 157210 195528
rect 158902 195880 158958 195936
rect 161386 195880 161442 195936
rect 159178 195744 159234 195800
rect 151450 193568 151506 193624
rect 153198 193568 153254 193624
rect 148782 190984 148838 191040
rect 149794 190576 149850 190632
rect 165434 196288 165490 196344
rect 144642 186904 144698 186960
rect 146114 180684 146116 180704
rect 146116 180684 146168 180704
rect 146168 180684 146170 180704
rect 146114 180648 146170 180684
rect 148046 179016 148102 179072
rect 142666 178744 142722 178800
rect 135258 173984 135314 174040
rect 137834 173984 137890 174040
rect 142066 176704 142122 176760
rect 144182 174528 144238 174584
rect 156050 174528 156106 174584
rect 145562 173848 145618 173904
rect 142710 173712 142766 173768
rect 142066 171128 142122 171184
rect 142066 170992 142122 171048
rect 142066 162152 142122 162208
rect 143538 142432 143594 142488
rect 142066 142160 142122 142216
rect 148690 173712 148746 173768
rect 146758 173576 146814 173632
rect 146482 143384 146538 143440
rect 148046 143248 148102 143304
rect 149610 143112 149666 143168
rect 151174 142976 151230 143032
rect 151358 142976 151414 143032
rect 151358 142568 151414 142624
rect 166170 196152 166226 196208
rect 166078 196016 166134 196072
rect 160558 142976 160614 143032
rect 164330 166368 164386 166424
rect 166998 166232 167054 166288
rect 171506 142840 171562 142896
rect 173070 142704 173126 142760
rect 179510 128152 179566 128208
rect 179602 126112 179658 126168
rect 179418 119312 179474 119368
rect 179694 116592 179750 116648
rect 179878 130464 179934 130520
rect 179786 112512 179842 112568
rect 123482 80144 123538 80200
rect 119342 79464 119398 79520
rect 122194 78240 122250 78296
rect 120722 75792 120778 75848
rect 122102 74432 122158 74488
rect 123850 76472 123906 76528
rect 125552 79906 125608 79962
rect 125736 79906 125792 79962
rect 125920 79906 125976 79962
rect 125874 79736 125930 79792
rect 125598 79636 125600 79656
rect 125600 79636 125652 79656
rect 125652 79636 125654 79656
rect 125598 79600 125654 79636
rect 125782 79600 125838 79656
rect 125690 78648 125746 78704
rect 125598 78512 125654 78568
rect 125966 78784 126022 78840
rect 125782 75792 125838 75848
rect 126748 79872 126804 79928
rect 126932 79906 126988 79962
rect 126058 77832 126114 77888
rect 126886 79736 126942 79792
rect 127392 79906 127448 79962
rect 127760 79906 127816 79962
rect 128036 79906 128092 79962
rect 127116 79736 127172 79792
rect 127714 79736 127770 79792
rect 127254 78648 127310 78704
rect 127346 78104 127402 78160
rect 127346 68176 127402 68232
rect 128312 79906 128368 79962
rect 128680 79872 128736 79928
rect 129048 79872 129104 79928
rect 128266 79600 128322 79656
rect 128450 77288 128506 77344
rect 129094 79736 129150 79792
rect 129508 79872 129564 79928
rect 128726 78104 128782 78160
rect 128542 76608 128598 76664
rect 128818 75928 128874 75984
rect 129692 79736 129748 79792
rect 129738 79600 129794 79656
rect 129968 79906 130024 79962
rect 130704 79906 130760 79962
rect 130106 79600 130162 79656
rect 129922 78648 129978 78704
rect 130198 78784 130254 78840
rect 130658 79636 130660 79656
rect 130660 79636 130712 79656
rect 130712 79636 130714 79656
rect 130980 79906 131036 79962
rect 131256 79872 131312 79928
rect 131440 79906 131496 79962
rect 130658 79600 130714 79636
rect 130290 76472 130346 76528
rect 130658 78784 130714 78840
rect 131118 79600 131174 79656
rect 131210 73888 131266 73944
rect 131808 79872 131864 79928
rect 131394 76608 131450 76664
rect 131578 79600 131634 79656
rect 131670 76608 131726 76664
rect 132360 79906 132416 79962
rect 132728 79872 132784 79928
rect 132636 79736 132692 79792
rect 133464 79872 133520 79928
rect 133648 79906 133704 79962
rect 133602 79600 133658 79656
rect 134016 79872 134072 79928
rect 134752 79906 134808 79962
rect 134246 76744 134302 76800
rect 134062 76608 134118 76664
rect 134798 79736 134854 79792
rect 135488 79906 135544 79962
rect 135672 79906 135728 79962
rect 134982 79600 135038 79656
rect 135626 79736 135682 79792
rect 135718 79600 135774 79656
rect 135902 78648 135958 78704
rect 136408 79872 136464 79928
rect 136776 79872 136832 79928
rect 136730 79736 136786 79792
rect 136960 79736 137016 79792
rect 136914 79600 136970 79656
rect 136914 76880 136970 76936
rect 137972 79872 138028 79928
rect 137880 79736 137936 79792
rect 137650 76472 137706 76528
rect 138616 79872 138672 79928
rect 138984 79906 139040 79962
rect 137926 76608 137982 76664
rect 138294 76472 138350 76528
rect 139628 79872 139684 79928
rect 138938 76608 138994 76664
rect 139122 76744 139178 76800
rect 139030 75792 139086 75848
rect 139214 75656 139270 75712
rect 140548 79872 140604 79928
rect 139950 79600 140006 79656
rect 140456 79736 140512 79792
rect 140824 79736 140880 79792
rect 140594 76608 140650 76664
rect 140686 74296 140742 74352
rect 141238 79600 141294 79656
rect 142112 79872 142168 79928
rect 142388 79906 142444 79962
rect 143124 79872 143180 79928
rect 142894 79736 142950 79792
rect 143492 79906 143548 79962
rect 144044 79906 144100 79962
rect 144504 79906 144560 79962
rect 142066 77152 142122 77208
rect 144780 79736 144836 79792
rect 143170 76608 143226 76664
rect 143262 76472 143318 76528
rect 143446 76608 143502 76664
rect 144458 79600 144514 79656
rect 144734 76744 144790 76800
rect 144550 76608 144606 76664
rect 144826 76472 144882 76528
rect 146160 79872 146216 79928
rect 146068 79736 146124 79792
rect 146620 79872 146676 79928
rect 146896 79872 146952 79928
rect 146712 79736 146768 79792
rect 147264 79872 147320 79928
rect 146298 76608 146354 76664
rect 146574 76744 146630 76800
rect 146482 76608 146538 76664
rect 146390 76472 146446 76528
rect 146298 76336 146354 76392
rect 147034 79600 147090 79656
rect 147034 77016 147090 77072
rect 147310 77832 147366 77888
rect 148092 79872 148148 79928
rect 147494 76880 147550 76936
rect 147402 74976 147458 75032
rect 147954 79600 148010 79656
rect 147862 74432 147918 74488
rect 148552 79872 148608 79928
rect 148920 79872 148976 79928
rect 149012 79736 149068 79792
rect 148506 74024 148562 74080
rect 149656 79872 149712 79928
rect 149610 79736 149666 79792
rect 148874 76608 148930 76664
rect 148966 73888 149022 73944
rect 148690 72392 148746 72448
rect 147126 3576 147182 3632
rect 150116 79872 150172 79928
rect 150300 79736 150356 79792
rect 150576 79838 150632 79894
rect 150162 75112 150218 75168
rect 150530 79600 150586 79656
rect 150346 73752 150402 73808
rect 151680 79872 151736 79928
rect 152048 79906 152104 79962
rect 152002 79736 152058 79792
rect 151542 78648 151598 78704
rect 151910 79620 151966 79656
rect 152416 79906 152472 79962
rect 151910 79600 151912 79620
rect 151912 79600 151964 79620
rect 151964 79600 151966 79620
rect 151726 78784 151782 78840
rect 151634 77560 151690 77616
rect 151726 77424 151782 77480
rect 152462 79600 152518 79656
rect 153060 79906 153116 79962
rect 152876 79736 152932 79792
rect 153244 79906 153300 79962
rect 153428 79906 153484 79962
rect 153198 77968 153254 78024
rect 153014 77288 153070 77344
rect 152462 43424 152518 43480
rect 153934 78104 153990 78160
rect 154348 79872 154404 79928
rect 154532 79736 154588 79792
rect 154486 79600 154542 79656
rect 154394 77832 154450 77888
rect 154670 79600 154726 79656
rect 154486 77560 154542 77616
rect 155268 79736 155324 79792
rect 155038 78648 155094 78704
rect 156418 79736 156474 79792
rect 155774 77288 155830 77344
rect 157108 79872 157164 79928
rect 156234 76744 156290 76800
rect 157200 79736 157256 79792
rect 157246 78784 157302 78840
rect 157154 77968 157210 78024
rect 158396 79906 158452 79962
rect 158304 79736 158360 79792
rect 159408 79906 159464 79962
rect 158442 77968 158498 78024
rect 158534 77832 158590 77888
rect 158718 77424 158774 77480
rect 159086 79736 159142 79792
rect 159270 79736 159326 79792
rect 158994 77968 159050 78024
rect 159178 77288 159234 77344
rect 159868 79906 159924 79962
rect 160512 79872 160568 79928
rect 159914 78648 159970 78704
rect 159914 78512 159970 78568
rect 159822 78104 159878 78160
rect 158902 6160 158958 6216
rect 156602 3440 156658 3496
rect 160006 78240 160062 78296
rect 160374 79736 160430 79792
rect 160098 76472 160154 76528
rect 160742 79736 160798 79792
rect 161248 79872 161304 79928
rect 160650 78512 160706 78568
rect 161110 76472 161166 76528
rect 161202 75384 161258 75440
rect 161984 79872 162040 79928
rect 162628 79872 162684 79928
rect 162122 76472 162178 76528
rect 162490 76472 162546 76528
rect 162996 79872 163052 79928
rect 162904 79736 162960 79792
rect 162674 77832 162730 77888
rect 162582 76336 162638 76392
rect 163134 78784 163190 78840
rect 163226 78240 163282 78296
rect 164008 79872 164064 79928
rect 164192 79872 164248 79928
rect 163502 76472 163558 76528
rect 164100 79736 164156 79792
rect 164054 74976 164110 75032
rect 165296 79872 165352 79928
rect 164882 79600 164938 79656
rect 164882 78376 164938 78432
rect 164974 77968 165030 78024
rect 164974 77560 165030 77616
rect 164882 77152 164938 77208
rect 164882 76200 164938 76256
rect 165158 79464 165214 79520
rect 165480 79736 165536 79792
rect 165756 79872 165812 79928
rect 165434 78648 165490 78704
rect 165342 76472 165398 76528
rect 165618 76336 165674 76392
rect 165894 79600 165950 79656
rect 161294 3304 161350 3360
rect 166768 79872 166824 79928
rect 166860 79736 166916 79792
rect 166722 76472 166778 76528
rect 167320 79872 167376 79928
rect 167688 79872 167744 79928
rect 166998 76336 167054 76392
rect 167182 79600 167238 79656
rect 167642 78512 167698 78568
rect 168056 79736 168112 79792
rect 168240 79872 168296 79928
rect 167826 76356 167882 76392
rect 167826 76336 167828 76356
rect 167828 76336 167880 76356
rect 167880 76336 167882 76356
rect 168102 79600 168158 79656
rect 168194 76472 168250 76528
rect 168792 79872 168848 79928
rect 168976 79872 169032 79928
rect 168746 79600 168802 79656
rect 168838 78648 168894 78704
rect 168654 78512 168710 78568
rect 168746 78376 168802 78432
rect 169712 79736 169768 79792
rect 170264 79872 170320 79928
rect 169666 76472 169722 76528
rect 169574 75112 169630 75168
rect 169850 77288 169906 77344
rect 169850 75928 169906 75984
rect 170908 79906 170964 79962
rect 171184 79906 171240 79962
rect 170816 79736 170872 79792
rect 170310 78648 170366 78704
rect 170494 77424 170550 77480
rect 170402 75928 170458 75984
rect 170678 78920 170734 78976
rect 170678 78648 170734 78704
rect 170954 78920 171010 78976
rect 170586 76064 170642 76120
rect 170954 77832 171010 77888
rect 171460 79906 171516 79962
rect 171736 79906 171792 79962
rect 172012 79906 172068 79962
rect 171414 78920 171470 78976
rect 171874 78784 171930 78840
rect 171782 78648 171838 78704
rect 171322 78376 171378 78432
rect 171506 78376 171562 78432
rect 171598 78240 171654 78296
rect 171230 78104 171286 78160
rect 171230 77832 171286 77888
rect 171230 77696 171286 77752
rect 172058 78240 172114 78296
rect 171598 77832 171654 77888
rect 172380 79906 172436 79962
rect 172242 77696 172298 77752
rect 172058 77560 172114 77616
rect 171966 75792 172022 75848
rect 172150 77152 172206 77208
rect 172150 74976 172206 75032
rect 172426 78920 172482 78976
rect 173208 79906 173264 79962
rect 172518 78784 172574 78840
rect 172978 79328 173034 79384
rect 173576 79872 173632 79928
rect 173346 79600 173402 79656
rect 173254 79464 173310 79520
rect 173346 79364 173348 79384
rect 173348 79364 173400 79384
rect 173400 79364 173402 79384
rect 173346 79328 173402 79364
rect 173070 79192 173126 79248
rect 173622 79464 173678 79520
rect 174036 79872 174092 79928
rect 173898 79600 173954 79656
rect 173162 76336 173218 76392
rect 172518 66952 172574 67008
rect 174542 79328 174598 79384
rect 178038 80144 178094 80200
rect 177394 79500 177396 79520
rect 177396 79500 177448 79520
rect 177448 79500 177450 79520
rect 177394 79464 177450 79500
rect 178590 78920 178646 78976
rect 179510 78920 179566 78976
rect 174542 78376 174598 78432
rect 179142 78104 179198 78160
rect 175922 76200 175978 76256
rect 174542 74296 174598 74352
rect 175278 69536 175334 69592
rect 176658 75656 176714 75712
rect 180062 80280 180118 80336
rect 180982 121488 181038 121544
rect 180890 117408 180946 117464
rect 181166 126928 181222 126984
rect 181258 114688 181314 114744
rect 181534 129648 181590 129704
rect 181442 120128 181498 120184
rect 181350 113328 181406 113384
rect 181074 109248 181130 109304
rect 182178 124208 182234 124264
rect 182178 98368 182234 98424
rect 182178 97008 182234 97064
rect 182454 122848 182510 122904
rect 182546 110608 182602 110664
rect 182638 101088 182694 101144
rect 182454 99728 182510 99784
rect 182822 92928 182878 92984
rect 182822 80688 182878 80744
rect 182362 78240 182418 78296
rect 176750 3848 176806 3904
rect 183282 107888 183338 107944
rect 183282 106528 183338 106584
rect 183282 105168 183338 105224
rect 183282 103808 183338 103864
rect 183466 102448 183522 102504
rect 183190 95648 183246 95704
rect 183466 94288 183522 94344
rect 183374 91568 183430 91624
rect 183466 90208 183522 90264
rect 183374 88848 183430 88904
rect 183466 87488 183522 87544
rect 183374 86128 183430 86184
rect 183466 84768 183522 84824
rect 183466 83408 183522 83464
rect 183006 82048 183062 82104
rect 193218 66816 193274 66872
rect 191838 47776 191894 47832
rect 193310 26968 193366 27024
rect 212538 17312 212594 17368
rect 230478 74160 230534 74216
rect 227718 61376 227774 61432
rect 226430 32680 226486 32736
rect 229374 13232 229430 13288
rect 247038 77016 247094 77072
rect 244278 74024 244334 74080
rect 245658 64232 245714 64288
rect 248418 20032 248474 20088
rect 266358 78920 266414 78976
rect 255962 77968 256018 78024
rect 263598 62872 263654 62928
rect 266358 51992 266414 52048
rect 264978 39208 265034 39264
rect 282918 76880 282974 76936
rect 279514 9560 279570 9616
rect 280710 9424 280766 9480
rect 281906 3712 281962 3768
rect 284390 73888 284446 73944
rect 298098 72392 298154 72448
rect 300858 17176 300914 17232
rect 299662 6568 299718 6624
rect 300766 6432 300822 6488
rect 354678 76744 354734 76800
rect 318798 73752 318854 73808
rect 316038 55936 316094 55992
rect 316130 42064 316186 42120
rect 317418 26832 317474 26888
rect 333978 51856 334034 51912
rect 336738 35264 336794 35320
rect 336278 11736 336334 11792
rect 353298 68312 353354 68368
rect 351918 47640 351974 47696
rect 350538 35128 350594 35184
rect 369858 51720 369914 51776
rect 372618 21528 372674 21584
rect 365810 15816 365866 15872
rect 371238 13096 371294 13152
rect 397458 78784 397514 78840
rect 389178 76608 389234 76664
rect 387798 55800 387854 55856
rect 402978 75520 403034 75576
rect 405738 47504 405794 47560
rect 407118 18536 407174 18592
rect 407210 9288 407266 9344
rect 423678 48864 423734 48920
rect 422298 19896 422354 19952
rect 420918 10240 420974 10296
rect 462318 78648 462374 78704
rect 423770 11600 423826 11656
rect 459558 75384 459614 75440
rect 441618 31048 441674 31104
rect 442998 21392 443054 21448
rect 456798 30912 456854 30968
rect 483018 77832 483074 77888
rect 459190 9152 459246 9208
rect 462226 4800 462282 4856
rect 474554 9016 474610 9072
rect 478142 8880 478198 8936
rect 476946 6296 477002 6352
rect 496818 75248 496874 75304
rect 494058 53080 494114 53136
rect 495438 43424 495494 43480
rect 580262 697176 580318 697232
rect 579618 683848 579674 683904
rect 580170 630808 580226 630864
rect 579986 617480 580042 617536
rect 579986 577632 580042 577688
rect 580170 564304 580226 564360
rect 579618 537784 579674 537840
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 579618 511264 579674 511320
rect 580170 484608 580226 484664
rect 579986 471416 580042 471472
rect 580170 458088 580226 458144
rect 579710 418240 579766 418296
rect 580170 404912 580226 404968
rect 580170 365064 580226 365120
rect 580170 351908 580172 351928
rect 580172 351908 580224 351928
rect 580224 351908 580226 351928
rect 580170 351872 580226 351908
rect 580170 312024 580226 312080
rect 580170 298696 580226 298752
rect 579618 272176 579674 272232
rect 580170 258848 580226 258904
rect 579618 245520 579674 245576
rect 579986 219000 580042 219056
rect 580170 205692 580226 205728
rect 580170 205672 580172 205692
rect 580172 205672 580224 205692
rect 580224 205672 580226 205692
rect 580170 179152 580226 179208
rect 579802 165824 579858 165880
rect 579986 152632 580042 152688
rect 580170 139304 580226 139360
rect 580170 125976 580226 126032
rect 580078 112784 580134 112840
rect 580078 99456 580134 99512
rect 511998 64096 512054 64152
rect 511262 14456 511318 14512
rect 514758 50224 514814 50280
rect 513378 21256 513434 21312
rect 549258 75112 549314 75168
rect 529938 68176 529994 68232
rect 528558 12960 528614 13016
rect 531318 28192 531374 28248
rect 531410 24112 531466 24168
rect 533710 3576 533766 3632
rect 547878 46144 547934 46200
rect 546498 32544 546554 32600
rect 549074 6160 549130 6216
rect 554962 3440 555018 3496
rect 565818 76472 565874 76528
rect 567198 32408 567254 32464
rect 569130 3304 569186 3360
rect 580170 80552 580226 80608
rect 580630 670656 580686 670712
rect 580354 644000 580410 644056
rect 580446 590960 580502 591016
rect 580538 431568 580594 431624
rect 580630 378392 580686 378448
rect 580722 325216 580778 325272
rect 580814 232328 580870 232384
rect 580906 192480 580962 192536
rect 580906 86128 580962 86184
rect 580722 80416 580778 80472
rect 580170 72936 580226 72992
rect 575478 62736 575534 62792
rect 580170 59608 580226 59664
rect 578238 58520 578294 58576
rect 580170 46280 580226 46336
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 579618 19760 579674 19816
rect 582378 22616 582434 22672
rect 580262 6568 580318 6624
<< metal3 >>
rect -960 697220 480 697460
rect 580257 697234 580323 697237
rect 583520 697234 584960 697324
rect 580257 697232 584960 697234
rect 580257 697176 580262 697232
rect 580318 697176 584960 697232
rect 580257 697174 584960 697176
rect 580257 697171 580323 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 2773 684314 2839 684317
rect -960 684312 2839 684314
rect -960 684256 2778 684312
rect 2834 684256 2839 684312
rect -960 684254 2839 684256
rect -960 684164 480 684254
rect 2773 684251 2839 684254
rect 579613 683906 579679 683909
rect 583520 683906 584960 683996
rect 579613 683904 584960 683906
rect 579613 683848 579618 683904
rect 579674 683848 584960 683904
rect 579613 683846 584960 683848
rect 579613 683843 579679 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580625 670714 580691 670717
rect 583520 670714 584960 670804
rect 580625 670712 584960 670714
rect 580625 670656 580630 670712
rect 580686 670656 584960 670712
rect 580625 670654 584960 670656
rect 580625 670651 580691 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580349 644058 580415 644061
rect 583520 644058 584960 644148
rect 580349 644056 584960 644058
rect 580349 644000 580354 644056
rect 580410 644000 584960 644056
rect 580349 643998 584960 644000
rect 580349 643995 580415 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3325 632090 3391 632093
rect -960 632088 3391 632090
rect -960 632032 3330 632088
rect 3386 632032 3391 632088
rect -960 632030 3391 632032
rect -960 631940 480 632030
rect 3325 632027 3391 632030
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3693 619170 3759 619173
rect -960 619168 3759 619170
rect -960 619112 3698 619168
rect 3754 619112 3759 619168
rect -960 619110 3759 619112
rect -960 619020 480 619110
rect 3693 619107 3759 619110
rect 579981 617538 580047 617541
rect 583520 617538 584960 617628
rect 579981 617536 584960 617538
rect 579981 617480 579986 617536
rect 580042 617480 584960 617536
rect 579981 617478 584960 617480
rect 579981 617475 580047 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3601 606114 3667 606117
rect -960 606112 3667 606114
rect -960 606056 3606 606112
rect 3662 606056 3667 606112
rect -960 606054 3667 606056
rect -960 605964 480 606054
rect 3601 606051 3667 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 580441 591018 580507 591021
rect 583520 591018 584960 591108
rect 580441 591016 584960 591018
rect 580441 590960 580446 591016
rect 580502 590960 584960 591016
rect 580441 590958 584960 590960
rect 580441 590955 580507 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3141 580002 3207 580005
rect -960 580000 3207 580002
rect -960 579944 3146 580000
rect 3202 579944 3207 580000
rect -960 579942 3207 579944
rect -960 579852 480 579942
rect 3141 579939 3207 579942
rect 579981 577690 580047 577693
rect 583520 577690 584960 577780
rect 579981 577688 584960 577690
rect 579981 577632 579986 577688
rect 580042 577632 584960 577688
rect 579981 577630 584960 577632
rect 579981 577627 580047 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3785 566946 3851 566949
rect -960 566944 3851 566946
rect -960 566888 3790 566944
rect 3846 566888 3851 566944
rect -960 566886 3851 566888
rect -960 566796 480 566886
rect 3785 566883 3851 566886
rect 580165 564362 580231 564365
rect 583520 564362 584960 564452
rect 580165 564360 584960 564362
rect 580165 564304 580170 564360
rect 580226 564304 584960 564360
rect 580165 564302 584960 564304
rect 580165 564299 580231 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3141 553890 3207 553893
rect -960 553888 3207 553890
rect -960 553832 3146 553888
rect 3202 553832 3207 553888
rect -960 553830 3207 553832
rect -960 553740 480 553830
rect 3141 553827 3207 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 579613 537842 579679 537845
rect 583520 537842 584960 537932
rect 579613 537840 584960 537842
rect 579613 537784 579618 537840
rect 579674 537784 584960 537840
rect 579613 537782 584960 537784
rect 579613 537779 579679 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 3325 527914 3391 527917
rect -960 527912 3391 527914
rect -960 527856 3330 527912
rect 3386 527856 3391 527912
rect -960 527854 3391 527856
rect -960 527764 480 527854
rect 3325 527851 3391 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3325 514858 3391 514861
rect -960 514856 3391 514858
rect -960 514800 3330 514856
rect 3386 514800 3391 514856
rect -960 514798 3391 514800
rect -960 514708 480 514798
rect 3325 514795 3391 514798
rect 579613 511322 579679 511325
rect 583520 511322 584960 511412
rect 579613 511320 584960 511322
rect 579613 511264 579618 511320
rect 579674 511264 584960 511320
rect 579613 511262 584960 511264
rect 579613 511259 579679 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 2773 501802 2839 501805
rect -960 501800 2839 501802
rect -960 501744 2778 501800
rect 2834 501744 2839 501800
rect -960 501742 2839 501744
rect -960 501652 480 501742
rect 2773 501739 2839 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3877 475690 3943 475693
rect -960 475688 3943 475690
rect -960 475632 3882 475688
rect 3938 475632 3943 475688
rect -960 475630 3943 475632
rect -960 475540 480 475630
rect 3877 475627 3943 475630
rect 579981 471474 580047 471477
rect 583520 471474 584960 471564
rect 579981 471472 584960 471474
rect 579981 471416 579986 471472
rect 580042 471416 584960 471472
rect 579981 471414 584960 471416
rect 579981 471411 580047 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3049 462634 3115 462637
rect -960 462632 3115 462634
rect -960 462576 3054 462632
rect 3110 462576 3115 462632
rect -960 462574 3115 462576
rect -960 462484 480 462574
rect 3049 462571 3115 462574
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 2957 449578 3023 449581
rect -960 449576 3023 449578
rect -960 449520 2962 449576
rect 3018 449520 3023 449576
rect -960 449518 3023 449520
rect -960 449428 480 449518
rect 2957 449515 3023 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 580533 431626 580599 431629
rect 583520 431626 584960 431716
rect 580533 431624 584960 431626
rect 580533 431568 580538 431624
rect 580594 431568 584960 431624
rect 580533 431566 584960 431568
rect 580533 431563 580599 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3325 423602 3391 423605
rect -960 423600 3391 423602
rect -960 423544 3330 423600
rect 3386 423544 3391 423600
rect -960 423542 3391 423544
rect -960 423452 480 423542
rect 3325 423539 3391 423542
rect 579705 418298 579771 418301
rect 583520 418298 584960 418388
rect 579705 418296 584960 418298
rect 579705 418240 579710 418296
rect 579766 418240 584960 418296
rect 579705 418238 584960 418240
rect 579705 418235 579771 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3877 410546 3943 410549
rect -960 410544 3943 410546
rect -960 410488 3882 410544
rect 3938 410488 3943 410544
rect -960 410486 3943 410488
rect -960 410396 480 410486
rect 3877 410483 3943 410486
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3325 397490 3391 397493
rect -960 397488 3391 397490
rect -960 397432 3330 397488
rect 3386 397432 3391 397488
rect -960 397430 3391 397432
rect -960 397340 480 397430
rect 3325 397427 3391 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580625 378450 580691 378453
rect 583520 378450 584960 378540
rect 580625 378448 584960 378450
rect 580625 378392 580630 378448
rect 580686 378392 584960 378448
rect 580625 378390 584960 378392
rect 580625 378387 580691 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 3325 371378 3391 371381
rect -960 371376 3391 371378
rect -960 371320 3330 371376
rect 3386 371320 3391 371376
rect -960 371318 3391 371320
rect -960 371228 480 371318
rect 3325 371315 3391 371318
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 3325 358458 3391 358461
rect -960 358456 3391 358458
rect -960 358400 3330 358456
rect 3386 358400 3391 358456
rect -960 358398 3391 358400
rect -960 358308 480 358398
rect 3325 358395 3391 358398
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 3325 345402 3391 345405
rect -960 345400 3391 345402
rect -960 345344 3330 345400
rect 3386 345344 3391 345400
rect -960 345342 3391 345344
rect -960 345252 480 345342
rect 3325 345339 3391 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 580717 325274 580783 325277
rect 583520 325274 584960 325364
rect 580717 325272 584960 325274
rect 580717 325216 580722 325272
rect 580778 325216 584960 325272
rect 580717 325214 584960 325216
rect 580717 325211 580783 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3141 319290 3207 319293
rect -960 319288 3207 319290
rect -960 319232 3146 319288
rect 3202 319232 3207 319288
rect -960 319230 3207 319232
rect -960 319140 480 319230
rect 3141 319227 3207 319230
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3325 306234 3391 306237
rect -960 306232 3391 306234
rect -960 306176 3330 306232
rect 3386 306176 3391 306232
rect -960 306174 3391 306176
rect -960 306084 480 306174
rect 3325 306171 3391 306174
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 3325 293178 3391 293181
rect -960 293176 3391 293178
rect -960 293120 3330 293176
rect 3386 293120 3391 293176
rect -960 293118 3391 293120
rect -960 293028 480 293118
rect 3325 293115 3391 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 579613 272234 579679 272237
rect 583520 272234 584960 272324
rect 579613 272232 584960 272234
rect 579613 272176 579618 272232
rect 579674 272176 584960 272232
rect 579613 272174 584960 272176
rect 579613 272171 579679 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 3233 267202 3299 267205
rect -960 267200 3299 267202
rect -960 267144 3238 267200
rect 3294 267144 3299 267200
rect -960 267142 3299 267144
rect -960 267052 480 267142
rect 3233 267139 3299 267142
rect 580165 258906 580231 258909
rect 583520 258906 584960 258996
rect 580165 258904 584960 258906
rect 580165 258848 580170 258904
rect 580226 258848 584960 258904
rect 580165 258846 584960 258848
rect 580165 258843 580231 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 2957 254146 3023 254149
rect -960 254144 3023 254146
rect -960 254088 2962 254144
rect 3018 254088 3023 254144
rect -960 254086 3023 254088
rect -960 253996 480 254086
rect 2957 254083 3023 254086
rect 579613 245578 579679 245581
rect 583520 245578 584960 245668
rect 579613 245576 584960 245578
rect 579613 245520 579618 245576
rect 579674 245520 584960 245576
rect 579613 245518 584960 245520
rect 579613 245515 579679 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 3969 241090 4035 241093
rect -960 241088 4035 241090
rect -960 241032 3974 241088
rect 4030 241032 4035 241088
rect -960 241030 4035 241032
rect -960 240940 480 241030
rect 3969 241027 4035 241030
rect 580809 232386 580875 232389
rect 583520 232386 584960 232476
rect 580809 232384 584960 232386
rect 580809 232328 580814 232384
rect 580870 232328 584960 232384
rect 580809 232326 584960 232328
rect 580809 232323 580875 232326
rect 583520 232236 584960 232326
rect -960 228034 480 228124
rect 2865 228034 2931 228037
rect -960 228032 2931 228034
rect -960 227976 2870 228032
rect 2926 227976 2931 228032
rect -960 227974 2931 227976
rect -960 227884 480 227974
rect 2865 227971 2931 227974
rect 579981 219058 580047 219061
rect 583520 219058 584960 219148
rect 579981 219056 584960 219058
rect 579981 219000 579986 219056
rect 580042 219000 584960 219056
rect 579981 218998 584960 219000
rect 579981 218995 580047 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 3325 214978 3391 214981
rect -960 214976 3391 214978
rect -960 214920 3330 214976
rect 3386 214920 3391 214976
rect -960 214918 3391 214920
rect -960 214828 480 214918
rect 3325 214915 3391 214918
rect 580165 205730 580231 205733
rect 583520 205730 584960 205820
rect 580165 205728 584960 205730
rect 580165 205672 580170 205728
rect 580226 205672 584960 205728
rect 580165 205670 584960 205672
rect 580165 205667 580231 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3325 201922 3391 201925
rect -960 201920 3391 201922
rect -960 201864 3330 201920
rect 3386 201864 3391 201920
rect -960 201862 3391 201864
rect -960 201772 480 201862
rect 3325 201859 3391 201862
rect 143533 200698 143599 200701
rect 144678 200698 144684 200700
rect 143533 200696 144684 200698
rect 143533 200640 143538 200696
rect 143594 200640 144684 200696
rect 143533 200638 144684 200640
rect 143533 200635 143599 200638
rect 144678 200636 144684 200638
rect 144748 200636 144754 200700
rect 149830 196284 149836 196348
rect 149900 196346 149906 196348
rect 165429 196346 165495 196349
rect 149900 196344 165495 196346
rect 149900 196288 165434 196344
rect 165490 196288 165495 196344
rect 149900 196286 165495 196288
rect 149900 196284 149906 196286
rect 165429 196283 165495 196286
rect 153193 196210 153259 196213
rect 166165 196210 166231 196213
rect 153193 196208 166231 196210
rect 153193 196152 153198 196208
rect 153254 196152 166170 196208
rect 166226 196152 166231 196208
rect 153193 196150 166231 196152
rect 153193 196147 153259 196150
rect 166165 196147 166231 196150
rect 151302 196012 151308 196076
rect 151372 196074 151378 196076
rect 166073 196074 166139 196077
rect 151372 196072 166139 196074
rect 151372 196016 166078 196072
rect 166134 196016 166139 196072
rect 151372 196014 166139 196016
rect 151372 196012 151378 196014
rect 166073 196011 166139 196014
rect 139393 195938 139459 195941
rect 142337 195938 142403 195941
rect 153469 195938 153535 195941
rect 139393 195936 142403 195938
rect 139393 195880 139398 195936
rect 139454 195880 142342 195936
rect 142398 195880 142403 195936
rect 139393 195878 142403 195880
rect 139393 195875 139459 195878
rect 142337 195875 142403 195878
rect 151126 195936 153535 195938
rect 151126 195880 153474 195936
rect 153530 195880 153535 195936
rect 151126 195878 153535 195880
rect 138105 195802 138171 195805
rect 140773 195802 140839 195805
rect 138105 195800 140839 195802
rect 138105 195744 138110 195800
rect 138166 195744 140778 195800
rect 140834 195744 140839 195800
rect 138105 195742 140839 195744
rect 138105 195739 138171 195742
rect 140773 195739 140839 195742
rect 146201 195802 146267 195805
rect 146201 195800 148426 195802
rect 146201 195744 146206 195800
rect 146262 195744 148426 195800
rect 146201 195742 148426 195744
rect 146201 195739 146267 195742
rect 148366 195712 148426 195742
rect 144678 195604 144684 195668
rect 144748 195604 144754 195668
rect 148366 195652 148948 195712
rect 151126 195696 151186 195878
rect 153469 195875 153535 195878
rect 153929 195938 153995 195941
rect 157241 195938 157307 195941
rect 153929 195936 157307 195938
rect 153929 195880 153934 195936
rect 153990 195880 157246 195936
rect 157302 195880 157307 195936
rect 153929 195878 157307 195880
rect 153929 195875 153995 195878
rect 157241 195875 157307 195878
rect 158897 195938 158963 195941
rect 161381 195938 161447 195941
rect 158897 195936 161447 195938
rect 158897 195880 158902 195936
rect 158958 195880 161386 195936
rect 161442 195880 161447 195936
rect 158897 195878 161447 195880
rect 158897 195875 158963 195878
rect 161381 195875 161447 195878
rect 159173 195802 159239 195805
rect 157750 195800 159239 195802
rect 157750 195744 159178 195800
rect 159234 195744 159239 195800
rect 157750 195742 159239 195744
rect 157750 195696 157810 195742
rect 159173 195739 159239 195742
rect 150604 195636 151186 195696
rect 157228 195636 157810 195696
rect 144686 195410 144746 195604
rect 157149 195530 157215 195533
rect 155910 195528 157215 195530
rect 155910 195472 157154 195528
rect 157210 195472 157215 195528
rect 155910 195470 157215 195472
rect 155910 195106 155970 195470
rect 157149 195467 157215 195470
rect 148777 194716 148843 194717
rect 148726 194714 148732 194716
rect 148686 194654 148732 194714
rect 148796 194712 148843 194716
rect 148838 194656 148843 194712
rect 148726 194652 148732 194654
rect 148796 194652 148843 194656
rect 148777 194651 148843 194652
rect 151445 193626 151511 193629
rect 153193 193626 153259 193629
rect 151445 193624 153259 193626
rect 151445 193568 151450 193624
rect 151506 193568 153198 193624
rect 153254 193568 153259 193624
rect 151445 193566 153259 193568
rect 151445 193563 151511 193566
rect 153193 193563 153259 193566
rect 580901 192538 580967 192541
rect 583520 192538 584960 192628
rect 580901 192536 584960 192538
rect 580901 192480 580906 192536
rect 580962 192480 584960 192536
rect 580901 192478 584960 192480
rect 580901 192475 580967 192478
rect 583520 192388 584960 192478
rect 143574 191744 143580 191808
rect 143644 191806 143650 191808
rect 143644 191746 143796 191806
rect 143644 191744 143650 191746
rect 143536 191336 144164 191396
rect 141734 191252 141740 191316
rect 141804 191314 141810 191316
rect 143536 191314 143596 191336
rect 151302 191316 151308 191318
rect 141804 191254 143596 191314
rect 151156 191256 151308 191316
rect 151302 191254 151308 191256
rect 151372 191254 151378 191318
rect 141804 191252 141810 191254
rect 141918 190572 141924 190636
rect 141988 190634 141994 190636
rect 144134 190634 144194 191226
rect 148777 191044 148843 191045
rect 148726 190980 148732 191044
rect 148796 191042 148843 191044
rect 148796 191040 148888 191042
rect 148838 190984 148888 191040
rect 148796 190982 148888 190984
rect 148796 190980 148843 190982
rect 148777 190979 148843 190980
rect 141988 190574 144194 190634
rect 149789 190636 149855 190637
rect 149789 190632 149836 190636
rect 149900 190634 149906 190636
rect 149789 190576 149794 190632
rect 141988 190572 141994 190574
rect 149789 190572 149836 190576
rect 149900 190574 149946 190634
rect 149900 190572 149906 190574
rect 149789 190571 149855 190572
rect -960 188866 480 188956
rect 3325 188866 3391 188869
rect -960 188864 3391 188866
rect -960 188808 3330 188864
rect 3386 188808 3391 188864
rect -960 188806 3391 188808
rect -960 188716 480 188806
rect 3325 188803 3391 188806
rect 140630 186900 140636 186964
rect 140700 186962 140706 186964
rect 144637 186962 144703 186965
rect 140700 186960 144703 186962
rect 140700 186904 144642 186960
rect 144698 186904 144703 186960
rect 140700 186902 144703 186904
rect 140700 186900 140706 186902
rect 144637 186899 144703 186902
rect 146109 180708 146175 180709
rect 146109 180704 146156 180708
rect 146220 180706 146226 180708
rect 146109 180648 146114 180704
rect 146109 180644 146156 180648
rect 146220 180646 146266 180706
rect 146220 180644 146226 180646
rect 146109 180643 146175 180644
rect 140446 179148 140452 179212
rect 140516 179210 140522 179212
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 140516 179150 148058 179210
rect 140516 179148 140522 179150
rect 147998 179077 148058 179150
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 147998 179072 148107 179077
rect 147998 179016 148046 179072
rect 148102 179016 148107 179072
rect 583520 179060 584960 179150
rect 147998 179014 148107 179016
rect 148041 179011 148107 179014
rect 142661 178804 142727 178805
rect 142654 178740 142660 178804
rect 142724 178802 142730 178804
rect 142724 178742 142816 178802
rect 142724 178740 142730 178742
rect 142661 178739 142727 178740
rect 142061 176762 142127 176765
rect 142654 176762 142660 176764
rect 142061 176760 142660 176762
rect 142061 176704 142066 176760
rect 142122 176704 142660 176760
rect 142061 176702 142660 176704
rect 142061 176699 142127 176702
rect 142654 176700 142660 176702
rect 142724 176700 142730 176764
rect -960 175946 480 176036
rect 3325 175946 3391 175949
rect -960 175944 3391 175946
rect -960 175888 3330 175944
rect 3386 175888 3391 175944
rect -960 175886 3391 175888
rect -960 175796 480 175886
rect 3325 175883 3391 175886
rect 144177 174586 144243 174589
rect 156045 174586 156111 174589
rect 144177 174584 156111 174586
rect 144177 174528 144182 174584
rect 144238 174528 156050 174584
rect 156106 174528 156111 174584
rect 144177 174526 156111 174528
rect 144177 174523 144243 174526
rect 156045 174523 156111 174526
rect 135253 174042 135319 174045
rect 137829 174042 137895 174045
rect 135253 174040 137895 174042
rect 135253 173984 135258 174040
rect 135314 173984 137834 174040
rect 137890 173984 137895 174040
rect 135253 173982 137895 173984
rect 135253 173979 135319 173982
rect 137829 173979 137895 173982
rect 142286 173844 142292 173908
rect 142356 173906 142362 173908
rect 145557 173906 145623 173909
rect 142356 173904 145623 173906
rect 142356 173848 145562 173904
rect 145618 173848 145623 173904
rect 142356 173846 145623 173848
rect 142356 173844 142362 173846
rect 145557 173843 145623 173846
rect 142705 173772 142771 173773
rect 142654 173770 142660 173772
rect 142614 173710 142660 173770
rect 142724 173768 142771 173772
rect 142766 173712 142771 173768
rect 142654 173708 142660 173710
rect 142724 173708 142771 173712
rect 144126 173708 144132 173772
rect 144196 173770 144202 173772
rect 148685 173770 148751 173773
rect 144196 173768 148751 173770
rect 144196 173712 148690 173768
rect 148746 173712 148751 173768
rect 144196 173710 148751 173712
rect 144196 173708 144202 173710
rect 142705 173707 142771 173708
rect 148685 173707 148751 173710
rect 142470 173572 142476 173636
rect 142540 173634 142546 173636
rect 146753 173634 146819 173637
rect 142540 173632 146819 173634
rect 142540 173576 146758 173632
rect 146814 173576 146819 173632
rect 142540 173574 146819 173576
rect 142540 173572 142546 173574
rect 146753 173571 146819 173574
rect 142102 171260 142108 171324
rect 142172 171260 142178 171324
rect 142110 171189 142170 171260
rect 142061 171186 142170 171189
rect 142016 171184 142170 171186
rect 142016 171128 142066 171184
rect 142122 171128 142170 171184
rect 142016 171126 142170 171128
rect 142061 171123 142127 171126
rect 142061 171050 142127 171053
rect 142016 171048 142170 171050
rect 142016 170992 142066 171048
rect 142122 170992 142170 171048
rect 142016 170990 142170 170992
rect 142061 170987 142170 170990
rect 142110 170916 142170 170987
rect 142102 170852 142108 170916
rect 142172 170852 142178 170916
rect 141734 166364 141740 166428
rect 141804 166426 141810 166428
rect 164325 166426 164391 166429
rect 141804 166424 164391 166426
rect 141804 166368 164330 166424
rect 164386 166368 164391 166424
rect 141804 166366 164391 166368
rect 141804 166364 141810 166366
rect 164325 166363 164391 166366
rect 141918 166228 141924 166292
rect 141988 166290 141994 166292
rect 166993 166290 167059 166293
rect 141988 166288 167059 166290
rect 141988 166232 166998 166288
rect 167054 166232 167059 166288
rect 141988 166230 167059 166232
rect 141988 166228 141994 166230
rect 166993 166227 167059 166230
rect 579797 165882 579863 165885
rect 583520 165882 584960 165972
rect 579797 165880 584960 165882
rect 579797 165824 579802 165880
rect 579858 165824 584960 165880
rect 579797 165822 584960 165824
rect 579797 165819 579863 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3325 162890 3391 162893
rect -960 162888 3391 162890
rect -960 162832 3330 162888
rect 3386 162832 3391 162888
rect -960 162830 3391 162832
rect -960 162740 480 162830
rect 3325 162827 3391 162830
rect 142061 162212 142127 162213
rect 142061 162210 142108 162212
rect 142016 162208 142108 162210
rect 142172 162210 142178 162212
rect 142016 162152 142066 162208
rect 142016 162150 142108 162152
rect 142061 162148 142108 162150
rect 142172 162150 142254 162210
rect 142172 162148 142178 162150
rect 142061 162147 142127 162148
rect 579981 152690 580047 152693
rect 583520 152690 584960 152780
rect 579981 152688 584960 152690
rect 579981 152632 579986 152688
rect 580042 152632 584960 152688
rect 579981 152630 584960 152632
rect 579981 152627 580047 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3509 149834 3575 149837
rect -960 149832 3575 149834
rect -960 149776 3514 149832
rect 3570 149776 3575 149832
rect -960 149774 3575 149776
rect -960 149684 480 149774
rect 3509 149771 3575 149774
rect 142286 143380 142292 143444
rect 142356 143442 142362 143444
rect 146477 143442 146543 143445
rect 142356 143440 146543 143442
rect 142356 143384 146482 143440
rect 146538 143384 146543 143440
rect 142356 143382 146543 143384
rect 142356 143380 142362 143382
rect 146477 143379 146543 143382
rect 142470 143244 142476 143308
rect 142540 143306 142546 143308
rect 148041 143306 148107 143309
rect 142540 143304 148107 143306
rect 142540 143248 148046 143304
rect 148102 143248 148107 143304
rect 142540 143246 148107 143248
rect 142540 143244 142546 143246
rect 148041 143243 148107 143246
rect 140446 143108 140452 143172
rect 140516 143170 140522 143172
rect 149605 143170 149671 143173
rect 140516 143168 149671 143170
rect 140516 143112 149610 143168
rect 149666 143112 149671 143168
rect 140516 143110 149671 143112
rect 140516 143108 140522 143110
rect 149605 143107 149671 143110
rect 144126 142972 144132 143036
rect 144196 143034 144202 143036
rect 151169 143034 151235 143037
rect 144196 143032 151235 143034
rect 144196 142976 151174 143032
rect 151230 142976 151235 143032
rect 144196 142974 151235 142976
rect 144196 142972 144202 142974
rect 151169 142971 151235 142974
rect 151353 143034 151419 143037
rect 160553 143034 160619 143037
rect 151353 143032 160619 143034
rect 151353 142976 151358 143032
rect 151414 142976 160558 143032
rect 160614 142976 160619 143032
rect 151353 142974 160619 142976
rect 151353 142971 151419 142974
rect 160553 142971 160619 142974
rect 146150 142836 146156 142900
rect 146220 142898 146226 142900
rect 171501 142898 171567 142901
rect 146220 142896 171567 142898
rect 146220 142840 171506 142896
rect 171562 142840 171567 142896
rect 146220 142838 171567 142840
rect 146220 142836 146226 142838
rect 171501 142835 171567 142838
rect 140630 142700 140636 142764
rect 140700 142762 140706 142764
rect 173065 142762 173131 142765
rect 140700 142760 173131 142762
rect 140700 142704 173070 142760
rect 173126 142704 173131 142760
rect 140700 142702 173131 142704
rect 140700 142700 140706 142702
rect 173065 142699 173131 142702
rect 143574 142564 143580 142628
rect 143644 142626 143650 142628
rect 151353 142626 151419 142629
rect 143644 142624 151419 142626
rect 143644 142568 151358 142624
rect 151414 142568 151419 142624
rect 143644 142566 151419 142568
rect 143644 142564 143650 142566
rect 151353 142563 151419 142566
rect 142102 142428 142108 142492
rect 142172 142490 142178 142492
rect 143533 142490 143599 142493
rect 142172 142488 143599 142490
rect 142172 142432 143538 142488
rect 143594 142432 143599 142488
rect 142172 142430 143599 142432
rect 142172 142428 142178 142430
rect 143533 142427 143599 142430
rect 142061 142218 142127 142221
rect 142654 142218 142660 142220
rect 142061 142216 142660 142218
rect 142061 142160 142066 142216
rect 142122 142160 142660 142216
rect 142061 142158 142660 142160
rect 142061 142155 142127 142158
rect 142654 142156 142660 142158
rect 142724 142156 142730 142220
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect 117313 137594 117379 137597
rect 117313 137592 120060 137594
rect 117313 137536 117318 137592
rect 117374 137536 120060 137592
rect 117313 137534 120060 137536
rect 117313 137531 117379 137534
rect -960 136778 480 136868
rect 2865 136778 2931 136781
rect -960 136776 2931 136778
rect -960 136720 2870 136776
rect 2926 136720 2931 136776
rect -960 136718 2931 136720
rect -960 136628 480 136718
rect 2865 136715 2931 136718
rect 117313 136098 117379 136101
rect 117313 136096 120060 136098
rect 117313 136040 117318 136096
rect 117374 136040 120060 136096
rect 117313 136038 120060 136040
rect 117313 136035 117379 136038
rect 117313 134602 117379 134605
rect 117313 134600 120060 134602
rect 117313 134544 117318 134600
rect 117374 134544 120060 134600
rect 117313 134542 120060 134544
rect 117313 134539 117379 134542
rect 117405 133106 117471 133109
rect 117405 133104 120060 133106
rect 117405 133048 117410 133104
rect 117466 133048 120060 133104
rect 117405 133046 120060 133048
rect 117405 133043 117471 133046
rect 117313 131610 117379 131613
rect 117313 131608 120060 131610
rect 117313 131552 117318 131608
rect 117374 131552 120060 131608
rect 117313 131550 120060 131552
rect 117313 131547 117379 131550
rect 179830 130525 179890 131036
rect 179830 130520 179939 130525
rect 179830 130464 179878 130520
rect 179934 130464 179939 130520
rect 179830 130462 179939 130464
rect 179873 130459 179939 130462
rect 117313 130114 117379 130117
rect 117313 130112 120060 130114
rect 117313 130056 117318 130112
rect 117374 130056 120060 130112
rect 117313 130054 120060 130056
rect 117313 130051 117379 130054
rect 181529 129706 181595 129709
rect 179860 129704 181595 129706
rect 179860 129648 181534 129704
rect 181590 129648 181595 129704
rect 179860 129646 181595 129648
rect 181529 129643 181595 129646
rect 117313 128618 117379 128621
rect 117313 128616 120060 128618
rect 117313 128560 117318 128616
rect 117374 128560 120060 128616
rect 117313 128558 120060 128560
rect 117313 128555 117379 128558
rect 179462 128213 179522 128316
rect 179462 128208 179571 128213
rect 179462 128152 179510 128208
rect 179566 128152 179571 128208
rect 179462 128150 179571 128152
rect 179505 128147 179571 128150
rect 117313 127122 117379 127125
rect 117313 127120 120060 127122
rect 117313 127064 117318 127120
rect 117374 127064 120060 127120
rect 117313 127062 120060 127064
rect 117313 127059 117379 127062
rect 181161 126986 181227 126989
rect 179860 126984 181227 126986
rect 179860 126928 181166 126984
rect 181222 126928 181227 126984
rect 179860 126926 181227 126928
rect 181161 126923 181227 126926
rect 179597 126170 179663 126173
rect 179597 126168 179706 126170
rect 179597 126112 179602 126168
rect 179658 126112 179706 126168
rect 179597 126107 179706 126112
rect 117313 125626 117379 125629
rect 117313 125624 120060 125626
rect 117313 125568 117318 125624
rect 117374 125568 120060 125624
rect 179646 125596 179706 126107
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect 117313 125566 120060 125568
rect 117313 125563 117379 125566
rect 182173 124266 182239 124269
rect 179860 124264 182239 124266
rect 179860 124208 182178 124264
rect 182234 124208 182239 124264
rect 179860 124206 182239 124208
rect 182173 124203 182239 124206
rect 117313 124130 117379 124133
rect 117313 124128 120060 124130
rect 117313 124072 117318 124128
rect 117374 124072 120060 124128
rect 117313 124070 120060 124072
rect 117313 124067 117379 124070
rect -960 123572 480 123812
rect 182449 122906 182515 122909
rect 179860 122904 182515 122906
rect 179860 122848 182454 122904
rect 182510 122848 182515 122904
rect 179860 122846 182515 122848
rect 182449 122843 182515 122846
rect 117313 122634 117379 122637
rect 117313 122632 120060 122634
rect 117313 122576 117318 122632
rect 117374 122576 120060 122632
rect 117313 122574 120060 122576
rect 117313 122571 117379 122574
rect 180977 121546 181043 121549
rect 179860 121544 181043 121546
rect 179860 121488 180982 121544
rect 181038 121488 181043 121544
rect 179860 121486 181043 121488
rect 180977 121483 181043 121486
rect 117313 121138 117379 121141
rect 117313 121136 120060 121138
rect 117313 121080 117318 121136
rect 117374 121080 120060 121136
rect 117313 121078 120060 121080
rect 117313 121075 117379 121078
rect 181437 120186 181503 120189
rect 179860 120184 181503 120186
rect 179860 120128 181442 120184
rect 181498 120128 181503 120184
rect 179860 120126 181503 120128
rect 181437 120123 181503 120126
rect 117313 119642 117379 119645
rect 117313 119640 120060 119642
rect 117313 119584 117318 119640
rect 117374 119584 120060 119640
rect 117313 119582 120060 119584
rect 117313 119579 117379 119582
rect 179413 119370 179479 119373
rect 179413 119368 179522 119370
rect 179413 119312 179418 119368
rect 179474 119312 179522 119368
rect 179413 119307 179522 119312
rect 179462 118796 179522 119307
rect 117313 118146 117379 118149
rect 117313 118144 120060 118146
rect 117313 118088 117318 118144
rect 117374 118088 120060 118144
rect 117313 118086 120060 118088
rect 117313 118083 117379 118086
rect 180885 117466 180951 117469
rect 179860 117464 180951 117466
rect 179860 117408 180890 117464
rect 180946 117408 180951 117464
rect 179860 117406 180951 117408
rect 180885 117403 180951 117406
rect 117313 116650 117379 116653
rect 179689 116650 179755 116653
rect 117313 116648 120060 116650
rect 117313 116592 117318 116648
rect 117374 116592 120060 116648
rect 117313 116590 120060 116592
rect 179646 116648 179755 116650
rect 179646 116592 179694 116648
rect 179750 116592 179755 116648
rect 117313 116587 117379 116590
rect 179646 116587 179755 116592
rect 179646 116076 179706 116587
rect 117313 115154 117379 115157
rect 117313 115152 120060 115154
rect 117313 115096 117318 115152
rect 117374 115096 120060 115152
rect 117313 115094 120060 115096
rect 117313 115091 117379 115094
rect 181253 114746 181319 114749
rect 179860 114744 181319 114746
rect 179860 114688 181258 114744
rect 181314 114688 181319 114744
rect 179860 114686 181319 114688
rect 181253 114683 181319 114686
rect 118049 113658 118115 113661
rect 118049 113656 120060 113658
rect 118049 113600 118054 113656
rect 118110 113600 120060 113656
rect 118049 113598 120060 113600
rect 118049 113595 118115 113598
rect 181345 113386 181411 113389
rect 179860 113384 181411 113386
rect 179860 113328 181350 113384
rect 181406 113328 181411 113384
rect 179860 113326 181411 113328
rect 181345 113323 181411 113326
rect 580073 112842 580139 112845
rect 583520 112842 584960 112932
rect 580073 112840 584960 112842
rect 580073 112784 580078 112840
rect 580134 112784 584960 112840
rect 580073 112782 584960 112784
rect 580073 112779 580139 112782
rect 583520 112692 584960 112782
rect 179781 112570 179847 112573
rect 179781 112568 179890 112570
rect 179781 112512 179786 112568
rect 179842 112512 179890 112568
rect 179781 112507 179890 112512
rect 119061 112162 119127 112165
rect 119061 112160 120060 112162
rect 119061 112104 119066 112160
rect 119122 112104 120060 112160
rect 119061 112102 120060 112104
rect 119061 112099 119127 112102
rect 179830 111996 179890 112507
rect -960 110666 480 110756
rect 3325 110666 3391 110669
rect -960 110664 3391 110666
rect -960 110608 3330 110664
rect 3386 110608 3391 110664
rect -960 110606 3391 110608
rect -960 110516 480 110606
rect 3325 110603 3391 110606
rect 119153 110666 119219 110669
rect 182541 110666 182607 110669
rect 119153 110664 120060 110666
rect 119153 110608 119158 110664
rect 119214 110608 120060 110664
rect 119153 110606 120060 110608
rect 179860 110664 182607 110666
rect 179860 110608 182546 110664
rect 182602 110608 182607 110664
rect 179860 110606 182607 110608
rect 119153 110603 119219 110606
rect 182541 110603 182607 110606
rect 181069 109306 181135 109309
rect 179860 109304 181135 109306
rect 179860 109248 181074 109304
rect 181130 109248 181135 109304
rect 179860 109246 181135 109248
rect 181069 109243 181135 109246
rect 119245 109170 119311 109173
rect 119245 109168 120060 109170
rect 119245 109112 119250 109168
rect 119306 109112 120060 109168
rect 119245 109110 120060 109112
rect 119245 109107 119311 109110
rect 183277 107946 183343 107949
rect 179860 107944 183343 107946
rect 179860 107888 183282 107944
rect 183338 107888 183343 107944
rect 179860 107886 183343 107888
rect 183277 107883 183343 107886
rect 118877 107674 118943 107677
rect 118877 107672 120060 107674
rect 118877 107616 118882 107672
rect 118938 107616 120060 107672
rect 118877 107614 120060 107616
rect 118877 107611 118943 107614
rect 183277 106586 183343 106589
rect 179860 106584 183343 106586
rect 179860 106528 183282 106584
rect 183338 106528 183343 106584
rect 179860 106526 183343 106528
rect 183277 106523 183343 106526
rect 118969 106178 119035 106181
rect 118969 106176 120060 106178
rect 118969 106120 118974 106176
rect 119030 106120 120060 106176
rect 118969 106118 120060 106120
rect 118969 106115 119035 106118
rect 183277 105226 183343 105229
rect 179860 105224 183343 105226
rect 179860 105168 183282 105224
rect 183338 105168 183343 105224
rect 179860 105166 183343 105168
rect 183277 105163 183343 105166
rect 118785 104682 118851 104685
rect 118785 104680 120060 104682
rect 118785 104624 118790 104680
rect 118846 104624 120060 104680
rect 118785 104622 120060 104624
rect 118785 104619 118851 104622
rect 183277 103866 183343 103869
rect 179860 103864 183343 103866
rect 179860 103808 183282 103864
rect 183338 103808 183343 103864
rect 179860 103806 183343 103808
rect 183277 103803 183343 103806
rect 118693 103186 118759 103189
rect 118693 103184 120060 103186
rect 118693 103128 118698 103184
rect 118754 103128 120060 103184
rect 118693 103126 120060 103128
rect 118693 103123 118759 103126
rect 183461 102506 183527 102509
rect 179860 102504 183527 102506
rect 179860 102448 183466 102504
rect 183522 102448 183527 102504
rect 179860 102446 183527 102448
rect 183461 102443 183527 102446
rect 120717 102098 120783 102101
rect 120582 102096 120783 102098
rect 120582 102040 120722 102096
rect 120778 102040 120783 102096
rect 120582 102038 120783 102040
rect 120582 101660 120642 102038
rect 120717 102035 120783 102038
rect 182633 101146 182699 101149
rect 179860 101144 182699 101146
rect 179860 101088 182638 101144
rect 182694 101088 182699 101144
rect 179860 101086 182699 101088
rect 182633 101083 182699 101086
rect 120809 100738 120875 100741
rect 120582 100736 120875 100738
rect 120582 100680 120814 100736
rect 120870 100680 120875 100736
rect 120582 100678 120875 100680
rect 120582 100164 120642 100678
rect 120809 100675 120875 100678
rect 182449 99786 182515 99789
rect 179860 99784 182515 99786
rect 179860 99728 182454 99784
rect 182510 99728 182515 99784
rect 179860 99726 182515 99728
rect 182449 99723 182515 99726
rect 580073 99514 580139 99517
rect 583520 99514 584960 99604
rect 580073 99512 584960 99514
rect 580073 99456 580078 99512
rect 580134 99456 584960 99512
rect 580073 99454 584960 99456
rect 580073 99451 580139 99454
rect 583520 99364 584960 99454
rect 120901 98698 120967 98701
rect 120612 98696 120967 98698
rect 120612 98640 120906 98696
rect 120962 98640 120967 98696
rect 120612 98638 120967 98640
rect 120901 98635 120967 98638
rect 182173 98426 182239 98429
rect 179860 98424 182239 98426
rect 179860 98368 182178 98424
rect 182234 98368 182239 98424
rect 179860 98366 182239 98368
rect 182173 98363 182239 98366
rect -960 97610 480 97700
rect 3509 97610 3575 97613
rect -960 97608 3575 97610
rect -960 97552 3514 97608
rect 3570 97552 3575 97608
rect -960 97550 3575 97552
rect -960 97460 480 97550
rect 3509 97547 3575 97550
rect 120993 97202 121059 97205
rect 120612 97200 121059 97202
rect 120612 97144 120998 97200
rect 121054 97144 121059 97200
rect 120612 97142 121059 97144
rect 120993 97139 121059 97142
rect 182173 97066 182239 97069
rect 179860 97064 182239 97066
rect 179860 97008 182178 97064
rect 182234 97008 182239 97064
rect 179860 97006 182239 97008
rect 182173 97003 182239 97006
rect 118601 95706 118667 95709
rect 183185 95706 183251 95709
rect 118601 95704 120060 95706
rect 118601 95648 118606 95704
rect 118662 95648 120060 95704
rect 118601 95646 120060 95648
rect 179860 95704 183251 95706
rect 179860 95648 183190 95704
rect 183246 95648 183251 95704
rect 179860 95646 183251 95648
rect 118601 95643 118667 95646
rect 183185 95643 183251 95646
rect 183461 94346 183527 94349
rect 179860 94344 183527 94346
rect 179860 94288 183466 94344
rect 183522 94288 183527 94344
rect 179860 94286 183527 94288
rect 183461 94283 183527 94286
rect 118509 94210 118575 94213
rect 118509 94208 120060 94210
rect 118509 94152 118514 94208
rect 118570 94152 120060 94208
rect 118509 94150 120060 94152
rect 118509 94147 118575 94150
rect 182817 92986 182883 92989
rect 179860 92984 182883 92986
rect 179860 92928 182822 92984
rect 182878 92928 182883 92984
rect 179860 92926 182883 92928
rect 182817 92923 182883 92926
rect 118233 92714 118299 92717
rect 118233 92712 120060 92714
rect 118233 92656 118238 92712
rect 118294 92656 120060 92712
rect 118233 92654 120060 92656
rect 118233 92651 118299 92654
rect 183369 91626 183435 91629
rect 179860 91624 183435 91626
rect 179860 91568 183374 91624
rect 183430 91568 183435 91624
rect 179860 91566 183435 91568
rect 183369 91563 183435 91566
rect 118141 91218 118207 91221
rect 118141 91216 120060 91218
rect 118141 91160 118146 91216
rect 118202 91160 120060 91216
rect 118141 91158 120060 91160
rect 118141 91155 118207 91158
rect 183461 90266 183527 90269
rect 179860 90264 183527 90266
rect 179860 90208 183466 90264
rect 183522 90208 183527 90264
rect 179860 90206 183527 90208
rect 183461 90203 183527 90206
rect 118325 89722 118391 89725
rect 118325 89720 120060 89722
rect 118325 89664 118330 89720
rect 118386 89664 120060 89720
rect 118325 89662 120060 89664
rect 118325 89659 118391 89662
rect 183369 88906 183435 88909
rect 179860 88904 183435 88906
rect 179860 88848 183374 88904
rect 183430 88848 183435 88904
rect 179860 88846 183435 88848
rect 183369 88843 183435 88846
rect 118417 88226 118483 88229
rect 118417 88224 120060 88226
rect 118417 88168 118422 88224
rect 118478 88168 120060 88224
rect 118417 88166 120060 88168
rect 118417 88163 118483 88166
rect 183461 87546 183527 87549
rect 179860 87544 183527 87546
rect 179860 87488 183466 87544
rect 183522 87488 183527 87544
rect 179860 87486 183527 87488
rect 183461 87483 183527 87486
rect 118417 86730 118483 86733
rect 118417 86728 120060 86730
rect 118417 86672 118422 86728
rect 118478 86672 120060 86728
rect 118417 86670 120060 86672
rect 118417 86667 118483 86670
rect 183369 86186 183435 86189
rect 179860 86184 183435 86186
rect 179860 86128 183374 86184
rect 183430 86128 183435 86184
rect 179860 86126 183435 86128
rect 183369 86123 183435 86126
rect 580901 86186 580967 86189
rect 583520 86186 584960 86276
rect 580901 86184 584960 86186
rect 580901 86128 580906 86184
rect 580962 86128 584960 86184
rect 580901 86126 584960 86128
rect 580901 86123 580967 86126
rect 583520 86036 584960 86126
rect 118601 85234 118667 85237
rect 118601 85232 120060 85234
rect 118601 85176 118606 85232
rect 118662 85176 120060 85232
rect 118601 85174 120060 85176
rect 118601 85171 118667 85174
rect 183461 84826 183527 84829
rect 179860 84824 183527 84826
rect -960 84690 480 84780
rect 179860 84768 183466 84824
rect 183522 84768 183527 84824
rect 179860 84766 183527 84768
rect 183461 84763 183527 84766
rect 3509 84690 3575 84693
rect -960 84688 3575 84690
rect -960 84632 3514 84688
rect 3570 84632 3575 84688
rect -960 84630 3575 84632
rect -960 84540 480 84630
rect 3509 84627 3575 84630
rect 118509 83738 118575 83741
rect 118509 83736 120060 83738
rect 118509 83680 118514 83736
rect 118570 83680 120060 83736
rect 118509 83678 120060 83680
rect 118509 83675 118575 83678
rect 183461 83466 183527 83469
rect 179860 83464 183527 83466
rect 179860 83408 183466 83464
rect 183522 83408 183527 83464
rect 179860 83406 183527 83408
rect 183461 83403 183527 83406
rect 118325 82242 118391 82245
rect 118325 82240 120060 82242
rect 118325 82184 118330 82240
rect 118386 82184 120060 82240
rect 118325 82182 120060 82184
rect 118325 82179 118391 82182
rect 183001 82106 183067 82109
rect 179860 82104 183067 82106
rect 179860 82048 183006 82104
rect 183062 82048 183067 82104
rect 179860 82046 183067 82048
rect 183001 82043 183067 82046
rect 182817 80746 182883 80749
rect 179860 80744 182883 80746
rect 179860 80688 182822 80744
rect 182878 80688 182883 80744
rect 179860 80686 182883 80688
rect 182817 80683 182883 80686
rect 118417 80610 118483 80613
rect 580165 80610 580231 80613
rect 118417 80608 580231 80610
rect 118417 80552 118422 80608
rect 118478 80552 580170 80608
rect 580226 80552 580231 80608
rect 118417 80550 580231 80552
rect 118417 80547 118483 80550
rect 580165 80547 580231 80550
rect 172278 80412 172284 80476
rect 172348 80474 172354 80476
rect 580717 80474 580783 80477
rect 172348 80472 580783 80474
rect 172348 80416 580722 80472
rect 580778 80416 580783 80472
rect 172348 80414 580783 80416
rect 172348 80412 172354 80414
rect 580717 80411 580783 80414
rect 171542 80276 171548 80340
rect 171612 80338 171618 80340
rect 180057 80338 180123 80341
rect 171612 80336 180123 80338
rect 171612 80280 180062 80336
rect 180118 80280 180123 80336
rect 171612 80278 180123 80280
rect 171612 80276 171618 80278
rect 180057 80275 180123 80278
rect 123477 80202 123543 80205
rect 123477 80200 132418 80202
rect 123477 80144 123482 80200
rect 123538 80144 132418 80200
rect 123477 80142 132418 80144
rect 123477 80139 123543 80142
rect 132358 79967 132418 80142
rect 159398 80140 159404 80204
rect 159468 80202 159474 80204
rect 171910 80202 171916 80204
rect 159468 80142 171916 80202
rect 159468 80140 159474 80142
rect 171910 80140 171916 80142
rect 171980 80140 171986 80204
rect 178033 80202 178099 80205
rect 172056 80200 178099 80202
rect 172056 80144 178038 80200
rect 178094 80144 178099 80200
rect 172056 80142 178099 80144
rect 167134 80006 167562 80066
rect 125547 79962 125613 79967
rect 125547 79906 125552 79962
rect 125608 79906 125613 79962
rect 125547 79901 125613 79906
rect 125731 79962 125797 79967
rect 125731 79906 125736 79962
rect 125792 79906 125797 79962
rect 125915 79962 125981 79967
rect 126927 79964 126993 79967
rect 125915 79932 125920 79962
rect 125976 79932 125981 79962
rect 126884 79962 126993 79964
rect 125731 79901 125797 79906
rect 125550 79661 125610 79901
rect 125734 79661 125794 79901
rect 125910 79868 125916 79932
rect 125980 79930 125986 79932
rect 126743 79930 126809 79933
rect 125980 79870 126038 79930
rect 126102 79928 126809 79930
rect 126102 79872 126748 79928
rect 126804 79872 126809 79928
rect 126102 79870 126809 79872
rect 125980 79868 125986 79870
rect 125869 79794 125935 79797
rect 126102 79794 126162 79870
rect 126743 79867 126809 79870
rect 126884 79906 126932 79962
rect 126988 79906 126993 79962
rect 126884 79901 126993 79906
rect 127387 79962 127453 79967
rect 127387 79906 127392 79962
rect 127448 79930 127453 79962
rect 127755 79962 127821 79967
rect 127566 79930 127572 79932
rect 127448 79906 127572 79930
rect 127387 79901 127572 79906
rect 126884 79797 126944 79901
rect 127390 79870 127572 79901
rect 127566 79868 127572 79870
rect 127636 79868 127642 79932
rect 127755 79906 127760 79962
rect 127816 79906 127821 79962
rect 127755 79901 127821 79906
rect 128031 79964 128097 79967
rect 128031 79962 128140 79964
rect 128031 79906 128036 79962
rect 128092 79906 128140 79962
rect 128307 79962 128373 79967
rect 128307 79932 128312 79962
rect 128368 79932 128373 79962
rect 129963 79962 130029 79967
rect 128031 79901 128140 79906
rect 127758 79797 127818 79901
rect 125869 79792 126162 79794
rect 125869 79736 125874 79792
rect 125930 79736 126162 79792
rect 125869 79734 126162 79736
rect 126881 79792 126947 79797
rect 126881 79736 126886 79792
rect 126942 79736 126947 79792
rect 125869 79731 125935 79734
rect 126881 79731 126947 79736
rect 127111 79794 127177 79797
rect 127382 79794 127388 79796
rect 127111 79792 127388 79794
rect 127111 79736 127116 79792
rect 127172 79736 127388 79792
rect 127111 79734 127388 79736
rect 127111 79731 127177 79734
rect 127382 79732 127388 79734
rect 127452 79732 127458 79796
rect 127709 79792 127818 79797
rect 127709 79736 127714 79792
rect 127770 79736 127818 79792
rect 127709 79734 127818 79736
rect 127709 79731 127775 79734
rect 125550 79656 125659 79661
rect 125550 79600 125598 79656
rect 125654 79600 125659 79656
rect 125550 79598 125659 79600
rect 125734 79656 125843 79661
rect 125734 79600 125782 79656
rect 125838 79600 125843 79656
rect 125734 79598 125843 79600
rect 128080 79658 128140 79901
rect 128302 79868 128308 79932
rect 128372 79930 128378 79932
rect 128675 79930 128741 79933
rect 129043 79932 129109 79933
rect 128854 79930 128860 79932
rect 128372 79870 128430 79930
rect 128675 79928 128860 79930
rect 128675 79872 128680 79928
rect 128736 79872 128860 79928
rect 128675 79870 128860 79872
rect 128372 79868 128378 79870
rect 128675 79867 128741 79870
rect 128854 79868 128860 79870
rect 128924 79868 128930 79932
rect 129038 79868 129044 79932
rect 129108 79930 129114 79932
rect 129503 79930 129569 79933
rect 129108 79870 129200 79930
rect 129276 79928 129569 79930
rect 129276 79872 129508 79928
rect 129564 79872 129569 79928
rect 129276 79870 129569 79872
rect 129108 79868 129114 79870
rect 129043 79867 129109 79868
rect 129089 79794 129155 79797
rect 129276 79794 129336 79870
rect 129503 79867 129569 79870
rect 129774 79868 129780 79932
rect 129844 79930 129850 79932
rect 129963 79930 129968 79962
rect 129844 79906 129968 79930
rect 130024 79906 130029 79962
rect 130699 79962 130765 79967
rect 130699 79932 130704 79962
rect 130760 79932 130765 79962
rect 130975 79962 131041 79967
rect 129844 79901 130029 79906
rect 129844 79870 130026 79901
rect 129844 79868 129850 79870
rect 130694 79868 130700 79932
rect 130764 79930 130770 79932
rect 130764 79870 130822 79930
rect 130975 79906 130980 79962
rect 131036 79906 131041 79962
rect 131435 79962 131501 79967
rect 131251 79932 131317 79933
rect 131246 79930 131252 79932
rect 130975 79901 131041 79906
rect 130764 79868 130770 79870
rect 129687 79794 129753 79797
rect 129089 79792 129336 79794
rect 129089 79736 129094 79792
rect 129150 79736 129336 79792
rect 129089 79734 129336 79736
rect 129552 79792 129753 79794
rect 129552 79736 129692 79792
rect 129748 79736 129753 79792
rect 129552 79734 129753 79736
rect 129089 79731 129155 79734
rect 128261 79658 128327 79661
rect 128080 79656 128327 79658
rect 128080 79600 128266 79656
rect 128322 79600 128327 79656
rect 128080 79598 128327 79600
rect 129552 79658 129612 79734
rect 129687 79731 129753 79734
rect 129733 79658 129799 79661
rect 129552 79656 129799 79658
rect 129552 79600 129738 79656
rect 129794 79600 129799 79656
rect 129552 79598 129799 79600
rect 125593 79595 125659 79598
rect 125777 79595 125843 79598
rect 128261 79595 128327 79598
rect 129733 79595 129799 79598
rect 130101 79660 130167 79661
rect 130101 79656 130148 79660
rect 130212 79658 130218 79660
rect 130101 79600 130106 79656
rect 130101 79596 130148 79600
rect 130212 79598 130258 79658
rect 130212 79596 130218 79598
rect 130510 79596 130516 79660
rect 130580 79658 130586 79660
rect 130653 79658 130719 79661
rect 130580 79656 130719 79658
rect 130580 79600 130658 79656
rect 130714 79600 130719 79656
rect 130580 79598 130719 79600
rect 130978 79658 131038 79901
rect 131160 79870 131252 79930
rect 131246 79868 131252 79870
rect 131316 79868 131322 79932
rect 131435 79906 131440 79962
rect 131496 79930 131501 79962
rect 132355 79962 132421 79967
rect 131803 79932 131869 79933
rect 131614 79930 131620 79932
rect 131496 79906 131620 79930
rect 131435 79901 131620 79906
rect 131438 79870 131620 79901
rect 131614 79868 131620 79870
rect 131684 79868 131690 79932
rect 131798 79868 131804 79932
rect 131868 79930 131874 79932
rect 131868 79870 131960 79930
rect 132355 79906 132360 79962
rect 132416 79906 132421 79962
rect 133643 79962 133709 79967
rect 132355 79901 132421 79906
rect 132723 79930 132789 79933
rect 133086 79930 133092 79932
rect 132723 79928 133092 79930
rect 132723 79872 132728 79928
rect 132784 79872 133092 79928
rect 132723 79870 133092 79872
rect 131868 79868 131874 79870
rect 131251 79867 131317 79868
rect 131803 79867 131869 79868
rect 132723 79867 132789 79870
rect 133086 79868 133092 79870
rect 133156 79868 133162 79932
rect 133459 79928 133525 79933
rect 133459 79872 133464 79928
rect 133520 79872 133525 79928
rect 133643 79906 133648 79962
rect 133704 79906 133709 79962
rect 134747 79962 134813 79967
rect 133643 79901 133709 79906
rect 133459 79867 133525 79872
rect 132631 79794 132697 79797
rect 133270 79794 133276 79796
rect 132631 79792 133276 79794
rect 132631 79736 132636 79792
rect 132692 79736 133276 79792
rect 132631 79734 133276 79736
rect 132631 79731 132697 79734
rect 133270 79732 133276 79734
rect 133340 79732 133346 79796
rect 131113 79658 131179 79661
rect 130978 79656 131179 79658
rect 130978 79600 131118 79656
rect 131174 79600 131179 79656
rect 130978 79598 131179 79600
rect 130580 79596 130586 79598
rect 130101 79595 130167 79596
rect 130653 79595 130719 79598
rect 131113 79595 131179 79598
rect 131573 79658 131639 79661
rect 133462 79658 133522 79867
rect 133646 79661 133706 79901
rect 133822 79868 133828 79932
rect 133892 79930 133898 79932
rect 134011 79930 134077 79933
rect 133892 79928 134077 79930
rect 133892 79872 134016 79928
rect 134072 79872 134077 79928
rect 134747 79906 134752 79962
rect 134808 79906 134813 79962
rect 135483 79962 135549 79967
rect 135483 79932 135488 79962
rect 135544 79932 135549 79962
rect 135667 79962 135733 79967
rect 134747 79901 134813 79906
rect 133892 79870 134077 79872
rect 133892 79868 133898 79870
rect 134011 79867 134077 79870
rect 134750 79797 134810 79901
rect 135118 79870 135362 79930
rect 134750 79792 134859 79797
rect 134750 79736 134798 79792
rect 134854 79736 134859 79792
rect 134750 79734 134859 79736
rect 134793 79731 134859 79734
rect 131573 79656 133522 79658
rect 131573 79600 131578 79656
rect 131634 79600 133522 79656
rect 131573 79598 133522 79600
rect 133597 79656 133706 79661
rect 133597 79600 133602 79656
rect 133658 79600 133706 79656
rect 133597 79598 133706 79600
rect 134977 79658 135043 79661
rect 135118 79658 135178 79870
rect 135302 79794 135362 79870
rect 135478 79868 135484 79932
rect 135548 79930 135554 79932
rect 135548 79870 135606 79930
rect 135667 79906 135672 79962
rect 135728 79930 135733 79962
rect 138979 79962 139045 79967
rect 135846 79930 135852 79932
rect 135728 79906 135852 79930
rect 135667 79901 135852 79906
rect 135670 79870 135852 79901
rect 135548 79868 135554 79870
rect 135846 79868 135852 79870
rect 135916 79868 135922 79932
rect 136403 79928 136469 79933
rect 136403 79872 136408 79928
rect 136464 79872 136469 79928
rect 136403 79867 136469 79872
rect 136771 79928 136837 79933
rect 136771 79872 136776 79928
rect 136832 79872 136837 79928
rect 136771 79867 136837 79872
rect 137686 79868 137692 79932
rect 137756 79930 137762 79932
rect 137967 79930 138033 79933
rect 137756 79928 138033 79930
rect 137756 79872 137972 79928
rect 138028 79872 138033 79928
rect 137756 79870 138033 79872
rect 137756 79868 137762 79870
rect 137967 79867 138033 79870
rect 138422 79868 138428 79932
rect 138492 79930 138498 79932
rect 138611 79930 138677 79933
rect 138492 79928 138677 79930
rect 138492 79872 138616 79928
rect 138672 79872 138677 79928
rect 138979 79906 138984 79962
rect 139040 79906 139045 79962
rect 142383 79964 142449 79967
rect 143487 79964 143553 79967
rect 144039 79964 144105 79967
rect 142383 79962 142722 79964
rect 138979 79901 139045 79906
rect 139623 79930 139689 79933
rect 139623 79928 139962 79930
rect 138492 79870 138677 79872
rect 138492 79868 138498 79870
rect 138611 79867 138677 79870
rect 135621 79794 135687 79797
rect 135302 79792 135687 79794
rect 135302 79736 135626 79792
rect 135682 79736 135687 79792
rect 135302 79734 135687 79736
rect 135621 79731 135687 79734
rect 134977 79656 135178 79658
rect 134977 79600 134982 79656
rect 135038 79600 135178 79656
rect 134977 79598 135178 79600
rect 135713 79658 135779 79661
rect 136406 79658 136466 79867
rect 136774 79797 136834 79867
rect 136725 79792 136834 79797
rect 136955 79794 137021 79797
rect 137875 79796 137941 79797
rect 137870 79794 137876 79796
rect 136725 79736 136730 79792
rect 136786 79736 136834 79792
rect 136725 79734 136834 79736
rect 136912 79792 137021 79794
rect 136912 79736 136960 79792
rect 137016 79736 137021 79792
rect 136725 79731 136791 79734
rect 136912 79731 137021 79736
rect 137784 79734 137876 79794
rect 137870 79732 137876 79734
rect 137940 79732 137946 79796
rect 138606 79732 138612 79796
rect 138676 79794 138682 79796
rect 138982 79794 139042 79901
rect 139623 79872 139628 79928
rect 139684 79872 139962 79928
rect 139623 79870 139962 79872
rect 139623 79867 139689 79870
rect 138676 79734 139042 79794
rect 138676 79732 138682 79734
rect 137875 79731 137941 79732
rect 136912 79661 136972 79731
rect 139902 79661 139962 79870
rect 140262 79868 140268 79932
rect 140332 79930 140338 79932
rect 140543 79930 140609 79933
rect 140332 79928 140609 79930
rect 140332 79872 140548 79928
rect 140604 79872 140609 79928
rect 140332 79870 140609 79872
rect 140332 79868 140338 79870
rect 140543 79867 140609 79870
rect 140998 79868 141004 79932
rect 141068 79930 141074 79932
rect 142107 79930 142173 79933
rect 141068 79928 142173 79930
rect 141068 79872 142112 79928
rect 142168 79872 142173 79928
rect 142383 79906 142388 79962
rect 142444 79932 142722 79962
rect 143487 79962 143826 79964
rect 142444 79906 142660 79932
rect 142383 79904 142660 79906
rect 142383 79901 142449 79904
rect 141068 79870 142173 79872
rect 141068 79868 141074 79870
rect 142107 79867 142173 79870
rect 142654 79868 142660 79904
rect 142724 79868 142730 79932
rect 143119 79930 143185 79933
rect 142846 79928 143185 79930
rect 142846 79872 143124 79928
rect 143180 79872 143185 79928
rect 143487 79906 143492 79962
rect 143548 79932 143826 79962
rect 144039 79962 144378 79964
rect 143548 79906 143764 79932
rect 143487 79904 143764 79906
rect 143487 79901 143553 79904
rect 142846 79870 143185 79872
rect 142846 79797 142906 79870
rect 143119 79867 143185 79870
rect 143758 79868 143764 79904
rect 143828 79868 143834 79932
rect 144039 79906 144044 79962
rect 144100 79932 144378 79962
rect 144499 79962 144565 79967
rect 144100 79906 144316 79932
rect 144039 79904 144316 79906
rect 144039 79901 144105 79904
rect 144310 79868 144316 79904
rect 144380 79868 144386 79932
rect 144499 79906 144504 79962
rect 144560 79906 144565 79962
rect 152043 79962 152109 79967
rect 144499 79901 144565 79906
rect 140451 79796 140517 79797
rect 140446 79794 140452 79796
rect 140360 79734 140452 79794
rect 140446 79732 140452 79734
rect 140516 79732 140522 79796
rect 140819 79792 140885 79797
rect 140819 79736 140824 79792
rect 140880 79736 140885 79792
rect 140451 79731 140517 79732
rect 140819 79731 140885 79736
rect 142846 79792 142955 79797
rect 142846 79736 142894 79792
rect 142950 79736 142955 79792
rect 142846 79734 142955 79736
rect 142889 79731 142955 79734
rect 135713 79656 136466 79658
rect 135713 79600 135718 79656
rect 135774 79600 136466 79656
rect 135713 79598 136466 79600
rect 136909 79656 136975 79661
rect 136909 79600 136914 79656
rect 136970 79600 136975 79656
rect 131573 79595 131639 79598
rect 133597 79595 133663 79598
rect 134977 79595 135043 79598
rect 135713 79595 135779 79598
rect 136909 79595 136975 79600
rect 139902 79656 140011 79661
rect 139902 79600 139950 79656
rect 140006 79600 140011 79656
rect 139902 79598 140011 79600
rect 140822 79658 140882 79731
rect 144502 79661 144562 79901
rect 145598 79868 145604 79932
rect 145668 79930 145674 79932
rect 146155 79930 146221 79933
rect 146615 79930 146681 79933
rect 146891 79932 146957 79933
rect 147259 79932 147325 79933
rect 146886 79930 146892 79932
rect 145668 79928 146221 79930
rect 145668 79872 146160 79928
rect 146216 79872 146221 79928
rect 145668 79870 146221 79872
rect 145668 79868 145674 79870
rect 146155 79867 146221 79870
rect 146342 79928 146681 79930
rect 146342 79872 146620 79928
rect 146676 79872 146681 79928
rect 146342 79870 146681 79872
rect 146800 79870 146892 79930
rect 144775 79794 144841 79797
rect 144775 79792 145114 79794
rect 144775 79736 144780 79792
rect 144836 79736 145114 79792
rect 144775 79734 145114 79736
rect 144775 79731 144841 79734
rect 141233 79658 141299 79661
rect 140822 79656 141299 79658
rect 140822 79600 141238 79656
rect 141294 79600 141299 79656
rect 140822 79598 141299 79600
rect 139945 79595 140011 79598
rect 141233 79595 141299 79598
rect 144453 79656 144562 79661
rect 144453 79600 144458 79656
rect 144514 79600 144562 79656
rect 144453 79598 144562 79600
rect 145054 79658 145114 79734
rect 145230 79732 145236 79796
rect 145300 79794 145306 79796
rect 146063 79794 146129 79797
rect 145300 79792 146129 79794
rect 145300 79736 146068 79792
rect 146124 79736 146129 79792
rect 145300 79734 146129 79736
rect 146342 79794 146402 79870
rect 146615 79867 146681 79870
rect 146886 79868 146892 79870
rect 146956 79868 146962 79932
rect 147254 79930 147260 79932
rect 147168 79870 147260 79930
rect 147254 79868 147260 79870
rect 147324 79868 147330 79932
rect 148087 79930 148153 79933
rect 147814 79928 148153 79930
rect 147814 79872 148092 79928
rect 148148 79872 148153 79928
rect 147814 79870 148153 79872
rect 146891 79867 146957 79868
rect 147259 79867 147325 79868
rect 146707 79796 146773 79797
rect 146518 79794 146524 79796
rect 146342 79734 146524 79794
rect 145300 79732 145306 79734
rect 146063 79731 146129 79734
rect 146518 79732 146524 79734
rect 146588 79732 146594 79796
rect 146702 79732 146708 79796
rect 146772 79794 146778 79796
rect 146772 79734 146864 79794
rect 146772 79732 146778 79734
rect 146707 79731 146773 79732
rect 147029 79658 147095 79661
rect 145054 79656 147095 79658
rect 145054 79600 147034 79656
rect 147090 79600 147095 79656
rect 145054 79598 147095 79600
rect 147814 79658 147874 79870
rect 148087 79867 148153 79870
rect 148358 79868 148364 79932
rect 148428 79930 148434 79932
rect 148547 79930 148613 79933
rect 148428 79928 148613 79930
rect 148428 79872 148552 79928
rect 148608 79872 148613 79928
rect 148428 79870 148613 79872
rect 148428 79868 148434 79870
rect 148547 79867 148613 79870
rect 148726 79868 148732 79932
rect 148796 79930 148802 79932
rect 148915 79930 148981 79933
rect 148796 79928 148981 79930
rect 148796 79872 148920 79928
rect 148976 79872 148981 79928
rect 148796 79870 148981 79872
rect 148796 79868 148802 79870
rect 148915 79867 148981 79870
rect 149651 79928 149717 79933
rect 149651 79872 149656 79928
rect 149712 79872 149717 79928
rect 149651 79867 149717 79872
rect 149830 79868 149836 79932
rect 149900 79930 149906 79932
rect 150111 79930 150177 79933
rect 151675 79932 151741 79933
rect 151670 79930 151676 79932
rect 149900 79928 150177 79930
rect 149900 79872 150116 79928
rect 150172 79872 150177 79928
rect 149900 79870 150177 79872
rect 149900 79868 149906 79870
rect 150111 79867 150177 79870
rect 150571 79894 150637 79899
rect 149654 79797 149714 79867
rect 150571 79838 150576 79894
rect 150632 79838 150637 79894
rect 151584 79870 151676 79930
rect 151670 79868 151676 79870
rect 151740 79868 151746 79932
rect 152043 79906 152048 79962
rect 152104 79906 152109 79962
rect 152411 79962 152477 79967
rect 153055 79964 153121 79967
rect 152411 79930 152416 79962
rect 152043 79901 152109 79906
rect 152276 79906 152416 79930
rect 152472 79906 152477 79962
rect 153012 79962 153121 79964
rect 153012 79932 153060 79962
rect 152276 79901 152477 79906
rect 151675 79867 151741 79868
rect 150571 79833 150637 79838
rect 148542 79732 148548 79796
rect 148612 79794 148618 79796
rect 149007 79794 149073 79797
rect 148612 79792 149073 79794
rect 148612 79736 149012 79792
rect 149068 79736 149073 79792
rect 148612 79734 149073 79736
rect 148612 79732 148618 79734
rect 149007 79731 149073 79734
rect 149605 79792 149714 79797
rect 149605 79736 149610 79792
rect 149666 79736 149714 79792
rect 149605 79734 149714 79736
rect 149605 79731 149671 79734
rect 150014 79732 150020 79796
rect 150084 79794 150090 79796
rect 150295 79794 150361 79797
rect 150084 79792 150361 79794
rect 150084 79736 150300 79792
rect 150356 79736 150361 79792
rect 150084 79734 150361 79736
rect 150084 79732 150090 79734
rect 150295 79731 150361 79734
rect 150574 79661 150634 79833
rect 152046 79797 152106 79901
rect 151997 79792 152106 79797
rect 151997 79736 152002 79792
rect 152058 79736 152106 79792
rect 151997 79734 152106 79736
rect 152276 79870 152474 79901
rect 151997 79731 152063 79734
rect 147949 79658 148015 79661
rect 147814 79656 148015 79658
rect 147814 79600 147954 79656
rect 148010 79600 148015 79656
rect 147814 79598 148015 79600
rect 144453 79595 144519 79598
rect 147029 79595 147095 79598
rect 147949 79595 148015 79598
rect 150525 79656 150634 79661
rect 151905 79660 151971 79661
rect 151854 79658 151860 79660
rect 150525 79600 150530 79656
rect 150586 79600 150634 79656
rect 150525 79598 150634 79600
rect 151814 79598 151860 79658
rect 151924 79656 151971 79660
rect 151966 79600 151971 79656
rect 150525 79595 150591 79598
rect 151854 79596 151860 79598
rect 151924 79596 151971 79600
rect 152276 79658 152336 79870
rect 152958 79868 152964 79932
rect 153028 79906 153060 79932
rect 153116 79906 153121 79962
rect 153028 79901 153121 79906
rect 153239 79962 153305 79967
rect 153239 79906 153244 79962
rect 153300 79906 153305 79962
rect 153239 79901 153305 79906
rect 153423 79962 153489 79967
rect 158391 79964 158457 79967
rect 153423 79906 153428 79962
rect 153484 79930 153489 79962
rect 158118 79962 158457 79964
rect 153694 79930 153700 79932
rect 153484 79906 153700 79930
rect 153423 79901 153700 79906
rect 153028 79870 153072 79901
rect 153028 79868 153034 79870
rect 152406 79732 152412 79796
rect 152476 79794 152482 79796
rect 152871 79794 152937 79797
rect 152476 79792 152937 79794
rect 152476 79736 152876 79792
rect 152932 79736 152937 79792
rect 152476 79734 152937 79736
rect 152476 79732 152482 79734
rect 152871 79731 152937 79734
rect 152457 79658 152523 79661
rect 152276 79656 152523 79658
rect 152276 79600 152462 79656
rect 152518 79600 152523 79656
rect 152276 79598 152523 79600
rect 153242 79658 153302 79901
rect 153426 79870 153700 79901
rect 153694 79868 153700 79870
rect 153764 79868 153770 79932
rect 153878 79868 153884 79932
rect 153948 79930 153954 79932
rect 154343 79930 154409 79933
rect 153948 79928 154409 79930
rect 153948 79872 154348 79928
rect 154404 79872 154409 79928
rect 153948 79870 154409 79872
rect 153948 79868 153954 79870
rect 154343 79867 154409 79870
rect 156822 79868 156828 79932
rect 156892 79930 156898 79932
rect 157103 79930 157169 79933
rect 158118 79932 158396 79962
rect 156892 79928 157169 79930
rect 156892 79872 157108 79928
rect 157164 79872 157169 79928
rect 156892 79870 157169 79872
rect 156892 79868 156898 79870
rect 157103 79867 157169 79870
rect 158110 79868 158116 79932
rect 158180 79906 158396 79932
rect 158452 79906 158457 79962
rect 158180 79904 158457 79906
rect 158180 79868 158186 79904
rect 158391 79901 158457 79904
rect 159403 79962 159469 79967
rect 159863 79964 159929 79967
rect 159403 79906 159408 79962
rect 159464 79906 159469 79962
rect 159403 79901 159469 79906
rect 159820 79962 159929 79964
rect 159820 79906 159868 79962
rect 159924 79930 159929 79962
rect 160134 79930 160140 79932
rect 159924 79906 160140 79930
rect 154062 79732 154068 79796
rect 154132 79794 154138 79796
rect 154527 79794 154593 79797
rect 154132 79792 154593 79794
rect 154132 79736 154532 79792
rect 154588 79736 154593 79792
rect 154132 79734 154593 79736
rect 154132 79732 154138 79734
rect 154527 79731 154593 79734
rect 154982 79732 154988 79796
rect 155052 79794 155058 79796
rect 155263 79794 155329 79797
rect 155052 79792 155329 79794
rect 155052 79736 155268 79792
rect 155324 79736 155329 79792
rect 155052 79734 155329 79736
rect 155052 79732 155058 79734
rect 155263 79731 155329 79734
rect 155902 79732 155908 79796
rect 155972 79794 155978 79796
rect 156413 79794 156479 79797
rect 155972 79792 156479 79794
rect 155972 79736 156418 79792
rect 156474 79736 156479 79792
rect 155972 79734 156479 79736
rect 155972 79732 155978 79734
rect 156413 79731 156479 79734
rect 156638 79732 156644 79796
rect 156708 79794 156714 79796
rect 157195 79794 157261 79797
rect 156708 79792 157261 79794
rect 156708 79736 157200 79792
rect 157256 79736 157261 79792
rect 156708 79734 157261 79736
rect 156708 79732 156714 79734
rect 157195 79731 157261 79734
rect 158299 79794 158365 79797
rect 158478 79794 158484 79796
rect 158299 79792 158484 79794
rect 158299 79736 158304 79792
rect 158360 79736 158484 79792
rect 158299 79734 158484 79736
rect 158299 79731 158365 79734
rect 158478 79732 158484 79734
rect 158548 79732 158554 79796
rect 159081 79794 159147 79797
rect 159265 79794 159331 79797
rect 159081 79792 159331 79794
rect 159081 79736 159086 79792
rect 159142 79736 159270 79792
rect 159326 79736 159331 79792
rect 159081 79734 159331 79736
rect 159406 79794 159466 79901
rect 159820 79870 160140 79906
rect 160134 79868 160140 79870
rect 160204 79868 160210 79932
rect 160507 79928 160573 79933
rect 160507 79872 160512 79928
rect 160568 79872 160573 79928
rect 160507 79867 160573 79872
rect 160686 79868 160692 79932
rect 160756 79930 160762 79932
rect 161243 79930 161309 79933
rect 161979 79932 162045 79933
rect 161974 79930 161980 79932
rect 160756 79928 161309 79930
rect 160756 79872 161248 79928
rect 161304 79872 161309 79928
rect 160756 79870 161309 79872
rect 161888 79870 161980 79930
rect 160756 79868 160762 79870
rect 161243 79867 161309 79870
rect 161974 79868 161980 79870
rect 162044 79868 162050 79932
rect 162158 79868 162164 79932
rect 162228 79930 162234 79932
rect 162623 79930 162689 79933
rect 162228 79928 162689 79930
rect 162228 79872 162628 79928
rect 162684 79872 162689 79928
rect 162228 79870 162689 79872
rect 162228 79868 162234 79870
rect 161979 79867 162045 79868
rect 162623 79867 162689 79870
rect 162991 79930 163057 79933
rect 163262 79930 163268 79932
rect 162991 79928 163268 79930
rect 162991 79872 162996 79928
rect 163052 79872 163268 79928
rect 162991 79870 163268 79872
rect 162991 79867 163057 79870
rect 163262 79868 163268 79870
rect 163332 79868 163338 79932
rect 163446 79868 163452 79932
rect 163516 79930 163522 79932
rect 164003 79930 164069 79933
rect 163516 79928 164069 79930
rect 163516 79872 164008 79928
rect 164064 79872 164069 79928
rect 163516 79870 164069 79872
rect 163516 79868 163522 79870
rect 164003 79867 164069 79870
rect 164187 79930 164253 79933
rect 164734 79930 164740 79932
rect 164187 79928 164740 79930
rect 164187 79872 164192 79928
rect 164248 79872 164740 79928
rect 164187 79870 164740 79872
rect 164187 79867 164253 79870
rect 164734 79868 164740 79870
rect 164804 79868 164810 79932
rect 165291 79930 165357 79933
rect 165470 79930 165476 79932
rect 165291 79928 165476 79930
rect 165291 79872 165296 79928
rect 165352 79872 165476 79928
rect 165291 79870 165476 79872
rect 165291 79867 165357 79870
rect 165470 79868 165476 79870
rect 165540 79868 165546 79932
rect 165751 79930 165817 79933
rect 165751 79928 166090 79930
rect 165751 79872 165756 79928
rect 165812 79872 166090 79928
rect 165751 79870 166090 79872
rect 165751 79867 165817 79870
rect 159766 79794 159772 79796
rect 159406 79734 159772 79794
rect 159081 79731 159147 79734
rect 159265 79731 159331 79734
rect 159766 79732 159772 79734
rect 159836 79732 159842 79796
rect 160369 79794 160435 79797
rect 160510 79794 160570 79867
rect 160369 79792 160570 79794
rect 160369 79736 160374 79792
rect 160430 79736 160570 79792
rect 160369 79734 160570 79736
rect 160737 79794 160803 79797
rect 162899 79796 162965 79797
rect 160870 79794 160876 79796
rect 160737 79792 160876 79794
rect 160737 79736 160742 79792
rect 160798 79736 160876 79792
rect 160737 79734 160876 79736
rect 160369 79731 160435 79734
rect 160737 79731 160803 79734
rect 160870 79732 160876 79734
rect 160940 79732 160946 79796
rect 162894 79794 162900 79796
rect 162808 79734 162900 79794
rect 162894 79732 162900 79734
rect 162964 79732 162970 79796
rect 163630 79732 163636 79796
rect 163700 79794 163706 79796
rect 164095 79794 164161 79797
rect 163700 79792 164161 79794
rect 163700 79736 164100 79792
rect 164156 79736 164161 79792
rect 163700 79734 164161 79736
rect 163700 79732 163706 79734
rect 162899 79731 162965 79732
rect 164095 79731 164161 79734
rect 165286 79732 165292 79796
rect 165356 79794 165362 79796
rect 165475 79794 165541 79797
rect 165356 79792 165541 79794
rect 165356 79736 165480 79792
rect 165536 79736 165541 79792
rect 165356 79734 165541 79736
rect 165356 79732 165362 79734
rect 165475 79731 165541 79734
rect 154481 79658 154547 79661
rect 153242 79656 154547 79658
rect 153242 79600 154486 79656
rect 154542 79600 154547 79656
rect 153242 79598 154547 79600
rect 151905 79595 151971 79596
rect 152457 79595 152523 79598
rect 154481 79595 154547 79598
rect 154665 79658 154731 79661
rect 164877 79658 164943 79661
rect 154665 79656 164943 79658
rect 154665 79600 154670 79656
rect 154726 79600 164882 79656
rect 164938 79600 164943 79656
rect 154665 79598 164943 79600
rect 154665 79595 154731 79598
rect 164877 79595 164943 79598
rect 165889 79658 165955 79661
rect 166030 79658 166090 79870
rect 166206 79868 166212 79932
rect 166276 79930 166282 79932
rect 166763 79930 166829 79933
rect 166276 79928 166829 79930
rect 166276 79872 166768 79928
rect 166824 79872 166829 79928
rect 166276 79870 166829 79872
rect 166276 79868 166282 79870
rect 166763 79867 166829 79870
rect 166574 79732 166580 79796
rect 166644 79794 166650 79796
rect 166855 79794 166921 79797
rect 166644 79792 166921 79794
rect 166644 79736 166860 79792
rect 166916 79736 166921 79792
rect 166644 79734 166921 79736
rect 166644 79732 166650 79734
rect 166855 79731 166921 79734
rect 165889 79656 166090 79658
rect 165889 79600 165894 79656
rect 165950 79600 166090 79656
rect 165889 79598 166090 79600
rect 167134 79661 167194 80006
rect 167315 79928 167381 79933
rect 167315 79872 167320 79928
rect 167376 79872 167381 79928
rect 167315 79867 167381 79872
rect 167502 79930 167562 80006
rect 172056 79967 172116 80142
rect 178033 80139 178099 80142
rect 170903 79964 170969 79967
rect 171179 79964 171245 79967
rect 171312 79964 171318 79966
rect 170903 79962 171012 79964
rect 167683 79930 167749 79933
rect 167502 79928 167749 79930
rect 167502 79872 167688 79928
rect 167744 79872 167749 79928
rect 167502 79870 167749 79872
rect 167683 79867 167749 79870
rect 168046 79868 168052 79932
rect 168116 79930 168122 79932
rect 168235 79930 168301 79933
rect 168787 79932 168853 79933
rect 168782 79930 168788 79932
rect 168116 79928 168301 79930
rect 168116 79872 168240 79928
rect 168296 79872 168301 79928
rect 168116 79870 168301 79872
rect 168696 79870 168788 79930
rect 168116 79868 168122 79870
rect 168235 79867 168301 79870
rect 168782 79868 168788 79870
rect 168852 79868 168858 79932
rect 168971 79930 169037 79933
rect 170259 79932 170325 79933
rect 169518 79930 169524 79932
rect 168971 79928 169524 79930
rect 168971 79872 168976 79928
rect 169032 79872 169524 79928
rect 168971 79870 169524 79872
rect 168787 79867 168853 79868
rect 168971 79867 169037 79870
rect 169518 79868 169524 79870
rect 169588 79868 169594 79932
rect 170254 79930 170260 79932
rect 170168 79870 170260 79930
rect 170254 79868 170260 79870
rect 170324 79868 170330 79932
rect 170903 79906 170908 79962
rect 170964 79906 171012 79962
rect 170903 79901 171012 79906
rect 171179 79962 171318 79964
rect 171179 79906 171184 79962
rect 171240 79906 171318 79962
rect 171179 79904 171318 79906
rect 171179 79901 171245 79904
rect 171312 79902 171318 79904
rect 171382 79902 171388 79966
rect 171455 79964 171521 79967
rect 171455 79962 171564 79964
rect 171455 79906 171460 79962
rect 171516 79932 171564 79962
rect 171731 79962 171797 79967
rect 171731 79932 171736 79962
rect 171792 79932 171797 79962
rect 172007 79962 172116 79967
rect 171516 79906 171548 79932
rect 171455 79901 171548 79906
rect 170259 79867 170325 79868
rect 167134 79656 167243 79661
rect 167134 79600 167182 79656
rect 167238 79600 167243 79656
rect 167134 79598 167243 79600
rect 167318 79658 167378 79867
rect 167862 79732 167868 79796
rect 167932 79794 167938 79796
rect 168051 79794 168117 79797
rect 167932 79792 168117 79794
rect 167932 79736 168056 79792
rect 168112 79736 168117 79792
rect 167932 79734 168117 79736
rect 167932 79732 167938 79734
rect 168051 79731 168117 79734
rect 169334 79732 169340 79796
rect 169404 79794 169410 79796
rect 169707 79794 169773 79797
rect 170811 79796 170877 79797
rect 170952 79796 171012 79901
rect 171504 79870 171548 79901
rect 171542 79868 171548 79870
rect 171612 79868 171618 79932
rect 171726 79868 171732 79932
rect 171796 79930 171802 79932
rect 171796 79870 171854 79930
rect 172007 79906 172012 79962
rect 172068 79906 172116 79962
rect 172007 79904 172116 79906
rect 172375 79962 172441 79967
rect 172375 79906 172380 79962
rect 172436 79930 172441 79962
rect 173203 79962 173269 79967
rect 173203 79932 173208 79962
rect 173264 79932 173269 79962
rect 173014 79930 173020 79932
rect 172436 79906 173020 79930
rect 172007 79901 172073 79904
rect 172375 79901 173020 79906
rect 172378 79870 173020 79901
rect 171796 79868 171802 79870
rect 173014 79868 173020 79870
rect 173084 79868 173090 79932
rect 173198 79868 173204 79932
rect 173268 79930 173274 79932
rect 173268 79870 173326 79930
rect 173571 79928 173637 79933
rect 174031 79930 174097 79933
rect 173571 79872 173576 79928
rect 173632 79872 173637 79928
rect 173268 79868 173274 79870
rect 173571 79867 173637 79872
rect 173758 79928 174097 79930
rect 173758 79872 174036 79928
rect 174092 79872 174097 79928
rect 173758 79870 174097 79872
rect 170806 79794 170812 79796
rect 169404 79792 169773 79794
rect 169404 79736 169712 79792
rect 169768 79736 169773 79792
rect 169404 79734 169773 79736
rect 170720 79734 170812 79794
rect 169404 79732 169410 79734
rect 169707 79731 169773 79734
rect 170806 79732 170812 79734
rect 170876 79732 170882 79796
rect 170952 79734 170996 79796
rect 170990 79732 170996 79734
rect 171060 79732 171066 79796
rect 171174 79732 171180 79796
rect 171244 79794 171250 79796
rect 173574 79794 173634 79867
rect 171244 79734 173634 79794
rect 171244 79732 171250 79734
rect 170811 79731 170877 79732
rect 168097 79658 168163 79661
rect 167318 79656 168163 79658
rect 167318 79600 168102 79656
rect 168158 79600 168163 79656
rect 167318 79598 168163 79600
rect 165889 79595 165955 79598
rect 167177 79595 167243 79598
rect 168097 79595 168163 79598
rect 168741 79658 168807 79661
rect 171910 79658 171916 79660
rect 168741 79656 171916 79658
rect 168741 79600 168746 79656
rect 168802 79600 171916 79656
rect 168741 79598 171916 79600
rect 168741 79595 168807 79598
rect 171910 79596 171916 79598
rect 171980 79596 171986 79660
rect 172094 79596 172100 79660
rect 172164 79658 172170 79660
rect 173341 79658 173407 79661
rect 172164 79656 173407 79658
rect 172164 79600 173346 79656
rect 173402 79600 173407 79656
rect 172164 79598 173407 79600
rect 173758 79658 173818 79870
rect 174031 79867 174097 79870
rect 173893 79658 173959 79661
rect 173758 79656 173959 79658
rect 173758 79600 173898 79656
rect 173954 79600 173959 79656
rect 173758 79598 173959 79600
rect 172164 79596 172170 79598
rect 173341 79595 173407 79598
rect 173893 79595 173959 79598
rect 119337 79522 119403 79525
rect 165153 79522 165219 79525
rect 173249 79522 173315 79525
rect 119337 79520 164986 79522
rect 119337 79464 119342 79520
rect 119398 79464 164986 79520
rect 119337 79462 164986 79464
rect 119337 79459 119403 79462
rect 115197 79386 115263 79389
rect 164926 79386 164986 79462
rect 165153 79520 173315 79522
rect 165153 79464 165158 79520
rect 165214 79464 173254 79520
rect 173310 79464 173315 79520
rect 165153 79462 173315 79464
rect 165153 79459 165219 79462
rect 173249 79459 173315 79462
rect 173617 79522 173683 79525
rect 177389 79522 177455 79525
rect 173617 79520 177455 79522
rect 173617 79464 173622 79520
rect 173678 79464 177394 79520
rect 177450 79464 177455 79520
rect 173617 79462 177455 79464
rect 173617 79459 173683 79462
rect 177389 79459 177455 79462
rect 172973 79386 173039 79389
rect 115197 79384 160110 79386
rect 115197 79328 115202 79384
rect 115258 79328 160110 79384
rect 115197 79326 160110 79328
rect 164926 79384 173039 79386
rect 164926 79328 172978 79384
rect 173034 79328 173039 79384
rect 164926 79326 173039 79328
rect 115197 79323 115263 79326
rect 4889 79250 4955 79253
rect 159398 79250 159404 79252
rect 4889 79248 159404 79250
rect 4889 79192 4894 79248
rect 4950 79192 159404 79248
rect 4889 79190 159404 79192
rect 4889 79187 4955 79190
rect 159398 79188 159404 79190
rect 159468 79188 159474 79252
rect 160050 79250 160110 79326
rect 172973 79323 173039 79326
rect 173341 79386 173407 79389
rect 174537 79386 174603 79389
rect 173341 79384 174603 79386
rect 173341 79328 173346 79384
rect 173402 79328 174542 79384
rect 174598 79328 174603 79384
rect 173341 79326 174603 79328
rect 173341 79323 173407 79326
rect 174537 79323 174603 79326
rect 173065 79250 173131 79253
rect 160050 79248 173131 79250
rect 160050 79192 173070 79248
rect 173126 79192 173131 79248
rect 160050 79190 173131 79192
rect 173065 79187 173131 79190
rect 3601 79114 3667 79117
rect 173198 79114 173204 79116
rect 3601 79112 173204 79114
rect 3601 79056 3606 79112
rect 3662 79056 173204 79112
rect 3601 79054 173204 79056
rect 3601 79051 3667 79054
rect 173198 79052 173204 79054
rect 173268 79052 173274 79116
rect 3417 78978 3483 78981
rect 170673 78978 170739 78981
rect 3417 78976 170739 78978
rect 3417 78920 3422 78976
rect 3478 78920 170678 78976
rect 170734 78920 170739 78976
rect 3417 78918 170739 78920
rect 3417 78915 3483 78918
rect 170673 78915 170739 78918
rect 170949 78978 171015 78981
rect 171174 78978 171180 78980
rect 170949 78976 171180 78978
rect 170949 78920 170954 78976
rect 171010 78920 171180 78976
rect 170949 78918 171180 78920
rect 170949 78915 171015 78918
rect 171174 78916 171180 78918
rect 171244 78916 171250 78980
rect 171409 78978 171475 78981
rect 172278 78978 172284 78980
rect 171409 78976 172284 78978
rect 171409 78920 171414 78976
rect 171470 78920 172284 78976
rect 171409 78918 172284 78920
rect 171409 78915 171475 78918
rect 172278 78916 172284 78918
rect 172348 78916 172354 78980
rect 172421 78978 172487 78981
rect 178585 78978 178651 78981
rect 172421 78976 178651 78978
rect 172421 78920 172426 78976
rect 172482 78920 178590 78976
rect 178646 78920 178651 78976
rect 172421 78918 178651 78920
rect 172421 78915 172487 78918
rect 178585 78915 178651 78918
rect 179505 78978 179571 78981
rect 266353 78978 266419 78981
rect 179505 78976 266419 78978
rect 179505 78920 179510 78976
rect 179566 78920 266358 78976
rect 266414 78920 266419 78976
rect 179505 78918 266419 78920
rect 179505 78915 179571 78918
rect 266353 78915 266419 78918
rect 125961 78842 126027 78845
rect 126094 78842 126100 78844
rect 125961 78840 126100 78842
rect 125961 78784 125966 78840
rect 126022 78784 126100 78840
rect 125961 78782 126100 78784
rect 125961 78779 126027 78782
rect 126094 78780 126100 78782
rect 126164 78780 126170 78844
rect 129958 78780 129964 78844
rect 130028 78842 130034 78844
rect 130193 78842 130259 78845
rect 130028 78840 130259 78842
rect 130028 78784 130198 78840
rect 130254 78784 130259 78840
rect 130028 78782 130259 78784
rect 130028 78780 130034 78782
rect 130193 78779 130259 78782
rect 130510 78780 130516 78844
rect 130580 78842 130586 78844
rect 130653 78842 130719 78845
rect 130580 78840 130719 78842
rect 130580 78784 130658 78840
rect 130714 78784 130719 78840
rect 130580 78782 130719 78784
rect 130580 78780 130586 78782
rect 130653 78779 130719 78782
rect 151486 78780 151492 78844
rect 151556 78842 151562 78844
rect 151721 78842 151787 78845
rect 151556 78840 151787 78842
rect 151556 78784 151726 78840
rect 151782 78784 151787 78840
rect 151556 78782 151787 78784
rect 151556 78780 151562 78782
rect 151721 78779 151787 78782
rect 157006 78780 157012 78844
rect 157076 78842 157082 78844
rect 157241 78842 157307 78845
rect 157076 78840 157307 78842
rect 157076 78784 157246 78840
rect 157302 78784 157307 78840
rect 157076 78782 157307 78784
rect 157076 78780 157082 78782
rect 157241 78779 157307 78782
rect 163129 78842 163195 78845
rect 171869 78842 171935 78845
rect 163129 78840 171935 78842
rect 163129 78784 163134 78840
rect 163190 78784 171874 78840
rect 171930 78784 171935 78840
rect 163129 78782 171935 78784
rect 163129 78779 163195 78782
rect 171869 78779 171935 78782
rect 172513 78842 172579 78845
rect 397453 78842 397519 78845
rect 172513 78840 397519 78842
rect 172513 78784 172518 78840
rect 172574 78784 397458 78840
rect 397514 78784 397519 78840
rect 172513 78782 397519 78784
rect 172513 78779 172579 78782
rect 397453 78779 397519 78782
rect 125685 78708 125751 78709
rect 127249 78708 127315 78709
rect 125685 78704 125732 78708
rect 125796 78706 125802 78708
rect 127198 78706 127204 78708
rect 125685 78648 125690 78704
rect 125685 78644 125732 78648
rect 125796 78646 125842 78706
rect 127158 78646 127204 78706
rect 127268 78704 127315 78708
rect 127310 78648 127315 78704
rect 125796 78644 125802 78646
rect 127198 78644 127204 78646
rect 127268 78644 127315 78648
rect 125685 78643 125751 78644
rect 127249 78643 127315 78644
rect 129917 78706 129983 78709
rect 135897 78708 135963 78709
rect 130326 78706 130332 78708
rect 129917 78704 130332 78706
rect 129917 78648 129922 78704
rect 129978 78648 130332 78704
rect 129917 78646 130332 78648
rect 129917 78643 129983 78646
rect 130326 78644 130332 78646
rect 130396 78644 130402 78708
rect 135846 78644 135852 78708
rect 135916 78706 135963 78708
rect 135916 78704 136008 78706
rect 135958 78648 136008 78704
rect 135916 78646 136008 78648
rect 135916 78644 135963 78646
rect 151302 78644 151308 78708
rect 151372 78706 151378 78708
rect 151537 78706 151603 78709
rect 155033 78708 155099 78709
rect 151372 78704 151603 78706
rect 151372 78648 151542 78704
rect 151598 78648 151603 78704
rect 151372 78646 151603 78648
rect 151372 78644 151378 78646
rect 135897 78643 135963 78644
rect 151537 78643 151603 78646
rect 154982 78644 154988 78708
rect 155052 78706 155099 78708
rect 155052 78704 155144 78706
rect 155094 78648 155144 78704
rect 155052 78646 155144 78648
rect 155052 78644 155099 78646
rect 159030 78644 159036 78708
rect 159100 78706 159106 78708
rect 159909 78706 159975 78709
rect 159100 78704 159975 78706
rect 159100 78648 159914 78704
rect 159970 78648 159975 78704
rect 159100 78646 159975 78648
rect 159100 78644 159106 78646
rect 155033 78643 155099 78644
rect 159909 78643 159975 78646
rect 162894 78644 162900 78708
rect 162964 78706 162970 78708
rect 165429 78706 165495 78709
rect 162964 78704 165495 78706
rect 162964 78648 165434 78704
rect 165490 78648 165495 78704
rect 162964 78646 165495 78648
rect 162964 78644 162970 78646
rect 165429 78643 165495 78646
rect 168833 78706 168899 78709
rect 170305 78706 170371 78709
rect 168833 78704 170371 78706
rect 168833 78648 168838 78704
rect 168894 78648 170310 78704
rect 170366 78648 170371 78704
rect 168833 78646 170371 78648
rect 168833 78643 168899 78646
rect 170305 78643 170371 78646
rect 170673 78706 170739 78709
rect 171777 78706 171843 78709
rect 170673 78704 171843 78706
rect 170673 78648 170678 78704
rect 170734 78648 171782 78704
rect 171838 78648 171843 78704
rect 170673 78646 171843 78648
rect 170673 78643 170739 78646
rect 171777 78643 171843 78646
rect 173014 78644 173020 78708
rect 173084 78706 173090 78708
rect 462313 78706 462379 78709
rect 173084 78704 462379 78706
rect 173084 78648 462318 78704
rect 462374 78648 462379 78704
rect 173084 78646 462379 78648
rect 173084 78644 173090 78646
rect 462313 78643 462379 78646
rect 125593 78570 125659 78573
rect 125593 78568 157350 78570
rect 125593 78512 125598 78568
rect 125654 78512 157350 78568
rect 125593 78510 157350 78512
rect 125593 78507 125659 78510
rect 157290 78434 157350 78510
rect 159766 78508 159772 78572
rect 159836 78570 159842 78572
rect 159909 78570 159975 78573
rect 159836 78568 159975 78570
rect 159836 78512 159914 78568
rect 159970 78512 159975 78568
rect 159836 78510 159975 78512
rect 159836 78508 159842 78510
rect 159909 78507 159975 78510
rect 160645 78570 160711 78573
rect 167637 78570 167703 78573
rect 160645 78568 167703 78570
rect 160645 78512 160650 78568
rect 160706 78512 167642 78568
rect 167698 78512 167703 78568
rect 160645 78510 167703 78512
rect 160645 78507 160711 78510
rect 167637 78507 167703 78510
rect 168649 78570 168715 78573
rect 172094 78570 172100 78572
rect 168649 78568 172100 78570
rect 168649 78512 168654 78568
rect 168710 78512 172100 78568
rect 168649 78510 172100 78512
rect 168649 78507 168715 78510
rect 172094 78508 172100 78510
rect 172164 78508 172170 78572
rect 164877 78434 164943 78437
rect 168741 78436 168807 78437
rect 171317 78436 171383 78437
rect 168741 78434 168788 78436
rect 157290 78432 164943 78434
rect 157290 78376 164882 78432
rect 164938 78376 164943 78432
rect 157290 78374 164943 78376
rect 168696 78432 168788 78434
rect 168696 78376 168746 78432
rect 168696 78374 168788 78376
rect 164877 78371 164943 78374
rect 168741 78372 168788 78374
rect 168852 78372 168858 78436
rect 171317 78434 171364 78436
rect 171272 78432 171364 78434
rect 171272 78376 171322 78432
rect 171272 78374 171364 78376
rect 171317 78372 171364 78374
rect 171428 78372 171434 78436
rect 171501 78434 171567 78437
rect 174537 78434 174603 78437
rect 171501 78432 174603 78434
rect 171501 78376 171506 78432
rect 171562 78376 174542 78432
rect 174598 78376 174603 78432
rect 171501 78374 174603 78376
rect 168741 78371 168807 78372
rect 171317 78371 171383 78372
rect 171501 78371 171567 78374
rect 174537 78371 174603 78374
rect 122189 78298 122255 78301
rect 127566 78298 127572 78300
rect 122189 78296 127572 78298
rect 122189 78240 122194 78296
rect 122250 78240 127572 78296
rect 122189 78238 127572 78240
rect 122189 78235 122255 78238
rect 127566 78236 127572 78238
rect 127636 78236 127642 78300
rect 158846 78236 158852 78300
rect 158916 78298 158922 78300
rect 160001 78298 160067 78301
rect 158916 78296 160067 78298
rect 158916 78240 160006 78296
rect 160062 78240 160067 78296
rect 158916 78238 160067 78240
rect 158916 78236 158922 78238
rect 160001 78235 160067 78238
rect 163221 78298 163287 78301
rect 171593 78298 171659 78301
rect 163221 78296 171659 78298
rect 163221 78240 163226 78296
rect 163282 78240 171598 78296
rect 171654 78240 171659 78296
rect 163221 78238 171659 78240
rect 163221 78235 163287 78238
rect 171593 78235 171659 78238
rect 172053 78298 172119 78301
rect 182357 78298 182423 78301
rect 172053 78296 182423 78298
rect 172053 78240 172058 78296
rect 172114 78240 182362 78296
rect 182418 78240 182423 78296
rect 172053 78238 182423 78240
rect 172053 78235 172119 78238
rect 182357 78235 182423 78238
rect 127341 78162 127407 78165
rect 128302 78162 128308 78164
rect 127341 78160 128308 78162
rect 127341 78104 127346 78160
rect 127402 78104 128308 78160
rect 127341 78102 128308 78104
rect 127341 78099 127407 78102
rect 128302 78100 128308 78102
rect 128372 78100 128378 78164
rect 128486 78100 128492 78164
rect 128556 78162 128562 78164
rect 128721 78162 128787 78165
rect 128556 78160 128787 78162
rect 128556 78104 128726 78160
rect 128782 78104 128787 78160
rect 128556 78102 128787 78104
rect 128556 78100 128562 78102
rect 128721 78099 128787 78102
rect 153929 78162 153995 78165
rect 154246 78162 154252 78164
rect 153929 78160 154252 78162
rect 153929 78104 153934 78160
rect 153990 78104 154252 78160
rect 153929 78102 154252 78104
rect 153929 78099 153995 78102
rect 154246 78100 154252 78102
rect 154316 78100 154322 78164
rect 159817 78162 159883 78165
rect 171225 78162 171291 78165
rect 159817 78160 171291 78162
rect 159817 78104 159822 78160
rect 159878 78104 171230 78160
rect 171286 78104 171291 78160
rect 159817 78102 171291 78104
rect 159817 78099 159883 78102
rect 171225 78099 171291 78102
rect 171726 78100 171732 78164
rect 171796 78162 171802 78164
rect 179137 78162 179203 78165
rect 171796 78160 179203 78162
rect 171796 78104 179142 78160
rect 179198 78104 179203 78160
rect 171796 78102 179203 78104
rect 171796 78100 171802 78102
rect 179137 78099 179203 78102
rect 153193 78026 153259 78029
rect 157149 78028 157215 78029
rect 153694 78026 153700 78028
rect 153193 78024 153700 78026
rect 153193 77968 153198 78024
rect 153254 77968 153700 78024
rect 153193 77966 153700 77968
rect 153193 77963 153259 77966
rect 153694 77964 153700 77966
rect 153764 77964 153770 78028
rect 157149 78024 157196 78028
rect 157260 78026 157266 78028
rect 157149 77968 157154 78024
rect 157149 77964 157196 77968
rect 157260 77966 157306 78026
rect 157260 77964 157266 77966
rect 157926 77964 157932 78028
rect 157996 78026 158002 78028
rect 158437 78026 158503 78029
rect 157996 78024 158503 78026
rect 157996 77968 158442 78024
rect 158498 77968 158503 78024
rect 157996 77966 158503 77968
rect 157996 77964 158002 77966
rect 157149 77963 157215 77964
rect 158437 77963 158503 77966
rect 158989 78026 159055 78029
rect 164969 78026 165035 78029
rect 255957 78026 256023 78029
rect 158989 78024 165035 78026
rect 158989 77968 158994 78024
rect 159050 77968 164974 78024
rect 165030 77968 165035 78024
rect 158989 77966 165035 77968
rect 158989 77963 159055 77966
rect 164969 77963 165035 77966
rect 169710 78024 256023 78026
rect 169710 77968 255962 78024
rect 256018 77968 256023 78024
rect 169710 77966 256023 77968
rect 10317 77890 10383 77893
rect 126053 77890 126119 77893
rect 10317 77888 126119 77890
rect 10317 77832 10322 77888
rect 10378 77832 126058 77888
rect 126114 77832 126119 77888
rect 10317 77830 126119 77832
rect 10317 77827 10383 77830
rect 126053 77827 126119 77830
rect 133638 77828 133644 77892
rect 133708 77890 133714 77892
rect 147305 77890 147371 77893
rect 133708 77888 147371 77890
rect 133708 77832 147310 77888
rect 147366 77832 147371 77888
rect 133708 77830 147371 77832
rect 133708 77828 133714 77830
rect 147305 77827 147371 77830
rect 154389 77892 154455 77893
rect 154389 77888 154436 77892
rect 154500 77890 154506 77892
rect 154389 77832 154394 77888
rect 154389 77828 154436 77832
rect 154500 77830 154546 77890
rect 154500 77828 154506 77830
rect 158294 77828 158300 77892
rect 158364 77890 158370 77892
rect 158529 77890 158595 77893
rect 158364 77888 158595 77890
rect 158364 77832 158534 77888
rect 158590 77832 158595 77888
rect 158364 77830 158595 77832
rect 158364 77828 158370 77830
rect 154389 77827 154455 77828
rect 158529 77827 158595 77830
rect 162669 77890 162735 77893
rect 169710 77890 169770 77966
rect 255957 77963 256023 77966
rect 170949 77892 171015 77893
rect 170949 77890 170996 77892
rect 162669 77888 169770 77890
rect 162669 77832 162674 77888
rect 162730 77832 169770 77888
rect 162669 77830 169770 77832
rect 170904 77888 170996 77890
rect 170904 77832 170954 77888
rect 170904 77830 170996 77832
rect 162669 77827 162735 77830
rect 170949 77828 170996 77830
rect 171060 77828 171066 77892
rect 171225 77890 171291 77893
rect 171593 77890 171659 77893
rect 483013 77890 483079 77893
rect 171225 77888 171426 77890
rect 171225 77832 171230 77888
rect 171286 77832 171426 77888
rect 171225 77830 171426 77832
rect 170949 77827 171015 77828
rect 171225 77827 171291 77830
rect 171225 77754 171291 77757
rect 160050 77752 171291 77754
rect 160050 77696 171230 77752
rect 171286 77696 171291 77752
rect 160050 77694 171291 77696
rect 171366 77754 171426 77830
rect 171593 77888 483079 77890
rect 171593 77832 171598 77888
rect 171654 77832 483018 77888
rect 483074 77832 483079 77888
rect 171593 77830 483079 77832
rect 171593 77827 171659 77830
rect 483013 77827 483079 77830
rect 172237 77754 172303 77757
rect 171366 77752 172303 77754
rect 171366 77696 172242 77752
rect 172298 77696 172303 77752
rect 171366 77694 172303 77696
rect 151629 77618 151695 77621
rect 154481 77618 154547 77621
rect 151629 77616 154547 77618
rect 151629 77560 151634 77616
rect 151690 77560 154486 77616
rect 154542 77560 154547 77616
rect 151629 77558 154547 77560
rect 151629 77555 151695 77558
rect 154481 77555 154547 77558
rect 151721 77482 151787 77485
rect 151854 77482 151860 77484
rect 151721 77480 151860 77482
rect 151721 77424 151726 77480
rect 151782 77424 151860 77480
rect 151721 77422 151860 77424
rect 151721 77419 151787 77422
rect 151854 77420 151860 77422
rect 151924 77420 151930 77484
rect 158713 77482 158779 77485
rect 160050 77482 160110 77694
rect 171225 77691 171291 77694
rect 172237 77691 172303 77694
rect 164969 77618 165035 77621
rect 172053 77618 172119 77621
rect 164969 77616 172119 77618
rect 164969 77560 164974 77616
rect 165030 77560 172058 77616
rect 172114 77560 172119 77616
rect 164969 77558 172119 77560
rect 164969 77555 165035 77558
rect 172053 77555 172119 77558
rect 158713 77480 160110 77482
rect 158713 77424 158718 77480
rect 158774 77424 160110 77480
rect 158713 77422 160110 77424
rect 170489 77482 170555 77485
rect 170990 77482 170996 77484
rect 170489 77480 170996 77482
rect 170489 77424 170494 77480
rect 170550 77424 170996 77480
rect 170489 77422 170996 77424
rect 158713 77419 158779 77422
rect 170489 77419 170555 77422
rect 170990 77420 170996 77422
rect 171060 77420 171066 77484
rect 128445 77346 128511 77349
rect 128670 77346 128676 77348
rect 128445 77344 128676 77346
rect 128445 77288 128450 77344
rect 128506 77288 128676 77344
rect 128445 77286 128676 77288
rect 128445 77283 128511 77286
rect 128670 77284 128676 77286
rect 128740 77284 128746 77348
rect 152774 77284 152780 77348
rect 152844 77346 152850 77348
rect 153009 77346 153075 77349
rect 155769 77348 155835 77349
rect 152844 77344 153075 77346
rect 152844 77288 153014 77344
rect 153070 77288 153075 77344
rect 152844 77286 153075 77288
rect 152844 77284 152850 77286
rect 153009 77283 153075 77286
rect 155718 77284 155724 77348
rect 155788 77346 155835 77348
rect 159173 77346 159239 77349
rect 160134 77346 160140 77348
rect 155788 77344 155880 77346
rect 155830 77288 155880 77344
rect 155788 77286 155880 77288
rect 159173 77344 160140 77346
rect 159173 77288 159178 77344
rect 159234 77288 160140 77344
rect 159173 77286 160140 77288
rect 155788 77284 155835 77286
rect 155769 77283 155835 77284
rect 159173 77283 159239 77286
rect 160134 77284 160140 77286
rect 160204 77284 160210 77348
rect 169845 77346 169911 77349
rect 172278 77346 172284 77348
rect 169845 77344 172284 77346
rect 169845 77288 169850 77344
rect 169906 77288 172284 77344
rect 169845 77286 172284 77288
rect 169845 77283 169911 77286
rect 172278 77284 172284 77286
rect 172348 77284 172354 77348
rect 142061 77210 142127 77213
rect 164877 77210 164943 77213
rect 142061 77208 164943 77210
rect 142061 77152 142066 77208
rect 142122 77152 164882 77208
rect 164938 77152 164943 77208
rect 142061 77150 164943 77152
rect 142061 77147 142127 77150
rect 164877 77147 164943 77150
rect 169518 77148 169524 77212
rect 169588 77210 169594 77212
rect 172145 77210 172211 77213
rect 169588 77208 172211 77210
rect 169588 77152 172150 77208
rect 172206 77152 172211 77208
rect 169588 77150 172211 77152
rect 169588 77148 169594 77150
rect 172145 77147 172211 77150
rect 147029 77074 147095 77077
rect 247033 77074 247099 77077
rect 147029 77072 247099 77074
rect 147029 77016 147034 77072
rect 147090 77016 247038 77072
rect 247094 77016 247099 77072
rect 147029 77014 247099 77016
rect 147029 77011 147095 77014
rect 247033 77011 247099 77014
rect 136214 76876 136220 76940
rect 136284 76938 136290 76940
rect 136909 76938 136975 76941
rect 136284 76936 136975 76938
rect 136284 76880 136914 76936
rect 136970 76880 136975 76936
rect 136284 76878 136975 76880
rect 136284 76876 136290 76878
rect 136909 76875 136975 76878
rect 147489 76938 147555 76941
rect 282913 76938 282979 76941
rect 147489 76936 282979 76938
rect 147489 76880 147494 76936
rect 147550 76880 282918 76936
rect 282974 76880 282979 76936
rect 147489 76878 282979 76880
rect 147489 76875 147555 76878
rect 282913 76875 282979 76878
rect 111793 76802 111859 76805
rect 134241 76802 134307 76805
rect 111793 76800 134307 76802
rect 111793 76744 111798 76800
rect 111854 76744 134246 76800
rect 134302 76744 134307 76800
rect 111793 76742 134307 76744
rect 111793 76739 111859 76742
rect 134241 76739 134307 76742
rect 136030 76740 136036 76804
rect 136100 76802 136106 76804
rect 139117 76802 139183 76805
rect 136100 76800 139183 76802
rect 136100 76744 139122 76800
rect 139178 76744 139183 76800
rect 136100 76742 139183 76744
rect 136100 76740 136106 76742
rect 139117 76739 139183 76742
rect 144494 76740 144500 76804
rect 144564 76802 144570 76804
rect 144729 76802 144795 76805
rect 144564 76800 144795 76802
rect 144564 76744 144734 76800
rect 144790 76744 144795 76800
rect 144564 76742 144795 76744
rect 144564 76740 144570 76742
rect 144729 76739 144795 76742
rect 146569 76802 146635 76805
rect 146702 76802 146708 76804
rect 146569 76800 146708 76802
rect 146569 76744 146574 76800
rect 146630 76744 146708 76800
rect 146569 76742 146708 76744
rect 146569 76739 146635 76742
rect 146702 76740 146708 76742
rect 146772 76740 146778 76804
rect 156229 76802 156295 76805
rect 354673 76802 354739 76805
rect 156229 76800 354739 76802
rect 156229 76744 156234 76800
rect 156290 76744 354678 76800
rect 354734 76744 354739 76800
rect 156229 76742 354739 76744
rect 156229 76739 156295 76742
rect 354673 76739 354739 76742
rect 37273 76666 37339 76669
rect 128537 76666 128603 76669
rect 37273 76664 128603 76666
rect 37273 76608 37278 76664
rect 37334 76608 128542 76664
rect 128598 76608 128603 76664
rect 37273 76606 128603 76608
rect 37273 76603 37339 76606
rect 128537 76603 128603 76606
rect 131389 76668 131455 76669
rect 131389 76664 131436 76668
rect 131500 76666 131506 76668
rect 131665 76666 131731 76669
rect 134057 76668 134123 76669
rect 131798 76666 131804 76668
rect 131389 76608 131394 76664
rect 131389 76604 131436 76608
rect 131500 76606 131546 76666
rect 131665 76664 131804 76666
rect 131665 76608 131670 76664
rect 131726 76608 131804 76664
rect 131665 76606 131804 76608
rect 131500 76604 131506 76606
rect 131389 76603 131455 76604
rect 131665 76603 131731 76606
rect 131798 76604 131804 76606
rect 131868 76604 131874 76668
rect 134006 76666 134012 76668
rect 133966 76606 134012 76666
rect 134076 76664 134123 76668
rect 134118 76608 134123 76664
rect 134006 76604 134012 76606
rect 134076 76604 134123 76608
rect 135110 76604 135116 76668
rect 135180 76666 135186 76668
rect 137921 76666 137987 76669
rect 135180 76664 137987 76666
rect 135180 76608 137926 76664
rect 137982 76608 137987 76664
rect 135180 76606 137987 76608
rect 135180 76604 135186 76606
rect 134057 76603 134123 76604
rect 137921 76603 137987 76606
rect 138933 76668 138999 76669
rect 138933 76664 138980 76668
rect 139044 76666 139050 76668
rect 138933 76608 138938 76664
rect 138933 76604 138980 76608
rect 139044 76606 139090 76666
rect 139044 76604 139050 76606
rect 140078 76604 140084 76668
rect 140148 76666 140154 76668
rect 140589 76666 140655 76669
rect 140148 76664 140655 76666
rect 140148 76608 140594 76664
rect 140650 76608 140655 76664
rect 140148 76606 140655 76608
rect 140148 76604 140154 76606
rect 138933 76603 138999 76604
rect 140589 76603 140655 76606
rect 143165 76668 143231 76669
rect 143441 76668 143507 76669
rect 143165 76664 143212 76668
rect 143276 76666 143282 76668
rect 143165 76608 143170 76664
rect 143165 76604 143212 76608
rect 143276 76606 143322 76666
rect 143276 76604 143282 76606
rect 143390 76604 143396 76668
rect 143460 76666 143507 76668
rect 143460 76664 143552 76666
rect 143502 76608 143552 76664
rect 143460 76606 143552 76608
rect 143460 76604 143507 76606
rect 144310 76604 144316 76668
rect 144380 76666 144386 76668
rect 144545 76666 144611 76669
rect 144380 76664 144611 76666
rect 144380 76608 144550 76664
rect 144606 76608 144611 76664
rect 144380 76606 144611 76608
rect 144380 76604 144386 76606
rect 143165 76603 143231 76604
rect 143441 76603 143507 76604
rect 144545 76603 144611 76606
rect 145414 76604 145420 76668
rect 145484 76666 145490 76668
rect 146293 76666 146359 76669
rect 145484 76664 146359 76666
rect 145484 76608 146298 76664
rect 146354 76608 146359 76664
rect 145484 76606 146359 76608
rect 145484 76604 145490 76606
rect 146293 76603 146359 76606
rect 146477 76666 146543 76669
rect 148869 76668 148935 76669
rect 146886 76666 146892 76668
rect 146477 76664 146892 76666
rect 146477 76608 146482 76664
rect 146538 76608 146892 76664
rect 146477 76606 146892 76608
rect 146477 76603 146543 76606
rect 146886 76604 146892 76606
rect 146956 76604 146962 76668
rect 148869 76664 148916 76668
rect 148980 76666 148986 76668
rect 148869 76608 148874 76664
rect 148869 76604 148916 76608
rect 148980 76606 149026 76666
rect 148980 76604 148986 76606
rect 155902 76604 155908 76668
rect 155972 76666 155978 76668
rect 389173 76666 389239 76669
rect 155972 76664 389239 76666
rect 155972 76608 389178 76664
rect 389234 76608 389239 76664
rect 155972 76606 389239 76608
rect 155972 76604 155978 76606
rect 148869 76603 148935 76604
rect 389173 76603 389239 76606
rect 20713 76530 20779 76533
rect 123845 76530 123911 76533
rect 20713 76528 123911 76530
rect 20713 76472 20718 76528
rect 20774 76472 123850 76528
rect 123906 76472 123911 76528
rect 20713 76470 123911 76472
rect 20713 76467 20779 76470
rect 123845 76467 123911 76470
rect 130285 76530 130351 76533
rect 130694 76530 130700 76532
rect 130285 76528 130700 76530
rect 130285 76472 130290 76528
rect 130346 76472 130700 76528
rect 130285 76470 130700 76472
rect 130285 76467 130351 76470
rect 130694 76468 130700 76470
rect 130764 76468 130770 76532
rect 136398 76468 136404 76532
rect 136468 76530 136474 76532
rect 137645 76530 137711 76533
rect 136468 76528 137711 76530
rect 136468 76472 137650 76528
rect 137706 76472 137711 76528
rect 136468 76470 137711 76472
rect 136468 76468 136474 76470
rect 137645 76467 137711 76470
rect 138289 76530 138355 76533
rect 138422 76530 138428 76532
rect 138289 76528 138428 76530
rect 138289 76472 138294 76528
rect 138350 76472 138428 76528
rect 138289 76470 138428 76472
rect 138289 76467 138355 76470
rect 138422 76468 138428 76470
rect 138492 76468 138498 76532
rect 143022 76468 143028 76532
rect 143092 76530 143098 76532
rect 143257 76530 143323 76533
rect 143092 76528 143323 76530
rect 143092 76472 143262 76528
rect 143318 76472 143323 76528
rect 143092 76470 143323 76472
rect 143092 76468 143098 76470
rect 143257 76467 143323 76470
rect 144126 76468 144132 76532
rect 144196 76530 144202 76532
rect 144821 76530 144887 76533
rect 144196 76528 144887 76530
rect 144196 76472 144826 76528
rect 144882 76472 144887 76528
rect 144196 76470 144887 76472
rect 144196 76468 144202 76470
rect 144821 76467 144887 76470
rect 146385 76530 146451 76533
rect 146518 76530 146524 76532
rect 146385 76528 146524 76530
rect 146385 76472 146390 76528
rect 146446 76472 146524 76528
rect 146385 76470 146524 76472
rect 146385 76467 146451 76470
rect 146518 76468 146524 76470
rect 146588 76468 146594 76532
rect 160093 76530 160159 76533
rect 161105 76532 161171 76533
rect 160870 76530 160876 76532
rect 160093 76528 160876 76530
rect 160093 76472 160098 76528
rect 160154 76472 160876 76528
rect 160093 76470 160876 76472
rect 160093 76467 160159 76470
rect 160870 76468 160876 76470
rect 160940 76468 160946 76532
rect 161054 76468 161060 76532
rect 161124 76530 161171 76532
rect 161124 76528 161216 76530
rect 161166 76472 161216 76528
rect 161124 76470 161216 76472
rect 161124 76468 161171 76470
rect 161974 76468 161980 76532
rect 162044 76530 162050 76532
rect 162117 76530 162183 76533
rect 162044 76528 162183 76530
rect 162044 76472 162122 76528
rect 162178 76472 162183 76528
rect 162044 76470 162183 76472
rect 162044 76468 162050 76470
rect 161105 76467 161171 76468
rect 162117 76467 162183 76470
rect 162485 76532 162551 76533
rect 162485 76528 162532 76532
rect 162596 76530 162602 76532
rect 162485 76472 162490 76528
rect 162485 76468 162532 76472
rect 162596 76470 162642 76530
rect 162596 76468 162602 76470
rect 163262 76468 163268 76532
rect 163332 76530 163338 76532
rect 163497 76530 163563 76533
rect 163332 76528 163563 76530
rect 163332 76472 163502 76528
rect 163558 76472 163563 76528
rect 163332 76470 163563 76472
rect 163332 76468 163338 76470
rect 162485 76467 162551 76468
rect 163497 76467 163563 76470
rect 164918 76468 164924 76532
rect 164988 76530 164994 76532
rect 165337 76530 165403 76533
rect 164988 76528 165403 76530
rect 164988 76472 165342 76528
rect 165398 76472 165403 76528
rect 164988 76470 165403 76472
rect 164988 76468 164994 76470
rect 165337 76467 165403 76470
rect 166717 76532 166783 76533
rect 166717 76528 166764 76532
rect 166828 76530 166834 76532
rect 166717 76472 166722 76528
rect 166717 76468 166764 76472
rect 166828 76470 166874 76530
rect 166828 76468 166834 76470
rect 167678 76468 167684 76532
rect 167748 76530 167754 76532
rect 168189 76530 168255 76533
rect 167748 76528 168255 76530
rect 167748 76472 168194 76528
rect 168250 76472 168255 76528
rect 167748 76470 168255 76472
rect 167748 76468 167754 76470
rect 166717 76467 166783 76468
rect 168189 76467 168255 76470
rect 169661 76530 169727 76533
rect 565813 76530 565879 76533
rect 169661 76528 565879 76530
rect 169661 76472 169666 76528
rect 169722 76472 565818 76528
rect 565874 76472 565879 76528
rect 169661 76470 565879 76472
rect 169661 76467 169727 76470
rect 565813 76467 565879 76470
rect 142654 76332 142660 76396
rect 142724 76394 142730 76396
rect 146293 76394 146359 76397
rect 142724 76392 146359 76394
rect 142724 76336 146298 76392
rect 146354 76336 146359 76392
rect 142724 76334 146359 76336
rect 142724 76332 142730 76334
rect 146293 76331 146359 76334
rect 162342 76332 162348 76396
rect 162412 76394 162418 76396
rect 162577 76394 162643 76397
rect 162412 76392 162643 76394
rect 162412 76336 162582 76392
rect 162638 76336 162643 76392
rect 162412 76334 162643 76336
rect 162412 76332 162418 76334
rect 162577 76331 162643 76334
rect 165102 76332 165108 76396
rect 165172 76394 165178 76396
rect 165613 76394 165679 76397
rect 165172 76392 165679 76394
rect 165172 76336 165618 76392
rect 165674 76336 165679 76392
rect 165172 76334 165679 76336
rect 165172 76332 165178 76334
rect 165613 76331 165679 76334
rect 166390 76332 166396 76396
rect 166460 76394 166466 76396
rect 166993 76394 167059 76397
rect 166460 76392 167059 76394
rect 166460 76336 166998 76392
rect 167054 76336 167059 76392
rect 166460 76334 167059 76336
rect 166460 76332 166466 76334
rect 166993 76331 167059 76334
rect 167821 76394 167887 76397
rect 173157 76394 173223 76397
rect 167821 76392 173223 76394
rect 167821 76336 167826 76392
rect 167882 76336 173162 76392
rect 173218 76336 173223 76392
rect 167821 76334 173223 76336
rect 167821 76331 167887 76334
rect 173157 76331 173223 76334
rect 164877 76258 164943 76261
rect 175917 76258 175983 76261
rect 164877 76256 175983 76258
rect 164877 76200 164882 76256
rect 164938 76200 175922 76256
rect 175978 76200 175983 76256
rect 164877 76198 175983 76200
rect 164877 76195 164943 76198
rect 175917 76195 175983 76198
rect 170581 76124 170647 76125
rect 170581 76120 170628 76124
rect 170692 76122 170698 76124
rect 170581 76064 170586 76120
rect 170581 76060 170628 76064
rect 170692 76062 170738 76122
rect 170692 76060 170698 76062
rect 170581 76059 170647 76060
rect 128813 75986 128879 75989
rect 129038 75986 129044 75988
rect 128813 75984 129044 75986
rect 128813 75928 128818 75984
rect 128874 75928 129044 75984
rect 128813 75926 129044 75928
rect 128813 75923 128879 75926
rect 129038 75924 129044 75926
rect 129108 75924 129114 75988
rect 169845 75986 169911 75989
rect 170397 75988 170463 75989
rect 170254 75986 170260 75988
rect 169845 75984 170260 75986
rect 169845 75928 169850 75984
rect 169906 75928 170260 75984
rect 169845 75926 170260 75928
rect 169845 75923 169911 75926
rect 170254 75924 170260 75926
rect 170324 75924 170330 75988
rect 170397 75984 170444 75988
rect 170508 75986 170514 75988
rect 170397 75928 170402 75984
rect 170397 75924 170444 75928
rect 170508 75926 170554 75986
rect 170508 75924 170514 75926
rect 170397 75923 170463 75924
rect 120717 75850 120783 75853
rect 125777 75850 125843 75853
rect 120717 75848 125843 75850
rect 120717 75792 120722 75848
rect 120778 75792 125782 75848
rect 125838 75792 125843 75848
rect 120717 75790 125843 75792
rect 120717 75787 120783 75790
rect 125777 75787 125843 75790
rect 139025 75850 139091 75853
rect 171961 75850 172027 75853
rect 139025 75848 172027 75850
rect 139025 75792 139030 75848
rect 139086 75792 171966 75848
rect 172022 75792 172027 75848
rect 139025 75790 172027 75792
rect 139025 75787 139091 75790
rect 171961 75787 172027 75790
rect 139209 75714 139275 75717
rect 176653 75714 176719 75717
rect 139209 75712 176719 75714
rect 139209 75656 139214 75712
rect 139270 75656 176658 75712
rect 176714 75656 176719 75712
rect 139209 75654 176719 75656
rect 139209 75651 139275 75654
rect 176653 75651 176719 75654
rect 157006 75516 157012 75580
rect 157076 75578 157082 75580
rect 402973 75578 403039 75581
rect 157076 75576 403039 75578
rect 157076 75520 402978 75576
rect 403034 75520 403039 75576
rect 157076 75518 403039 75520
rect 157076 75516 157082 75518
rect 402973 75515 403039 75518
rect 161197 75442 161263 75445
rect 459553 75442 459619 75445
rect 161197 75440 459619 75442
rect 161197 75384 161202 75440
rect 161258 75384 459558 75440
rect 459614 75384 459619 75440
rect 161197 75382 459619 75384
rect 161197 75379 161263 75382
rect 459553 75379 459619 75382
rect 164734 75244 164740 75308
rect 164804 75306 164810 75308
rect 496813 75306 496879 75309
rect 164804 75304 496879 75306
rect 164804 75248 496818 75304
rect 496874 75248 496879 75304
rect 164804 75246 496879 75248
rect 164804 75244 164810 75246
rect 496813 75243 496879 75246
rect 75913 75170 75979 75173
rect 131614 75170 131620 75172
rect 75913 75168 131620 75170
rect 75913 75112 75918 75168
rect 75974 75112 131620 75168
rect 75913 75110 131620 75112
rect 75913 75107 75979 75110
rect 131614 75108 131620 75110
rect 131684 75108 131690 75172
rect 149646 75108 149652 75172
rect 149716 75170 149722 75172
rect 150157 75170 150223 75173
rect 149716 75168 150223 75170
rect 149716 75112 150162 75168
rect 150218 75112 150223 75168
rect 149716 75110 150223 75112
rect 149716 75108 149722 75110
rect 150157 75107 150223 75110
rect 169569 75170 169635 75173
rect 549253 75170 549319 75173
rect 169569 75168 549319 75170
rect 169569 75112 169574 75168
rect 169630 75112 549258 75168
rect 549314 75112 549319 75168
rect 169569 75110 549319 75112
rect 169569 75107 169635 75110
rect 549253 75107 549319 75110
rect 147070 74972 147076 75036
rect 147140 75034 147146 75036
rect 147397 75034 147463 75037
rect 147140 75032 147463 75034
rect 147140 74976 147402 75032
rect 147458 74976 147463 75032
rect 147140 74974 147463 74976
rect 147140 74972 147146 74974
rect 147397 74971 147463 74974
rect 164049 75034 164115 75037
rect 172145 75034 172211 75037
rect 164049 75032 172211 75034
rect 164049 74976 164054 75032
rect 164110 74976 172150 75032
rect 172206 74976 172211 75032
rect 164049 74974 172211 74976
rect 164049 74971 164115 74974
rect 172145 74971 172211 74974
rect 122097 74490 122163 74493
rect 125910 74490 125916 74492
rect 122097 74488 125916 74490
rect 122097 74432 122102 74488
rect 122158 74432 125916 74488
rect 122097 74430 125916 74432
rect 122097 74427 122163 74430
rect 125910 74428 125916 74430
rect 125980 74428 125986 74492
rect 147857 74490 147923 74493
rect 148358 74490 148364 74492
rect 147857 74488 148364 74490
rect 147857 74432 147862 74488
rect 147918 74432 148364 74488
rect 147857 74430 148364 74432
rect 147857 74427 147923 74430
rect 148358 74428 148364 74430
rect 148428 74428 148434 74492
rect 140681 74354 140747 74357
rect 174537 74354 174603 74357
rect 140681 74352 174603 74354
rect 140681 74296 140686 74352
rect 140742 74296 174542 74352
rect 174598 74296 174603 74352
rect 140681 74294 174603 74296
rect 140681 74291 140747 74294
rect 174537 74291 174603 74294
rect 143758 74156 143764 74220
rect 143828 74218 143834 74220
rect 230473 74218 230539 74221
rect 143828 74216 230539 74218
rect 143828 74160 230478 74216
rect 230534 74160 230539 74216
rect 143828 74158 230539 74160
rect 143828 74156 143834 74158
rect 230473 74155 230539 74158
rect 148501 74082 148567 74085
rect 244273 74082 244339 74085
rect 148501 74080 244339 74082
rect 148501 74024 148506 74080
rect 148562 74024 244278 74080
rect 244334 74024 244339 74080
rect 148501 74022 244339 74024
rect 148501 74019 148567 74022
rect 244273 74019 244339 74022
rect 71773 73946 71839 73949
rect 131205 73946 131271 73949
rect 71773 73944 131271 73946
rect 71773 73888 71778 73944
rect 71834 73888 131210 73944
rect 131266 73888 131271 73944
rect 71773 73886 131271 73888
rect 71773 73883 71839 73886
rect 131205 73883 131271 73886
rect 148961 73946 149027 73949
rect 284385 73946 284451 73949
rect 148961 73944 284451 73946
rect 148961 73888 148966 73944
rect 149022 73888 284390 73944
rect 284446 73888 284451 73944
rect 148961 73886 284451 73888
rect 148961 73883 149027 73886
rect 284385 73883 284451 73886
rect 35893 73810 35959 73813
rect 128670 73810 128676 73812
rect 35893 73808 128676 73810
rect 35893 73752 35898 73808
rect 35954 73752 128676 73808
rect 35893 73750 128676 73752
rect 35893 73747 35959 73750
rect 128670 73748 128676 73750
rect 128740 73748 128746 73812
rect 150341 73810 150407 73813
rect 318793 73810 318859 73813
rect 150341 73808 318859 73810
rect 150341 73752 150346 73808
rect 150402 73752 318798 73808
rect 318854 73752 318859 73808
rect 150341 73750 318859 73752
rect 150341 73747 150407 73750
rect 318793 73747 318859 73750
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 583520 72844 584960 72934
rect 40033 72586 40099 72589
rect 128854 72586 128860 72588
rect 40033 72584 128860 72586
rect 40033 72528 40038 72584
rect 40094 72528 128860 72584
rect 40033 72526 128860 72528
rect 40033 72523 40099 72526
rect 128854 72524 128860 72526
rect 128924 72524 128930 72588
rect 1393 72450 1459 72453
rect 125726 72450 125732 72452
rect 1393 72448 125732 72450
rect 1393 72392 1398 72448
rect 1454 72392 125732 72448
rect 1393 72390 125732 72392
rect 1393 72387 1459 72390
rect 125726 72388 125732 72390
rect 125796 72388 125802 72452
rect 148685 72450 148751 72453
rect 298093 72450 298159 72453
rect 148685 72448 298159 72450
rect 148685 72392 148690 72448
rect 148746 72392 298098 72448
rect 298154 72392 298159 72448
rect 148685 72390 298159 72392
rect 148685 72387 148751 72390
rect 298093 72387 298159 72390
rect -960 71634 480 71724
rect 3417 71634 3483 71637
rect -960 71632 3483 71634
rect -960 71576 3422 71632
rect 3478 71576 3483 71632
rect -960 71574 3483 71576
rect -960 71484 480 71574
rect 3417 71571 3483 71574
rect 91093 69730 91159 69733
rect 133270 69730 133276 69732
rect 91093 69728 133276 69730
rect 91093 69672 91098 69728
rect 91154 69672 133276 69728
rect 91093 69670 133276 69672
rect 91093 69667 91159 69670
rect 133270 69668 133276 69670
rect 133340 69668 133346 69732
rect 55213 69594 55279 69597
rect 130326 69594 130332 69596
rect 55213 69592 130332 69594
rect 55213 69536 55218 69592
rect 55274 69536 130332 69592
rect 55213 69534 130332 69536
rect 55213 69531 55279 69534
rect 130326 69532 130332 69534
rect 130396 69532 130402 69596
rect 138974 69532 138980 69596
rect 139044 69594 139050 69596
rect 175273 69594 175339 69597
rect 139044 69592 175339 69594
rect 139044 69536 175278 69592
rect 175334 69536 175339 69592
rect 139044 69534 175339 69536
rect 139044 69532 139050 69534
rect 175273 69531 175339 69534
rect 57973 68370 58039 68373
rect 130142 68370 130148 68372
rect 57973 68368 130148 68370
rect 57973 68312 57978 68368
rect 58034 68312 130148 68368
rect 57973 68310 130148 68312
rect 57973 68307 58039 68310
rect 130142 68308 130148 68310
rect 130212 68308 130218 68372
rect 152590 68308 152596 68372
rect 152660 68370 152666 68372
rect 353293 68370 353359 68373
rect 152660 68368 353359 68370
rect 152660 68312 353298 68368
rect 353354 68312 353359 68368
rect 152660 68310 353359 68312
rect 152660 68308 152666 68310
rect 353293 68307 353359 68310
rect 22093 68234 22159 68237
rect 127198 68234 127204 68236
rect 22093 68232 127204 68234
rect 22093 68176 22098 68232
rect 22154 68176 127204 68232
rect 22093 68174 127204 68176
rect 22093 68171 22159 68174
rect 127198 68172 127204 68174
rect 127268 68172 127274 68236
rect 127341 68234 127407 68237
rect 135294 68234 135300 68236
rect 127341 68232 135300 68234
rect 127341 68176 127346 68232
rect 127402 68176 135300 68232
rect 127341 68174 135300 68176
rect 127341 68171 127407 68174
rect 135294 68172 135300 68174
rect 135364 68172 135370 68236
rect 166206 68172 166212 68236
rect 166276 68234 166282 68236
rect 529933 68234 529999 68237
rect 166276 68232 529999 68234
rect 166276 68176 529938 68232
rect 529994 68176 529999 68232
rect 166276 68174 529999 68176
rect 166276 68172 166282 68174
rect 529933 68171 529999 68174
rect 138606 66948 138612 67012
rect 138676 67010 138682 67012
rect 172513 67010 172579 67013
rect 138676 67008 172579 67010
rect 138676 66952 172518 67008
rect 172574 66952 172579 67008
rect 138676 66950 172579 66952
rect 138676 66948 138682 66950
rect 172513 66947 172579 66950
rect 140262 66812 140268 66876
rect 140332 66874 140338 66876
rect 193213 66874 193279 66877
rect 140332 66872 193279 66874
rect 140332 66816 193218 66872
rect 193274 66816 193279 66872
rect 140332 66814 193279 66816
rect 140332 66812 140338 66814
rect 193213 66811 193279 66814
rect 73153 65514 73219 65517
rect 131246 65514 131252 65516
rect 73153 65512 131252 65514
rect 73153 65456 73158 65512
rect 73214 65456 131252 65512
rect 73153 65454 131252 65456
rect 73153 65451 73219 65454
rect 131246 65452 131252 65454
rect 131316 65452 131322 65516
rect 144494 64228 144500 64292
rect 144564 64290 144570 64292
rect 245653 64290 245719 64293
rect 144564 64288 245719 64290
rect 144564 64232 245658 64288
rect 245714 64232 245719 64288
rect 144564 64230 245719 64232
rect 144564 64228 144570 64230
rect 245653 64227 245719 64230
rect 164918 64092 164924 64156
rect 164988 64154 164994 64156
rect 511993 64154 512059 64157
rect 164988 64152 512059 64154
rect 164988 64096 511998 64152
rect 512054 64096 512059 64152
rect 164988 64094 512059 64096
rect 164988 64092 164994 64094
rect 511993 64091 512059 64094
rect 145230 62868 145236 62932
rect 145300 62930 145306 62932
rect 263593 62930 263659 62933
rect 145300 62928 263659 62930
rect 145300 62872 263598 62928
rect 263654 62872 263659 62928
rect 145300 62870 263659 62872
rect 145300 62868 145306 62870
rect 263593 62867 263659 62870
rect 170438 62732 170444 62796
rect 170508 62794 170514 62796
rect 575473 62794 575539 62797
rect 170508 62792 575539 62794
rect 170508 62736 575478 62792
rect 575534 62736 575539 62792
rect 170508 62734 575539 62736
rect 170508 62732 170514 62734
rect 575473 62731 575539 62734
rect 143022 61372 143028 61436
rect 143092 61434 143098 61436
rect 227713 61434 227779 61437
rect 143092 61432 227779 61434
rect 143092 61376 227718 61432
rect 227774 61376 227779 61432
rect 143092 61374 227779 61376
rect 143092 61372 143098 61374
rect 227713 61371 227779 61374
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3049 58578 3115 58581
rect -960 58576 3115 58578
rect -960 58520 3054 58576
rect 3110 58520 3115 58576
rect -960 58518 3115 58520
rect -960 58428 480 58518
rect 3049 58515 3115 58518
rect 170622 58516 170628 58580
rect 170692 58578 170698 58580
rect 578233 58578 578299 58581
rect 170692 58576 578299 58578
rect 170692 58520 578238 58576
rect 578294 58520 578299 58576
rect 170692 58518 578299 58520
rect 170692 58516 170698 58518
rect 578233 58515 578299 58518
rect 149646 55932 149652 55996
rect 149716 55994 149722 55996
rect 316033 55994 316099 55997
rect 149716 55992 316099 55994
rect 149716 55936 316038 55992
rect 316094 55936 316099 55992
rect 149716 55934 316099 55936
rect 149716 55932 149722 55934
rect 316033 55931 316099 55934
rect 155718 55796 155724 55860
rect 155788 55858 155794 55860
rect 387793 55858 387859 55861
rect 155788 55856 387859 55858
rect 155788 55800 387798 55856
rect 387854 55800 387859 55856
rect 155788 55798 387859 55800
rect 155788 55796 155794 55798
rect 387793 55795 387859 55798
rect 163446 53076 163452 53140
rect 163516 53138 163522 53140
rect 494053 53138 494119 53141
rect 163516 53136 494119 53138
rect 163516 53080 494058 53136
rect 494114 53080 494119 53136
rect 163516 53078 494119 53080
rect 163516 53076 163522 53078
rect 494053 53075 494119 53078
rect 145414 51988 145420 52052
rect 145484 52050 145490 52052
rect 266353 52050 266419 52053
rect 145484 52048 266419 52050
rect 145484 51992 266358 52048
rect 266414 51992 266419 52048
rect 145484 51990 266419 51992
rect 145484 51988 145490 51990
rect 266353 51987 266419 51990
rect 151302 51852 151308 51916
rect 151372 51914 151378 51916
rect 333973 51914 334039 51917
rect 151372 51912 334039 51914
rect 151372 51856 333978 51912
rect 334034 51856 334039 51912
rect 151372 51854 334039 51856
rect 151372 51852 151378 51854
rect 333973 51851 334039 51854
rect 153878 51716 153884 51780
rect 153948 51778 153954 51780
rect 369853 51778 369919 51781
rect 153948 51776 369919 51778
rect 153948 51720 369858 51776
rect 369914 51720 369919 51776
rect 153948 51718 369919 51720
rect 153948 51716 153954 51718
rect 369853 51715 369919 51718
rect 165102 50220 165108 50284
rect 165172 50282 165178 50284
rect 514753 50282 514819 50285
rect 165172 50280 514819 50282
rect 165172 50224 514758 50280
rect 514814 50224 514819 50280
rect 165172 50222 514819 50224
rect 165172 50220 165178 50222
rect 514753 50219 514819 50222
rect 157926 48860 157932 48924
rect 157996 48922 158002 48924
rect 423673 48922 423739 48925
rect 157996 48920 423739 48922
rect 157996 48864 423678 48920
rect 423734 48864 423739 48920
rect 157996 48862 423739 48864
rect 157996 48860 158002 48862
rect 423673 48859 423739 48862
rect 140446 47772 140452 47836
rect 140516 47834 140522 47836
rect 191833 47834 191899 47837
rect 140516 47832 191899 47834
rect 140516 47776 191838 47832
rect 191894 47776 191899 47832
rect 140516 47774 191899 47776
rect 140516 47772 140522 47774
rect 191833 47771 191899 47774
rect 152774 47636 152780 47700
rect 152844 47698 152850 47700
rect 351913 47698 351979 47701
rect 152844 47696 351979 47698
rect 152844 47640 351918 47696
rect 351974 47640 351979 47696
rect 152844 47638 351979 47640
rect 152844 47636 152850 47638
rect 351913 47635 351979 47638
rect 156822 47500 156828 47564
rect 156892 47562 156898 47564
rect 405733 47562 405799 47565
rect 156892 47560 405799 47562
rect 156892 47504 405738 47560
rect 405794 47504 405799 47560
rect 156892 47502 405799 47504
rect 156892 47500 156898 47502
rect 405733 47499 405799 47502
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 167678 46140 167684 46204
rect 167748 46202 167754 46204
rect 547873 46202 547939 46205
rect 167748 46200 547939 46202
rect 167748 46144 547878 46200
rect 547934 46144 547939 46200
rect 583520 46188 584960 46278
rect 167748 46142 547939 46144
rect 167748 46140 167754 46142
rect 547873 46139 547939 46142
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 74533 44842 74599 44845
rect 131430 44842 131436 44844
rect 74533 44840 131436 44842
rect 74533 44784 74538 44840
rect 74594 44784 131436 44840
rect 74533 44782 131436 44784
rect 74533 44779 74599 44782
rect 131430 44780 131436 44782
rect 131500 44780 131506 44844
rect 137686 43420 137692 43484
rect 137756 43482 137762 43484
rect 152457 43482 152523 43485
rect 137756 43480 152523 43482
rect 137756 43424 152462 43480
rect 152518 43424 152523 43480
rect 137756 43422 152523 43424
rect 137756 43420 137762 43422
rect 152457 43419 152523 43422
rect 163630 43420 163636 43484
rect 163700 43482 163706 43484
rect 495433 43482 495499 43485
rect 163700 43480 495499 43482
rect 163700 43424 495438 43480
rect 495494 43424 495499 43480
rect 163700 43422 495499 43424
rect 163700 43420 163706 43422
rect 495433 43419 495499 43422
rect 149830 42060 149836 42124
rect 149900 42122 149906 42124
rect 316125 42122 316191 42125
rect 149900 42120 316191 42122
rect 149900 42064 316130 42120
rect 316186 42064 316191 42120
rect 149900 42062 316191 42064
rect 149900 42060 149906 42062
rect 316125 42059 316191 42062
rect 145598 39204 145604 39268
rect 145668 39266 145674 39268
rect 264973 39266 265039 39269
rect 145668 39264 265039 39266
rect 145668 39208 264978 39264
rect 265034 39208 265039 39264
rect 145668 39206 265039 39208
rect 145668 39204 145674 39206
rect 264973 39203 265039 39206
rect 151486 35260 151492 35324
rect 151556 35322 151562 35324
rect 336733 35322 336799 35325
rect 151556 35320 336799 35322
rect 151556 35264 336738 35320
rect 336794 35264 336799 35320
rect 151556 35262 336799 35264
rect 151556 35260 151562 35262
rect 336733 35259 336799 35262
rect 152406 35124 152412 35188
rect 152476 35186 152482 35188
rect 350533 35186 350599 35189
rect 152476 35184 350599 35186
rect 152476 35128 350538 35184
rect 350594 35128 350599 35184
rect 152476 35126 350599 35128
rect 152476 35124 152482 35126
rect 350533 35123 350599 35126
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect 143206 32676 143212 32740
rect 143276 32738 143282 32740
rect 226425 32738 226491 32741
rect 143276 32736 226491 32738
rect 143276 32680 226430 32736
rect 226486 32680 226491 32736
rect 143276 32678 226491 32680
rect 143276 32676 143282 32678
rect 226425 32675 226491 32678
rect -960 32466 480 32556
rect 167862 32540 167868 32604
rect 167932 32602 167938 32604
rect 546493 32602 546559 32605
rect 167932 32600 546559 32602
rect 167932 32544 546498 32600
rect 546554 32544 546559 32600
rect 167932 32542 546559 32544
rect 167932 32540 167938 32542
rect 546493 32539 546559 32542
rect 3141 32466 3207 32469
rect -960 32464 3207 32466
rect -960 32408 3146 32464
rect 3202 32408 3207 32464
rect -960 32406 3207 32408
rect -960 32316 480 32406
rect 3141 32403 3207 32406
rect 169334 32404 169340 32468
rect 169404 32466 169410 32468
rect 567193 32466 567259 32469
rect 169404 32464 567259 32466
rect 169404 32408 567198 32464
rect 567254 32408 567259 32464
rect 169404 32406 567259 32408
rect 169404 32404 169410 32406
rect 567193 32403 567259 32406
rect 158846 31044 158852 31108
rect 158916 31106 158922 31108
rect 441613 31106 441679 31109
rect 158916 31104 441679 31106
rect 158916 31048 441618 31104
rect 441674 31048 441679 31104
rect 158916 31046 441679 31048
rect 158916 31044 158922 31046
rect 441613 31043 441679 31046
rect 161054 30908 161060 30972
rect 161124 30970 161130 30972
rect 456793 30970 456859 30973
rect 161124 30968 456859 30970
rect 161124 30912 456798 30968
rect 456854 30912 456859 30968
rect 161124 30910 456859 30912
rect 161124 30908 161130 30910
rect 456793 30907 456859 30910
rect 166390 28188 166396 28252
rect 166460 28250 166466 28252
rect 531313 28250 531379 28253
rect 166460 28248 531379 28250
rect 166460 28192 531318 28248
rect 531374 28192 531379 28248
rect 166460 28190 531379 28192
rect 166460 28188 166466 28190
rect 531313 28187 531379 28190
rect 140078 26964 140084 27028
rect 140148 27026 140154 27028
rect 193305 27026 193371 27029
rect 140148 27024 193371 27026
rect 140148 26968 193310 27024
rect 193366 26968 193371 27024
rect 140148 26966 193371 26968
rect 140148 26964 140154 26966
rect 193305 26963 193371 26966
rect 150014 26828 150020 26892
rect 150084 26890 150090 26892
rect 317413 26890 317479 26893
rect 150084 26888 317479 26890
rect 150084 26832 317418 26888
rect 317474 26832 317479 26888
rect 150084 26830 317479 26832
rect 150084 26828 150090 26830
rect 317413 26827 317479 26830
rect 19333 25530 19399 25533
rect 127382 25530 127388 25532
rect 19333 25528 127388 25530
rect 19333 25472 19338 25528
rect 19394 25472 127388 25528
rect 19333 25470 127388 25472
rect 19333 25467 19399 25470
rect 127382 25468 127388 25470
rect 127452 25468 127458 25532
rect 166574 24108 166580 24172
rect 166644 24170 166650 24172
rect 531405 24170 531471 24173
rect 166644 24168 531471 24170
rect 166644 24112 531410 24168
rect 531466 24112 531471 24168
rect 166644 24110 531471 24112
rect 166644 24108 166650 24110
rect 531405 24107 531471 24110
rect 170806 22612 170812 22676
rect 170876 22674 170882 22676
rect 582373 22674 582439 22677
rect 170876 22672 582439 22674
rect 170876 22616 582378 22672
rect 582434 22616 582439 22672
rect 170876 22614 582439 22616
rect 170876 22612 170882 22614
rect 582373 22611 582439 22614
rect 154062 21524 154068 21588
rect 154132 21586 154138 21588
rect 372613 21586 372679 21589
rect 154132 21584 372679 21586
rect 154132 21528 372618 21584
rect 372674 21528 372679 21584
rect 154132 21526 372679 21528
rect 154132 21524 154138 21526
rect 372613 21523 372679 21526
rect 159030 21388 159036 21452
rect 159100 21450 159106 21452
rect 442993 21450 443059 21453
rect 159100 21448 443059 21450
rect 159100 21392 442998 21448
rect 443054 21392 443059 21448
rect 159100 21390 443059 21392
rect 159100 21388 159106 21390
rect 442993 21387 443059 21390
rect 165286 21252 165292 21316
rect 165356 21314 165362 21316
rect 513373 21314 513439 21317
rect 165356 21312 513439 21314
rect 165356 21256 513378 21312
rect 513434 21256 513439 21312
rect 165356 21254 513439 21256
rect 165356 21252 165362 21254
rect 513373 21251 513439 21254
rect 144126 20028 144132 20092
rect 144196 20090 144202 20092
rect 248413 20090 248479 20093
rect 144196 20088 248479 20090
rect 144196 20032 248418 20088
rect 248474 20032 248479 20088
rect 144196 20030 248479 20032
rect 144196 20028 144202 20030
rect 248413 20027 248479 20030
rect 158110 19892 158116 19956
rect 158180 19954 158186 19956
rect 422293 19954 422359 19957
rect 158180 19952 422359 19954
rect 158180 19896 422298 19952
rect 422354 19896 422359 19952
rect 158180 19894 422359 19896
rect 158180 19892 158186 19894
rect 422293 19891 422359 19894
rect 579613 19818 579679 19821
rect 583520 19818 584960 19908
rect 579613 19816 584960 19818
rect 579613 19760 579618 19816
rect 579674 19760 584960 19816
rect 579613 19758 584960 19760
rect 579613 19755 579679 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3325 19410 3391 19413
rect -960 19408 3391 19410
rect -960 19352 3330 19408
rect 3386 19352 3391 19408
rect -960 19350 3391 19352
rect -960 19260 480 19350
rect 3325 19347 3391 19350
rect 157006 18532 157012 18596
rect 157076 18594 157082 18596
rect 407113 18594 407179 18597
rect 157076 18592 407179 18594
rect 157076 18536 407118 18592
rect 407174 18536 407179 18592
rect 157076 18534 407179 18536
rect 157076 18532 157082 18534
rect 407113 18531 407179 18534
rect 140998 17308 141004 17372
rect 141068 17370 141074 17372
rect 212533 17370 212599 17373
rect 141068 17368 212599 17370
rect 141068 17312 212538 17368
rect 212594 17312 212599 17368
rect 141068 17310 212599 17312
rect 141068 17308 141074 17310
rect 212533 17307 212599 17310
rect 148542 17172 148548 17236
rect 148612 17234 148618 17236
rect 300853 17234 300919 17237
rect 148612 17232 300919 17234
rect 148612 17176 300858 17232
rect 300914 17176 300919 17232
rect 148612 17174 300919 17176
rect 148612 17172 148618 17174
rect 300853 17171 300919 17174
rect 154246 15812 154252 15876
rect 154316 15874 154322 15876
rect 365805 15874 365871 15877
rect 154316 15872 365871 15874
rect 154316 15816 365810 15872
rect 365866 15816 365871 15872
rect 154316 15814 365871 15816
rect 154316 15812 154322 15814
rect 365805 15811 365871 15814
rect 165470 14452 165476 14516
rect 165540 14514 165546 14516
rect 511257 14514 511323 14517
rect 165540 14512 511323 14514
rect 165540 14456 511262 14512
rect 511318 14456 511323 14512
rect 165540 14454 511323 14456
rect 165540 14452 165546 14454
rect 511257 14451 511323 14454
rect 143390 13228 143396 13292
rect 143460 13290 143466 13292
rect 229369 13290 229435 13293
rect 143460 13288 229435 13290
rect 143460 13232 229374 13288
rect 229430 13232 229435 13288
rect 143460 13230 229435 13232
rect 143460 13228 143466 13230
rect 229369 13227 229435 13230
rect 154430 13092 154436 13156
rect 154500 13154 154506 13156
rect 371233 13154 371299 13157
rect 154500 13152 371299 13154
rect 154500 13096 371238 13152
rect 371294 13096 371299 13152
rect 154500 13094 371299 13096
rect 154500 13092 154506 13094
rect 371233 13091 371299 13094
rect 166758 12956 166764 13020
rect 166828 13018 166834 13020
rect 528553 13018 528619 13021
rect 166828 13016 528619 13018
rect 166828 12960 528558 13016
rect 528614 12960 528619 13016
rect 166828 12958 528619 12960
rect 166828 12956 166834 12958
rect 528553 12955 528619 12958
rect 151670 11732 151676 11796
rect 151740 11794 151746 11796
rect 336273 11794 336339 11797
rect 151740 11792 336339 11794
rect 151740 11736 336278 11792
rect 336334 11736 336339 11792
rect 151740 11734 336339 11736
rect 151740 11732 151746 11734
rect 336273 11731 336339 11734
rect 158294 11596 158300 11660
rect 158364 11658 158370 11660
rect 423765 11658 423831 11661
rect 158364 11656 423831 11658
rect 158364 11600 423770 11656
rect 423826 11600 423831 11656
rect 158364 11598 423831 11600
rect 158364 11596 158370 11598
rect 423765 11595 423831 11598
rect 110505 10298 110571 10301
rect 134006 10298 134012 10300
rect 110505 10296 134012 10298
rect 110505 10240 110510 10296
rect 110566 10240 134012 10296
rect 110505 10238 134012 10240
rect 110505 10235 110571 10238
rect 134006 10236 134012 10238
rect 134076 10236 134082 10300
rect 158478 10236 158484 10300
rect 158548 10298 158554 10300
rect 420913 10298 420979 10301
rect 158548 10296 420979 10298
rect 158548 10240 420918 10296
rect 420974 10240 420979 10296
rect 158548 10238 420979 10240
rect 158548 10236 158554 10238
rect 420913 10235 420979 10238
rect 147254 9556 147260 9620
rect 147324 9618 147330 9620
rect 279509 9618 279575 9621
rect 147324 9616 279575 9618
rect 147324 9560 279514 9616
rect 279570 9560 279575 9616
rect 147324 9558 279575 9560
rect 147324 9556 147330 9558
rect 279509 9555 279575 9558
rect 133638 9420 133644 9484
rect 133708 9482 133714 9484
rect 280705 9482 280771 9485
rect 133708 9480 280771 9482
rect 133708 9424 280710 9480
rect 280766 9424 280771 9480
rect 133708 9422 280771 9424
rect 133708 9420 133714 9422
rect 280705 9419 280771 9422
rect 156638 9284 156644 9348
rect 156708 9346 156714 9348
rect 407205 9346 407271 9349
rect 156708 9344 407271 9346
rect 156708 9288 407210 9344
rect 407266 9288 407271 9344
rect 156708 9286 407271 9288
rect 156708 9284 156714 9286
rect 407205 9283 407271 9286
rect 92749 9210 92815 9213
rect 133086 9210 133092 9212
rect 92749 9208 133092 9210
rect 92749 9152 92754 9208
rect 92810 9152 133092 9208
rect 92749 9150 133092 9152
rect 92749 9147 92815 9150
rect 133086 9148 133092 9150
rect 133156 9148 133162 9212
rect 160686 9148 160692 9212
rect 160756 9210 160762 9212
rect 459185 9210 459251 9213
rect 160756 9208 459251 9210
rect 160756 9152 459190 9208
rect 459246 9152 459251 9208
rect 160756 9150 459251 9152
rect 160756 9148 160762 9150
rect 459185 9147 459251 9150
rect 59629 9074 59695 9077
rect 129958 9074 129964 9076
rect 59629 9072 129964 9074
rect 59629 9016 59634 9072
rect 59690 9016 129964 9072
rect 59629 9014 129964 9016
rect 59629 9011 59695 9014
rect 129958 9012 129964 9014
rect 130028 9012 130034 9076
rect 162526 9012 162532 9076
rect 162596 9074 162602 9076
rect 474549 9074 474615 9077
rect 162596 9072 474615 9074
rect 162596 9016 474554 9072
rect 474610 9016 474615 9072
rect 162596 9014 474615 9016
rect 162596 9012 162602 9014
rect 474549 9011 474615 9014
rect 57237 8938 57303 8941
rect 129774 8938 129780 8940
rect 57237 8936 129780 8938
rect 57237 8880 57242 8936
rect 57298 8880 129780 8936
rect 57237 8878 129780 8880
rect 57237 8875 57303 8878
rect 129774 8876 129780 8878
rect 129844 8876 129850 8940
rect 162342 8876 162348 8940
rect 162412 8938 162418 8940
rect 478137 8938 478203 8941
rect 162412 8936 478203 8938
rect 162412 8880 478142 8936
rect 478198 8880 478203 8936
rect 162412 8878 478203 8880
rect 162412 8876 162418 8878
rect 478137 8875 478203 8878
rect 109309 7714 109375 7717
rect 133822 7714 133828 7716
rect 109309 7712 133828 7714
rect 109309 7656 109314 7712
rect 109370 7656 133828 7712
rect 109309 7654 133828 7656
rect 109309 7651 109375 7654
rect 133822 7652 133828 7654
rect 133892 7652 133898 7716
rect 41873 7578 41939 7581
rect 128670 7578 128676 7580
rect 41873 7576 128676 7578
rect 41873 7520 41878 7576
rect 41934 7520 128676 7576
rect 41873 7518 128676 7520
rect 41873 7515 41939 7518
rect 128670 7516 128676 7518
rect 128740 7516 128746 7580
rect -960 6490 480 6580
rect 148910 6564 148916 6628
rect 148980 6626 148986 6628
rect 299657 6626 299723 6629
rect 148980 6624 299723 6626
rect 148980 6568 299662 6624
rect 299718 6568 299723 6624
rect 148980 6566 299723 6568
rect 148980 6564 148986 6566
rect 299657 6563 299723 6566
rect 580257 6626 580323 6629
rect 583520 6626 584960 6716
rect 580257 6624 584960 6626
rect 580257 6568 580262 6624
rect 580318 6568 584960 6624
rect 580257 6566 584960 6568
rect 580257 6563 580323 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 148726 6428 148732 6492
rect 148796 6490 148802 6492
rect 300761 6490 300827 6493
rect 148796 6488 300827 6490
rect 148796 6432 300766 6488
rect 300822 6432 300827 6488
rect 583520 6476 584960 6566
rect 148796 6430 300827 6432
rect 148796 6428 148802 6430
rect 300761 6427 300827 6430
rect 162158 6292 162164 6356
rect 162228 6354 162234 6356
rect 476941 6354 477007 6357
rect 162228 6352 477007 6354
rect 162228 6296 476946 6352
rect 477002 6296 477007 6352
rect 162228 6294 477007 6296
rect 162228 6292 162234 6294
rect 476941 6291 477007 6294
rect 137870 6156 137876 6220
rect 137940 6218 137946 6220
rect 158897 6218 158963 6221
rect 137940 6216 158963 6218
rect 137940 6160 158902 6216
rect 158958 6160 158963 6216
rect 137940 6158 158963 6160
rect 137940 6156 137946 6158
rect 158897 6155 158963 6158
rect 168046 6156 168052 6220
rect 168116 6218 168122 6220
rect 549069 6218 549135 6221
rect 168116 6216 549135 6218
rect 168116 6160 549074 6216
rect 549130 6160 549135 6216
rect 168116 6158 549135 6160
rect 168116 6156 168122 6158
rect 549069 6155 549135 6158
rect 4061 4858 4127 4861
rect 126094 4858 126100 4860
rect 4061 4856 126100 4858
rect 4061 4800 4066 4856
rect 4122 4800 126100 4856
rect 4061 4798 126100 4800
rect 4061 4795 4127 4798
rect 126094 4796 126100 4798
rect 126164 4796 126170 4860
rect 170990 4796 170996 4860
rect 171060 4858 171066 4860
rect 462221 4858 462287 4861
rect 171060 4856 462287 4858
rect 171060 4800 462226 4856
rect 462282 4800 462287 4856
rect 171060 4798 462287 4800
rect 171060 4796 171066 4798
rect 462221 4795 462287 4798
rect 136030 3844 136036 3908
rect 136100 3906 136106 3908
rect 176745 3906 176811 3909
rect 136100 3904 176811 3906
rect 136100 3848 176750 3904
rect 176806 3848 176811 3904
rect 136100 3846 176811 3848
rect 136100 3844 136106 3846
rect 176745 3843 176811 3846
rect 147070 3708 147076 3772
rect 147140 3770 147146 3772
rect 281901 3770 281967 3773
rect 147140 3768 281967 3770
rect 147140 3712 281906 3768
rect 281962 3712 281967 3768
rect 147140 3710 281967 3712
rect 147140 3708 147146 3710
rect 281901 3707 281967 3710
rect 136214 3572 136220 3636
rect 136284 3634 136290 3636
rect 147121 3634 147187 3637
rect 136284 3632 147187 3634
rect 136284 3576 147126 3632
rect 147182 3576 147187 3632
rect 136284 3574 147187 3576
rect 136284 3572 136290 3574
rect 147121 3571 147187 3574
rect 172094 3572 172100 3636
rect 172164 3634 172170 3636
rect 533705 3634 533771 3637
rect 172164 3632 533771 3634
rect 172164 3576 533710 3632
rect 533766 3576 533771 3632
rect 172164 3574 533771 3576
rect 172164 3572 172170 3574
rect 533705 3571 533771 3574
rect 136398 3436 136404 3500
rect 136468 3498 136474 3500
rect 156597 3498 156663 3501
rect 136468 3496 156663 3498
rect 136468 3440 156602 3496
rect 156658 3440 156663 3496
rect 136468 3438 156663 3440
rect 136468 3436 136474 3438
rect 156597 3435 156663 3438
rect 171910 3436 171916 3500
rect 171980 3498 171986 3500
rect 554957 3498 555023 3501
rect 171980 3496 555023 3498
rect 171980 3440 554962 3496
rect 555018 3440 555023 3496
rect 171980 3438 555023 3440
rect 171980 3436 171986 3438
rect 554957 3435 555023 3438
rect 135110 3300 135116 3364
rect 135180 3362 135186 3364
rect 161289 3362 161355 3365
rect 135180 3360 161355 3362
rect 135180 3304 161294 3360
rect 161350 3304 161355 3360
rect 135180 3302 161355 3304
rect 135180 3300 135186 3302
rect 161289 3299 161355 3302
rect 172278 3300 172284 3364
rect 172348 3362 172354 3364
rect 569125 3362 569191 3365
rect 172348 3360 569191 3362
rect 172348 3304 569130 3360
rect 569186 3304 569191 3360
rect 172348 3302 569191 3304
rect 172348 3300 172354 3302
rect 569125 3299 569191 3302
<< via3 >>
rect 144684 200636 144748 200700
rect 149836 196284 149900 196348
rect 151308 196012 151372 196076
rect 144684 195604 144748 195668
rect 148732 194712 148796 194716
rect 148732 194656 148782 194712
rect 148782 194656 148796 194712
rect 148732 194652 148796 194656
rect 143580 191744 143644 191808
rect 141740 191252 141804 191316
rect 151308 191254 151372 191318
rect 141924 190572 141988 190636
rect 148732 191040 148796 191044
rect 148732 190984 148782 191040
rect 148782 190984 148796 191040
rect 148732 190980 148796 190984
rect 149836 190632 149900 190636
rect 149836 190576 149850 190632
rect 149850 190576 149900 190632
rect 149836 190572 149900 190576
rect 140636 186900 140700 186964
rect 146156 180704 146220 180708
rect 146156 180648 146170 180704
rect 146170 180648 146220 180704
rect 146156 180644 146220 180648
rect 140452 179148 140516 179212
rect 142660 178800 142724 178804
rect 142660 178744 142666 178800
rect 142666 178744 142722 178800
rect 142722 178744 142724 178800
rect 142660 178740 142724 178744
rect 142660 176700 142724 176764
rect 142292 173844 142356 173908
rect 142660 173768 142724 173772
rect 142660 173712 142710 173768
rect 142710 173712 142724 173768
rect 142660 173708 142724 173712
rect 144132 173708 144196 173772
rect 142476 173572 142540 173636
rect 142108 171260 142172 171324
rect 142108 170852 142172 170916
rect 141740 166364 141804 166428
rect 141924 166228 141988 166292
rect 142108 162208 142172 162212
rect 142108 162152 142122 162208
rect 142122 162152 142172 162208
rect 142108 162148 142172 162152
rect 142292 143380 142356 143444
rect 142476 143244 142540 143308
rect 140452 143108 140516 143172
rect 144132 142972 144196 143036
rect 146156 142836 146220 142900
rect 140636 142700 140700 142764
rect 143580 142564 143644 142628
rect 142108 142428 142172 142492
rect 142660 142156 142724 142220
rect 172284 80412 172348 80476
rect 171548 80276 171612 80340
rect 159404 80140 159468 80204
rect 171916 80140 171980 80204
rect 125916 79906 125920 79932
rect 125920 79906 125976 79932
rect 125976 79906 125980 79932
rect 125916 79868 125980 79906
rect 127572 79868 127636 79932
rect 127388 79732 127452 79796
rect 128308 79906 128312 79932
rect 128312 79906 128368 79932
rect 128368 79906 128372 79932
rect 128308 79868 128372 79906
rect 128860 79868 128924 79932
rect 129044 79928 129108 79932
rect 129044 79872 129048 79928
rect 129048 79872 129104 79928
rect 129104 79872 129108 79928
rect 129044 79868 129108 79872
rect 129780 79868 129844 79932
rect 130700 79906 130704 79932
rect 130704 79906 130760 79932
rect 130760 79906 130764 79932
rect 130700 79868 130764 79906
rect 130148 79656 130212 79660
rect 130148 79600 130162 79656
rect 130162 79600 130212 79656
rect 130148 79596 130212 79600
rect 130516 79596 130580 79660
rect 131252 79928 131316 79932
rect 131252 79872 131256 79928
rect 131256 79872 131312 79928
rect 131312 79872 131316 79928
rect 131252 79868 131316 79872
rect 131620 79868 131684 79932
rect 131804 79928 131868 79932
rect 131804 79872 131808 79928
rect 131808 79872 131864 79928
rect 131864 79872 131868 79928
rect 131804 79868 131868 79872
rect 133092 79868 133156 79932
rect 133276 79732 133340 79796
rect 133828 79868 133892 79932
rect 135484 79906 135488 79932
rect 135488 79906 135544 79932
rect 135544 79906 135548 79932
rect 135484 79868 135548 79906
rect 135852 79868 135916 79932
rect 137692 79868 137756 79932
rect 138428 79868 138492 79932
rect 137876 79792 137940 79796
rect 137876 79736 137880 79792
rect 137880 79736 137936 79792
rect 137936 79736 137940 79792
rect 137876 79732 137940 79736
rect 138612 79732 138676 79796
rect 140268 79868 140332 79932
rect 141004 79868 141068 79932
rect 142660 79868 142724 79932
rect 143764 79868 143828 79932
rect 144316 79868 144380 79932
rect 140452 79792 140516 79796
rect 140452 79736 140456 79792
rect 140456 79736 140512 79792
rect 140512 79736 140516 79792
rect 140452 79732 140516 79736
rect 145604 79868 145668 79932
rect 146892 79928 146956 79932
rect 146892 79872 146896 79928
rect 146896 79872 146952 79928
rect 146952 79872 146956 79928
rect 145236 79732 145300 79796
rect 146892 79868 146956 79872
rect 147260 79928 147324 79932
rect 147260 79872 147264 79928
rect 147264 79872 147320 79928
rect 147320 79872 147324 79928
rect 147260 79868 147324 79872
rect 146524 79732 146588 79796
rect 146708 79792 146772 79796
rect 146708 79736 146712 79792
rect 146712 79736 146768 79792
rect 146768 79736 146772 79792
rect 146708 79732 146772 79736
rect 148364 79868 148428 79932
rect 148732 79868 148796 79932
rect 149836 79868 149900 79932
rect 151676 79928 151740 79932
rect 151676 79872 151680 79928
rect 151680 79872 151736 79928
rect 151736 79872 151740 79928
rect 151676 79868 151740 79872
rect 148548 79732 148612 79796
rect 150020 79732 150084 79796
rect 151860 79656 151924 79660
rect 151860 79600 151910 79656
rect 151910 79600 151924 79656
rect 151860 79596 151924 79600
rect 152964 79868 153028 79932
rect 152412 79732 152476 79796
rect 153700 79868 153764 79932
rect 153884 79868 153948 79932
rect 156828 79868 156892 79932
rect 158116 79868 158180 79932
rect 154068 79732 154132 79796
rect 154988 79732 155052 79796
rect 155908 79732 155972 79796
rect 156644 79732 156708 79796
rect 158484 79732 158548 79796
rect 160140 79868 160204 79932
rect 160692 79868 160756 79932
rect 161980 79928 162044 79932
rect 161980 79872 161984 79928
rect 161984 79872 162040 79928
rect 162040 79872 162044 79928
rect 161980 79868 162044 79872
rect 162164 79868 162228 79932
rect 163268 79868 163332 79932
rect 163452 79868 163516 79932
rect 164740 79868 164804 79932
rect 165476 79868 165540 79932
rect 159772 79732 159836 79796
rect 160876 79732 160940 79796
rect 162900 79792 162964 79796
rect 162900 79736 162904 79792
rect 162904 79736 162960 79792
rect 162960 79736 162964 79792
rect 162900 79732 162964 79736
rect 163636 79732 163700 79796
rect 165292 79732 165356 79796
rect 166212 79868 166276 79932
rect 166580 79732 166644 79796
rect 168052 79868 168116 79932
rect 168788 79928 168852 79932
rect 168788 79872 168792 79928
rect 168792 79872 168848 79928
rect 168848 79872 168852 79928
rect 168788 79868 168852 79872
rect 169524 79868 169588 79932
rect 170260 79928 170324 79932
rect 170260 79872 170264 79928
rect 170264 79872 170320 79928
rect 170320 79872 170324 79928
rect 170260 79868 170324 79872
rect 171318 79902 171382 79966
rect 167868 79732 167932 79796
rect 169340 79732 169404 79796
rect 171548 79868 171612 79932
rect 171732 79906 171736 79932
rect 171736 79906 171792 79932
rect 171792 79906 171796 79932
rect 171732 79868 171796 79906
rect 173020 79868 173084 79932
rect 173204 79906 173208 79932
rect 173208 79906 173264 79932
rect 173264 79906 173268 79932
rect 173204 79868 173268 79906
rect 170812 79792 170876 79796
rect 170812 79736 170816 79792
rect 170816 79736 170872 79792
rect 170872 79736 170876 79792
rect 170812 79732 170876 79736
rect 170996 79732 171060 79796
rect 171180 79732 171244 79796
rect 171916 79596 171980 79660
rect 172100 79596 172164 79660
rect 159404 79188 159468 79252
rect 173204 79052 173268 79116
rect 171180 78916 171244 78980
rect 172284 78916 172348 78980
rect 126100 78780 126164 78844
rect 129964 78780 130028 78844
rect 130516 78780 130580 78844
rect 151492 78780 151556 78844
rect 157012 78780 157076 78844
rect 125732 78704 125796 78708
rect 125732 78648 125746 78704
rect 125746 78648 125796 78704
rect 125732 78644 125796 78648
rect 127204 78704 127268 78708
rect 127204 78648 127254 78704
rect 127254 78648 127268 78704
rect 127204 78644 127268 78648
rect 130332 78644 130396 78708
rect 135852 78704 135916 78708
rect 135852 78648 135902 78704
rect 135902 78648 135916 78704
rect 135852 78644 135916 78648
rect 151308 78644 151372 78708
rect 154988 78704 155052 78708
rect 154988 78648 155038 78704
rect 155038 78648 155052 78704
rect 154988 78644 155052 78648
rect 159036 78644 159100 78708
rect 162900 78644 162964 78708
rect 173020 78644 173084 78708
rect 159772 78508 159836 78572
rect 172100 78508 172164 78572
rect 168788 78432 168852 78436
rect 168788 78376 168802 78432
rect 168802 78376 168852 78432
rect 168788 78372 168852 78376
rect 171364 78432 171428 78436
rect 171364 78376 171378 78432
rect 171378 78376 171428 78432
rect 171364 78372 171428 78376
rect 127572 78236 127636 78300
rect 158852 78236 158916 78300
rect 128308 78100 128372 78164
rect 128492 78100 128556 78164
rect 154252 78100 154316 78164
rect 171732 78100 171796 78164
rect 153700 77964 153764 78028
rect 157196 78024 157260 78028
rect 157196 77968 157210 78024
rect 157210 77968 157260 78024
rect 157196 77964 157260 77968
rect 157932 77964 157996 78028
rect 133644 77828 133708 77892
rect 154436 77888 154500 77892
rect 154436 77832 154450 77888
rect 154450 77832 154500 77888
rect 154436 77828 154500 77832
rect 158300 77828 158364 77892
rect 170996 77888 171060 77892
rect 170996 77832 171010 77888
rect 171010 77832 171060 77888
rect 170996 77828 171060 77832
rect 151860 77420 151924 77484
rect 170996 77420 171060 77484
rect 128676 77284 128740 77348
rect 152780 77284 152844 77348
rect 155724 77344 155788 77348
rect 155724 77288 155774 77344
rect 155774 77288 155788 77344
rect 155724 77284 155788 77288
rect 160140 77284 160204 77348
rect 172284 77284 172348 77348
rect 169524 77148 169588 77212
rect 136220 76876 136284 76940
rect 136036 76740 136100 76804
rect 144500 76740 144564 76804
rect 146708 76740 146772 76804
rect 131436 76664 131500 76668
rect 131436 76608 131450 76664
rect 131450 76608 131500 76664
rect 131436 76604 131500 76608
rect 131804 76604 131868 76668
rect 134012 76664 134076 76668
rect 134012 76608 134062 76664
rect 134062 76608 134076 76664
rect 134012 76604 134076 76608
rect 135116 76604 135180 76668
rect 138980 76664 139044 76668
rect 138980 76608 138994 76664
rect 138994 76608 139044 76664
rect 138980 76604 139044 76608
rect 140084 76604 140148 76668
rect 143212 76664 143276 76668
rect 143212 76608 143226 76664
rect 143226 76608 143276 76664
rect 143212 76604 143276 76608
rect 143396 76664 143460 76668
rect 143396 76608 143446 76664
rect 143446 76608 143460 76664
rect 143396 76604 143460 76608
rect 144316 76604 144380 76668
rect 145420 76604 145484 76668
rect 146892 76604 146956 76668
rect 148916 76664 148980 76668
rect 148916 76608 148930 76664
rect 148930 76608 148980 76664
rect 148916 76604 148980 76608
rect 155908 76604 155972 76668
rect 130700 76468 130764 76532
rect 136404 76468 136468 76532
rect 138428 76468 138492 76532
rect 143028 76468 143092 76532
rect 144132 76468 144196 76532
rect 146524 76468 146588 76532
rect 160876 76468 160940 76532
rect 161060 76528 161124 76532
rect 161060 76472 161110 76528
rect 161110 76472 161124 76528
rect 161060 76468 161124 76472
rect 161980 76468 162044 76532
rect 162532 76528 162596 76532
rect 162532 76472 162546 76528
rect 162546 76472 162596 76528
rect 162532 76468 162596 76472
rect 163268 76468 163332 76532
rect 164924 76468 164988 76532
rect 166764 76528 166828 76532
rect 166764 76472 166778 76528
rect 166778 76472 166828 76528
rect 166764 76468 166828 76472
rect 167684 76468 167748 76532
rect 142660 76332 142724 76396
rect 162348 76332 162412 76396
rect 165108 76332 165172 76396
rect 166396 76332 166460 76396
rect 170628 76120 170692 76124
rect 170628 76064 170642 76120
rect 170642 76064 170692 76120
rect 170628 76060 170692 76064
rect 129044 75924 129108 75988
rect 170260 75924 170324 75988
rect 170444 75984 170508 75988
rect 170444 75928 170458 75984
rect 170458 75928 170508 75984
rect 170444 75924 170508 75928
rect 157012 75516 157076 75580
rect 164740 75244 164804 75308
rect 131620 75108 131684 75172
rect 149652 75108 149716 75172
rect 147076 74972 147140 75036
rect 125916 74428 125980 74492
rect 148364 74428 148428 74492
rect 143764 74156 143828 74220
rect 128676 73748 128740 73812
rect 128860 72524 128924 72588
rect 125732 72388 125796 72452
rect 133276 69668 133340 69732
rect 130332 69532 130396 69596
rect 138980 69532 139044 69596
rect 130148 68308 130212 68372
rect 152596 68308 152660 68372
rect 127204 68172 127268 68236
rect 135300 68172 135364 68236
rect 166212 68172 166276 68236
rect 138612 66948 138676 67012
rect 140268 66812 140332 66876
rect 131252 65452 131316 65516
rect 144500 64228 144564 64292
rect 164924 64092 164988 64156
rect 145236 62868 145300 62932
rect 170444 62732 170508 62796
rect 143028 61372 143092 61436
rect 170628 58516 170692 58580
rect 149652 55932 149716 55996
rect 155724 55796 155788 55860
rect 163452 53076 163516 53140
rect 145420 51988 145484 52052
rect 151308 51852 151372 51916
rect 153884 51716 153948 51780
rect 165108 50220 165172 50284
rect 157932 48860 157996 48924
rect 140452 47772 140516 47836
rect 152780 47636 152844 47700
rect 156828 47500 156892 47564
rect 167684 46140 167748 46204
rect 131436 44780 131500 44844
rect 137692 43420 137756 43484
rect 163636 43420 163700 43484
rect 149836 42060 149900 42124
rect 145604 39204 145668 39268
rect 151492 35260 151556 35324
rect 152412 35124 152476 35188
rect 143212 32676 143276 32740
rect 167868 32540 167932 32604
rect 169340 32404 169404 32468
rect 158852 31044 158916 31108
rect 161060 30908 161124 30972
rect 166396 28188 166460 28252
rect 140084 26964 140148 27028
rect 150020 26828 150084 26892
rect 127388 25468 127452 25532
rect 166580 24108 166644 24172
rect 170812 22612 170876 22676
rect 154068 21524 154132 21588
rect 159036 21388 159100 21452
rect 165292 21252 165356 21316
rect 144132 20028 144196 20092
rect 158116 19892 158180 19956
rect 157012 18532 157076 18596
rect 141004 17308 141068 17372
rect 148548 17172 148612 17236
rect 154252 15812 154316 15876
rect 165476 14452 165540 14516
rect 143396 13228 143460 13292
rect 154436 13092 154500 13156
rect 166764 12956 166828 13020
rect 151676 11732 151740 11796
rect 158300 11596 158364 11660
rect 134012 10236 134076 10300
rect 158484 10236 158548 10300
rect 147260 9556 147324 9620
rect 133644 9420 133708 9484
rect 156644 9284 156708 9348
rect 133092 9148 133156 9212
rect 160692 9148 160756 9212
rect 129964 9012 130028 9076
rect 162532 9012 162596 9076
rect 129780 8876 129844 8940
rect 162348 8876 162412 8940
rect 133828 7652 133892 7716
rect 128676 7516 128740 7580
rect 148916 6564 148980 6628
rect 148732 6428 148796 6492
rect 162164 6292 162228 6356
rect 137876 6156 137940 6220
rect 168052 6156 168116 6220
rect 126100 4796 126164 4860
rect 170996 4796 171060 4860
rect 136036 3844 136100 3908
rect 147076 3708 147140 3772
rect 136220 3572 136284 3636
rect 172100 3572 172164 3636
rect 136404 3436 136468 3500
rect 171916 3436 171980 3500
rect 135116 3300 135180 3364
rect 172284 3300 172348 3364
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 682954 -8106 711002
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 -8106 682954
rect -8726 682634 -8106 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 -8106 682634
rect -8726 646954 -8106 682398
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 -8106 646954
rect -8726 646634 -8106 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 -8106 646634
rect -8726 610954 -8106 646398
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 -8106 610954
rect -8726 610634 -8106 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 -8106 610634
rect -8726 574954 -8106 610398
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 -8106 574954
rect -8726 574634 -8106 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 -8106 574634
rect -8726 538954 -8106 574398
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 -8106 538954
rect -8726 538634 -8106 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 -8106 538634
rect -8726 502954 -8106 538398
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 -8106 502954
rect -8726 502634 -8106 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 -8106 502634
rect -8726 466954 -8106 502398
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 -8106 466954
rect -8726 466634 -8106 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 -8106 466634
rect -8726 430954 -8106 466398
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 -8106 430954
rect -8726 430634 -8106 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 -8106 430634
rect -8726 394954 -8106 430398
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 -8106 394954
rect -8726 394634 -8106 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 -8106 394634
rect -8726 358954 -8106 394398
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 -8106 358954
rect -8726 358634 -8106 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 -8106 358634
rect -8726 322954 -8106 358398
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 -8106 322954
rect -8726 322634 -8106 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 -8106 322634
rect -8726 286954 -8106 322398
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 -8106 286954
rect -8726 286634 -8106 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 -8106 286634
rect -8726 250954 -8106 286398
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 -8106 250954
rect -8726 250634 -8106 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 -8106 250634
rect -8726 214954 -8106 250398
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 -8106 214954
rect -8726 214634 -8106 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 -8106 214634
rect -8726 178954 -8106 214398
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 -8106 178954
rect -8726 178634 -8106 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 -8106 178634
rect -8726 142954 -8106 178398
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 -8106 142954
rect -8726 142634 -8106 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 -8106 142634
rect -8726 106954 -8106 142398
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 -8106 106954
rect -8726 106634 -8106 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 -8106 106634
rect -8726 70954 -8106 106398
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 -8106 70954
rect -8726 70634 -8106 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 -8106 70634
rect -8726 34954 -8106 70398
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 -8106 34954
rect -8726 34634 -8106 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 -8106 34634
rect -8726 -7066 -8106 34398
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 678454 -7146 710042
rect -7766 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 -7146 678454
rect -7766 678134 -7146 678218
rect -7766 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 -7146 678134
rect -7766 642454 -7146 677898
rect -7766 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 -7146 642454
rect -7766 642134 -7146 642218
rect -7766 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 -7146 642134
rect -7766 606454 -7146 641898
rect -7766 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 -7146 606454
rect -7766 606134 -7146 606218
rect -7766 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 -7146 606134
rect -7766 570454 -7146 605898
rect -7766 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 -7146 570454
rect -7766 570134 -7146 570218
rect -7766 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 -7146 570134
rect -7766 534454 -7146 569898
rect -7766 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 -7146 534454
rect -7766 534134 -7146 534218
rect -7766 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 -7146 534134
rect -7766 498454 -7146 533898
rect -7766 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 -7146 498454
rect -7766 498134 -7146 498218
rect -7766 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 -7146 498134
rect -7766 462454 -7146 497898
rect -7766 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 -7146 462454
rect -7766 462134 -7146 462218
rect -7766 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 -7146 462134
rect -7766 426454 -7146 461898
rect -7766 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 -7146 426454
rect -7766 426134 -7146 426218
rect -7766 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 -7146 426134
rect -7766 390454 -7146 425898
rect -7766 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 -7146 390454
rect -7766 390134 -7146 390218
rect -7766 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 -7146 390134
rect -7766 354454 -7146 389898
rect -7766 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 -7146 354454
rect -7766 354134 -7146 354218
rect -7766 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 -7146 354134
rect -7766 318454 -7146 353898
rect -7766 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 -7146 318454
rect -7766 318134 -7146 318218
rect -7766 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 -7146 318134
rect -7766 282454 -7146 317898
rect -7766 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 -7146 282454
rect -7766 282134 -7146 282218
rect -7766 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 -7146 282134
rect -7766 246454 -7146 281898
rect -7766 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 -7146 246454
rect -7766 246134 -7146 246218
rect -7766 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 -7146 246134
rect -7766 210454 -7146 245898
rect -7766 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 -7146 210454
rect -7766 210134 -7146 210218
rect -7766 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 -7146 210134
rect -7766 174454 -7146 209898
rect -7766 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 -7146 174454
rect -7766 174134 -7146 174218
rect -7766 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 -7146 174134
rect -7766 138454 -7146 173898
rect -7766 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 -7146 138454
rect -7766 138134 -7146 138218
rect -7766 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 -7146 138134
rect -7766 102454 -7146 137898
rect -7766 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 -7146 102454
rect -7766 102134 -7146 102218
rect -7766 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 -7146 102134
rect -7766 66454 -7146 101898
rect -7766 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 -7146 66454
rect -7766 66134 -7146 66218
rect -7766 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 -7146 66134
rect -7766 30454 -7146 65898
rect -7766 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 -7146 30454
rect -7766 30134 -7146 30218
rect -7766 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 -7146 30134
rect -7766 -6106 -7146 29898
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 673954 -6186 709082
rect -6806 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 -6186 673954
rect -6806 673634 -6186 673718
rect -6806 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 -6186 673634
rect -6806 637954 -6186 673398
rect -6806 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 -6186 637954
rect -6806 637634 -6186 637718
rect -6806 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 -6186 637634
rect -6806 601954 -6186 637398
rect -6806 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 -6186 601954
rect -6806 601634 -6186 601718
rect -6806 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 -6186 601634
rect -6806 565954 -6186 601398
rect -6806 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 -6186 565954
rect -6806 565634 -6186 565718
rect -6806 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 -6186 565634
rect -6806 529954 -6186 565398
rect -6806 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 -6186 529954
rect -6806 529634 -6186 529718
rect -6806 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 -6186 529634
rect -6806 493954 -6186 529398
rect -6806 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 -6186 493954
rect -6806 493634 -6186 493718
rect -6806 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 -6186 493634
rect -6806 457954 -6186 493398
rect -6806 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 -6186 457954
rect -6806 457634 -6186 457718
rect -6806 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 -6186 457634
rect -6806 421954 -6186 457398
rect -6806 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 -6186 421954
rect -6806 421634 -6186 421718
rect -6806 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 -6186 421634
rect -6806 385954 -6186 421398
rect -6806 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 -6186 385954
rect -6806 385634 -6186 385718
rect -6806 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 -6186 385634
rect -6806 349954 -6186 385398
rect -6806 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 -6186 349954
rect -6806 349634 -6186 349718
rect -6806 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 -6186 349634
rect -6806 313954 -6186 349398
rect -6806 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 -6186 313954
rect -6806 313634 -6186 313718
rect -6806 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 -6186 313634
rect -6806 277954 -6186 313398
rect -6806 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 -6186 277954
rect -6806 277634 -6186 277718
rect -6806 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 -6186 277634
rect -6806 241954 -6186 277398
rect -6806 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 -6186 241954
rect -6806 241634 -6186 241718
rect -6806 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 -6186 241634
rect -6806 205954 -6186 241398
rect -6806 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 -6186 205954
rect -6806 205634 -6186 205718
rect -6806 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 -6186 205634
rect -6806 169954 -6186 205398
rect -6806 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 -6186 169954
rect -6806 169634 -6186 169718
rect -6806 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 -6186 169634
rect -6806 133954 -6186 169398
rect -6806 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 -6186 133954
rect -6806 133634 -6186 133718
rect -6806 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 -6186 133634
rect -6806 97954 -6186 133398
rect -6806 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 -6186 97954
rect -6806 97634 -6186 97718
rect -6806 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 -6186 97634
rect -6806 61954 -6186 97398
rect -6806 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 -6186 61954
rect -6806 61634 -6186 61718
rect -6806 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 -6186 61634
rect -6806 25954 -6186 61398
rect -6806 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 -6186 25954
rect -6806 25634 -6186 25718
rect -6806 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 -6186 25634
rect -6806 -5146 -6186 25398
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 669454 -5226 708122
rect -5846 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 -5226 669454
rect -5846 669134 -5226 669218
rect -5846 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 -5226 669134
rect -5846 633454 -5226 668898
rect -5846 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 -5226 633454
rect -5846 633134 -5226 633218
rect -5846 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 -5226 633134
rect -5846 597454 -5226 632898
rect -5846 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 -5226 597454
rect -5846 597134 -5226 597218
rect -5846 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 -5226 597134
rect -5846 561454 -5226 596898
rect -5846 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 -5226 561454
rect -5846 561134 -5226 561218
rect -5846 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 -5226 561134
rect -5846 525454 -5226 560898
rect -5846 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 -5226 525454
rect -5846 525134 -5226 525218
rect -5846 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 -5226 525134
rect -5846 489454 -5226 524898
rect -5846 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 -5226 489454
rect -5846 489134 -5226 489218
rect -5846 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 -5226 489134
rect -5846 453454 -5226 488898
rect -5846 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 -5226 453454
rect -5846 453134 -5226 453218
rect -5846 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 -5226 453134
rect -5846 417454 -5226 452898
rect -5846 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 -5226 417454
rect -5846 417134 -5226 417218
rect -5846 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 -5226 417134
rect -5846 381454 -5226 416898
rect -5846 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 -5226 381454
rect -5846 381134 -5226 381218
rect -5846 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 -5226 381134
rect -5846 345454 -5226 380898
rect -5846 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 -5226 345454
rect -5846 345134 -5226 345218
rect -5846 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 -5226 345134
rect -5846 309454 -5226 344898
rect -5846 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 -5226 309454
rect -5846 309134 -5226 309218
rect -5846 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 -5226 309134
rect -5846 273454 -5226 308898
rect -5846 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 -5226 273454
rect -5846 273134 -5226 273218
rect -5846 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 -5226 273134
rect -5846 237454 -5226 272898
rect -5846 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 -5226 237454
rect -5846 237134 -5226 237218
rect -5846 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 -5226 237134
rect -5846 201454 -5226 236898
rect -5846 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 -5226 201454
rect -5846 201134 -5226 201218
rect -5846 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 -5226 201134
rect -5846 165454 -5226 200898
rect -5846 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 -5226 165454
rect -5846 165134 -5226 165218
rect -5846 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 -5226 165134
rect -5846 129454 -5226 164898
rect -5846 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 -5226 129454
rect -5846 129134 -5226 129218
rect -5846 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 -5226 129134
rect -5846 93454 -5226 128898
rect -5846 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 -5226 93454
rect -5846 93134 -5226 93218
rect -5846 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 -5226 93134
rect -5846 57454 -5226 92898
rect -5846 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 -5226 57454
rect -5846 57134 -5226 57218
rect -5846 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 -5226 57134
rect -5846 21454 -5226 56898
rect -5846 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 -5226 21454
rect -5846 21134 -5226 21218
rect -5846 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 -5226 21134
rect -5846 -4186 -5226 20898
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 700954 -4266 707162
rect -4886 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 -4266 700954
rect -4886 700634 -4266 700718
rect -4886 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 -4266 700634
rect -4886 664954 -4266 700398
rect -4886 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 -4266 664954
rect -4886 664634 -4266 664718
rect -4886 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 -4266 664634
rect -4886 628954 -4266 664398
rect -4886 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 -4266 628954
rect -4886 628634 -4266 628718
rect -4886 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 -4266 628634
rect -4886 592954 -4266 628398
rect -4886 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 -4266 592954
rect -4886 592634 -4266 592718
rect -4886 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 -4266 592634
rect -4886 556954 -4266 592398
rect -4886 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 -4266 556954
rect -4886 556634 -4266 556718
rect -4886 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 -4266 556634
rect -4886 520954 -4266 556398
rect -4886 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 -4266 520954
rect -4886 520634 -4266 520718
rect -4886 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 -4266 520634
rect -4886 484954 -4266 520398
rect -4886 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 -4266 484954
rect -4886 484634 -4266 484718
rect -4886 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 -4266 484634
rect -4886 448954 -4266 484398
rect -4886 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 -4266 448954
rect -4886 448634 -4266 448718
rect -4886 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 -4266 448634
rect -4886 412954 -4266 448398
rect -4886 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 -4266 412954
rect -4886 412634 -4266 412718
rect -4886 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 -4266 412634
rect -4886 376954 -4266 412398
rect -4886 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 -4266 376954
rect -4886 376634 -4266 376718
rect -4886 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 -4266 376634
rect -4886 340954 -4266 376398
rect -4886 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 -4266 340954
rect -4886 340634 -4266 340718
rect -4886 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 -4266 340634
rect -4886 304954 -4266 340398
rect -4886 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 -4266 304954
rect -4886 304634 -4266 304718
rect -4886 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 -4266 304634
rect -4886 268954 -4266 304398
rect -4886 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 -4266 268954
rect -4886 268634 -4266 268718
rect -4886 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 -4266 268634
rect -4886 232954 -4266 268398
rect -4886 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 -4266 232954
rect -4886 232634 -4266 232718
rect -4886 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 -4266 232634
rect -4886 196954 -4266 232398
rect -4886 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 -4266 196954
rect -4886 196634 -4266 196718
rect -4886 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 -4266 196634
rect -4886 160954 -4266 196398
rect -4886 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 -4266 160954
rect -4886 160634 -4266 160718
rect -4886 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 -4266 160634
rect -4886 124954 -4266 160398
rect -4886 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 -4266 124954
rect -4886 124634 -4266 124718
rect -4886 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 -4266 124634
rect -4886 88954 -4266 124398
rect -4886 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 -4266 88954
rect -4886 88634 -4266 88718
rect -4886 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 -4266 88634
rect -4886 52954 -4266 88398
rect -4886 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 -4266 52954
rect -4886 52634 -4266 52718
rect -4886 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 -4266 52634
rect -4886 16954 -4266 52398
rect -4886 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 -4266 16954
rect -4886 16634 -4266 16718
rect -4886 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 -4266 16634
rect -4886 -3226 -4266 16398
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 696454 -3306 706202
rect -3926 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 -3306 696454
rect -3926 696134 -3306 696218
rect -3926 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 -3306 696134
rect -3926 660454 -3306 695898
rect -3926 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 -3306 660454
rect -3926 660134 -3306 660218
rect -3926 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 -3306 660134
rect -3926 624454 -3306 659898
rect -3926 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 -3306 624454
rect -3926 624134 -3306 624218
rect -3926 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 -3306 624134
rect -3926 588454 -3306 623898
rect -3926 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 -3306 588454
rect -3926 588134 -3306 588218
rect -3926 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 -3306 588134
rect -3926 552454 -3306 587898
rect -3926 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 -3306 552454
rect -3926 552134 -3306 552218
rect -3926 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 -3306 552134
rect -3926 516454 -3306 551898
rect -3926 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 -3306 516454
rect -3926 516134 -3306 516218
rect -3926 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 -3306 516134
rect -3926 480454 -3306 515898
rect -3926 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 -3306 480454
rect -3926 480134 -3306 480218
rect -3926 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 -3306 480134
rect -3926 444454 -3306 479898
rect -3926 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 -3306 444454
rect -3926 444134 -3306 444218
rect -3926 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 -3306 444134
rect -3926 408454 -3306 443898
rect -3926 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 -3306 408454
rect -3926 408134 -3306 408218
rect -3926 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 -3306 408134
rect -3926 372454 -3306 407898
rect -3926 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 -3306 372454
rect -3926 372134 -3306 372218
rect -3926 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 -3306 372134
rect -3926 336454 -3306 371898
rect -3926 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 -3306 336454
rect -3926 336134 -3306 336218
rect -3926 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 -3306 336134
rect -3926 300454 -3306 335898
rect -3926 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 -3306 300454
rect -3926 300134 -3306 300218
rect -3926 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 -3306 300134
rect -3926 264454 -3306 299898
rect -3926 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 -3306 264454
rect -3926 264134 -3306 264218
rect -3926 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 -3306 264134
rect -3926 228454 -3306 263898
rect -3926 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 -3306 228454
rect -3926 228134 -3306 228218
rect -3926 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 -3306 228134
rect -3926 192454 -3306 227898
rect -3926 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 -3306 192454
rect -3926 192134 -3306 192218
rect -3926 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 -3306 192134
rect -3926 156454 -3306 191898
rect -3926 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 -3306 156454
rect -3926 156134 -3306 156218
rect -3926 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 -3306 156134
rect -3926 120454 -3306 155898
rect -3926 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 -3306 120454
rect -3926 120134 -3306 120218
rect -3926 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 -3306 120134
rect -3926 84454 -3306 119898
rect -3926 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 -3306 84454
rect -3926 84134 -3306 84218
rect -3926 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 -3306 84134
rect -3926 48454 -3306 83898
rect -3926 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 -3306 48454
rect -3926 48134 -3306 48218
rect -3926 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 -3306 48134
rect -3926 12454 -3306 47898
rect -3926 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 -3306 12454
rect -3926 12134 -3306 12218
rect -3926 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 -3306 12134
rect -3926 -2266 -3306 11898
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691954 -2346 705242
rect -2966 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 -2346 691954
rect -2966 691634 -2346 691718
rect -2966 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 -2346 691634
rect -2966 655954 -2346 691398
rect -2966 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 -2346 655954
rect -2966 655634 -2346 655718
rect -2966 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 -2346 655634
rect -2966 619954 -2346 655398
rect -2966 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 -2346 619954
rect -2966 619634 -2346 619718
rect -2966 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 -2346 619634
rect -2966 583954 -2346 619398
rect -2966 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 -2346 583954
rect -2966 583634 -2346 583718
rect -2966 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 -2346 583634
rect -2966 547954 -2346 583398
rect -2966 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 -2346 547954
rect -2966 547634 -2346 547718
rect -2966 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 -2346 547634
rect -2966 511954 -2346 547398
rect -2966 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 -2346 511954
rect -2966 511634 -2346 511718
rect -2966 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 -2346 511634
rect -2966 475954 -2346 511398
rect -2966 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 -2346 475954
rect -2966 475634 -2346 475718
rect -2966 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 -2346 475634
rect -2966 439954 -2346 475398
rect -2966 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 -2346 439954
rect -2966 439634 -2346 439718
rect -2966 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 -2346 439634
rect -2966 403954 -2346 439398
rect -2966 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 -2346 403954
rect -2966 403634 -2346 403718
rect -2966 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 -2346 403634
rect -2966 367954 -2346 403398
rect -2966 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 -2346 367954
rect -2966 367634 -2346 367718
rect -2966 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 -2346 367634
rect -2966 331954 -2346 367398
rect -2966 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 -2346 331954
rect -2966 331634 -2346 331718
rect -2966 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 -2346 331634
rect -2966 295954 -2346 331398
rect -2966 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 -2346 295954
rect -2966 295634 -2346 295718
rect -2966 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 -2346 295634
rect -2966 259954 -2346 295398
rect -2966 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 -2346 259954
rect -2966 259634 -2346 259718
rect -2966 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 -2346 259634
rect -2966 223954 -2346 259398
rect -2966 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 -2346 223954
rect -2966 223634 -2346 223718
rect -2966 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 -2346 223634
rect -2966 187954 -2346 223398
rect -2966 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 -2346 187954
rect -2966 187634 -2346 187718
rect -2966 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 -2346 187634
rect -2966 151954 -2346 187398
rect -2966 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 -2346 151954
rect -2966 151634 -2346 151718
rect -2966 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 -2346 151634
rect -2966 115954 -2346 151398
rect -2966 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 -2346 115954
rect -2966 115634 -2346 115718
rect -2966 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 -2346 115634
rect -2966 79954 -2346 115398
rect -2966 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 -2346 79954
rect -2966 79634 -2346 79718
rect -2966 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 -2346 79634
rect -2966 43954 -2346 79398
rect -2966 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 -2346 43954
rect -2966 43634 -2346 43718
rect -2966 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 -2346 43634
rect -2966 7954 -2346 43398
rect -2966 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 -2346 7954
rect -2966 7634 -2346 7718
rect -2966 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 -2346 7634
rect -2966 -1306 -2346 7398
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 6294 705798 6914 711590
rect 6294 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 6914 705798
rect 6294 705478 6914 705562
rect 6294 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 6914 705478
rect 6294 691954 6914 705242
rect 6294 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 6914 691954
rect 6294 691634 6914 691718
rect 6294 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 6914 691634
rect 6294 655954 6914 691398
rect 6294 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 6914 655954
rect 6294 655634 6914 655718
rect 6294 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 6914 655634
rect 6294 619954 6914 655398
rect 6294 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 6914 619954
rect 6294 619634 6914 619718
rect 6294 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 6914 619634
rect 6294 583954 6914 619398
rect 6294 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 6914 583954
rect 6294 583634 6914 583718
rect 6294 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 6914 583634
rect 6294 547954 6914 583398
rect 6294 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 6914 547954
rect 6294 547634 6914 547718
rect 6294 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 6914 547634
rect 6294 511954 6914 547398
rect 6294 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 6914 511954
rect 6294 511634 6914 511718
rect 6294 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 6914 511634
rect 6294 475954 6914 511398
rect 6294 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 6914 475954
rect 6294 475634 6914 475718
rect 6294 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 6914 475634
rect 6294 439954 6914 475398
rect 6294 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 6914 439954
rect 6294 439634 6914 439718
rect 6294 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 6914 439634
rect 6294 403954 6914 439398
rect 6294 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 6914 403954
rect 6294 403634 6914 403718
rect 6294 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 6914 403634
rect 6294 367954 6914 403398
rect 6294 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 6914 367954
rect 6294 367634 6914 367718
rect 6294 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 6914 367634
rect 6294 331954 6914 367398
rect 6294 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 6914 331954
rect 6294 331634 6914 331718
rect 6294 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 6914 331634
rect 6294 295954 6914 331398
rect 6294 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 6914 295954
rect 6294 295634 6914 295718
rect 6294 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 6914 295634
rect 6294 259954 6914 295398
rect 6294 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 6914 259954
rect 6294 259634 6914 259718
rect 6294 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 6914 259634
rect 6294 223954 6914 259398
rect 6294 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 6914 223954
rect 6294 223634 6914 223718
rect 6294 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 6914 223634
rect 6294 187954 6914 223398
rect 6294 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 6914 187954
rect 6294 187634 6914 187718
rect 6294 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 6914 187634
rect 6294 151954 6914 187398
rect 6294 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 6914 151954
rect 6294 151634 6914 151718
rect 6294 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 6914 151634
rect 6294 115954 6914 151398
rect 6294 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 6914 115954
rect 6294 115634 6914 115718
rect 6294 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 6914 115634
rect 6294 79954 6914 115398
rect 6294 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 6914 79954
rect 6294 79634 6914 79718
rect 6294 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 6914 79634
rect 6294 43954 6914 79398
rect 6294 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 6914 43954
rect 6294 43634 6914 43718
rect 6294 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 6914 43634
rect 6294 7954 6914 43398
rect 6294 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 6914 7954
rect 6294 7634 6914 7718
rect 6294 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 6914 7634
rect 6294 -1306 6914 7398
rect 6294 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 6914 -1306
rect 6294 -1626 6914 -1542
rect 6294 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 6914 -1626
rect 6294 -7654 6914 -1862
rect 10794 706758 11414 711590
rect 10794 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 11414 706758
rect 10794 706438 11414 706522
rect 10794 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 11414 706438
rect 10794 696454 11414 706202
rect 10794 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 11414 696454
rect 10794 696134 11414 696218
rect 10794 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 11414 696134
rect 10794 660454 11414 695898
rect 10794 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 11414 660454
rect 10794 660134 11414 660218
rect 10794 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 11414 660134
rect 10794 624454 11414 659898
rect 10794 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 11414 624454
rect 10794 624134 11414 624218
rect 10794 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 11414 624134
rect 10794 588454 11414 623898
rect 10794 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 11414 588454
rect 10794 588134 11414 588218
rect 10794 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 11414 588134
rect 10794 552454 11414 587898
rect 10794 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 11414 552454
rect 10794 552134 11414 552218
rect 10794 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 11414 552134
rect 10794 516454 11414 551898
rect 10794 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 11414 516454
rect 10794 516134 11414 516218
rect 10794 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 11414 516134
rect 10794 480454 11414 515898
rect 10794 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 11414 480454
rect 10794 480134 11414 480218
rect 10794 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 11414 480134
rect 10794 444454 11414 479898
rect 10794 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 11414 444454
rect 10794 444134 11414 444218
rect 10794 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 11414 444134
rect 10794 408454 11414 443898
rect 10794 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 11414 408454
rect 10794 408134 11414 408218
rect 10794 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 11414 408134
rect 10794 372454 11414 407898
rect 10794 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 11414 372454
rect 10794 372134 11414 372218
rect 10794 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 11414 372134
rect 10794 336454 11414 371898
rect 10794 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 11414 336454
rect 10794 336134 11414 336218
rect 10794 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 11414 336134
rect 10794 300454 11414 335898
rect 10794 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 11414 300454
rect 10794 300134 11414 300218
rect 10794 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 11414 300134
rect 10794 264454 11414 299898
rect 10794 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 11414 264454
rect 10794 264134 11414 264218
rect 10794 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 11414 264134
rect 10794 228454 11414 263898
rect 10794 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 11414 228454
rect 10794 228134 11414 228218
rect 10794 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 11414 228134
rect 10794 192454 11414 227898
rect 10794 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 11414 192454
rect 10794 192134 11414 192218
rect 10794 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 11414 192134
rect 10794 156454 11414 191898
rect 10794 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 11414 156454
rect 10794 156134 11414 156218
rect 10794 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 11414 156134
rect 10794 120454 11414 155898
rect 10794 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 11414 120454
rect 10794 120134 11414 120218
rect 10794 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 11414 120134
rect 10794 84454 11414 119898
rect 10794 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 11414 84454
rect 10794 84134 11414 84218
rect 10794 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 11414 84134
rect 10794 48454 11414 83898
rect 10794 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 11414 48454
rect 10794 48134 11414 48218
rect 10794 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 11414 48134
rect 10794 12454 11414 47898
rect 10794 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 11414 12454
rect 10794 12134 11414 12218
rect 10794 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 11414 12134
rect 10794 -2266 11414 11898
rect 10794 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 11414 -2266
rect 10794 -2586 11414 -2502
rect 10794 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 11414 -2586
rect 10794 -7654 11414 -2822
rect 15294 707718 15914 711590
rect 15294 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 15914 707718
rect 15294 707398 15914 707482
rect 15294 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 15914 707398
rect 15294 700954 15914 707162
rect 15294 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 15914 700954
rect 15294 700634 15914 700718
rect 15294 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 15914 700634
rect 15294 664954 15914 700398
rect 15294 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 15914 664954
rect 15294 664634 15914 664718
rect 15294 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 15914 664634
rect 15294 628954 15914 664398
rect 15294 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 15914 628954
rect 15294 628634 15914 628718
rect 15294 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 15914 628634
rect 15294 592954 15914 628398
rect 15294 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 15914 592954
rect 15294 592634 15914 592718
rect 15294 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 15914 592634
rect 15294 556954 15914 592398
rect 15294 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 15914 556954
rect 15294 556634 15914 556718
rect 15294 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 15914 556634
rect 15294 520954 15914 556398
rect 15294 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 15914 520954
rect 15294 520634 15914 520718
rect 15294 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 15914 520634
rect 15294 484954 15914 520398
rect 15294 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 15914 484954
rect 15294 484634 15914 484718
rect 15294 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 15914 484634
rect 15294 448954 15914 484398
rect 15294 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 15914 448954
rect 15294 448634 15914 448718
rect 15294 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 15914 448634
rect 15294 412954 15914 448398
rect 15294 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 15914 412954
rect 15294 412634 15914 412718
rect 15294 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 15914 412634
rect 15294 376954 15914 412398
rect 15294 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 15914 376954
rect 15294 376634 15914 376718
rect 15294 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 15914 376634
rect 15294 340954 15914 376398
rect 15294 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 15914 340954
rect 15294 340634 15914 340718
rect 15294 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 15914 340634
rect 15294 304954 15914 340398
rect 15294 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 15914 304954
rect 15294 304634 15914 304718
rect 15294 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 15914 304634
rect 15294 268954 15914 304398
rect 15294 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 15914 268954
rect 15294 268634 15914 268718
rect 15294 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 15914 268634
rect 15294 232954 15914 268398
rect 15294 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 15914 232954
rect 15294 232634 15914 232718
rect 15294 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 15914 232634
rect 15294 196954 15914 232398
rect 15294 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 15914 196954
rect 15294 196634 15914 196718
rect 15294 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 15914 196634
rect 15294 160954 15914 196398
rect 15294 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 15914 160954
rect 15294 160634 15914 160718
rect 15294 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 15914 160634
rect 15294 124954 15914 160398
rect 15294 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 15914 124954
rect 15294 124634 15914 124718
rect 15294 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 15914 124634
rect 15294 88954 15914 124398
rect 15294 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 15914 88954
rect 15294 88634 15914 88718
rect 15294 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 15914 88634
rect 15294 52954 15914 88398
rect 15294 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 15914 52954
rect 15294 52634 15914 52718
rect 15294 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 15914 52634
rect 15294 16954 15914 52398
rect 15294 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 15914 16954
rect 15294 16634 15914 16718
rect 15294 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 15914 16634
rect 15294 -3226 15914 16398
rect 15294 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 15914 -3226
rect 15294 -3546 15914 -3462
rect 15294 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 15914 -3546
rect 15294 -7654 15914 -3782
rect 19794 708678 20414 711590
rect 19794 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 20414 708678
rect 19794 708358 20414 708442
rect 19794 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 20414 708358
rect 19794 669454 20414 708122
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -4186 20414 20898
rect 19794 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 20414 -4186
rect 19794 -4506 20414 -4422
rect 19794 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 20414 -4506
rect 19794 -7654 20414 -4742
rect 24294 709638 24914 711590
rect 24294 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 24914 709638
rect 24294 709318 24914 709402
rect 24294 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 24914 709318
rect 24294 673954 24914 709082
rect 24294 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 24914 673954
rect 24294 673634 24914 673718
rect 24294 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 24914 673634
rect 24294 637954 24914 673398
rect 24294 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 24914 637954
rect 24294 637634 24914 637718
rect 24294 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 24914 637634
rect 24294 601954 24914 637398
rect 24294 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 24914 601954
rect 24294 601634 24914 601718
rect 24294 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 24914 601634
rect 24294 565954 24914 601398
rect 24294 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 24914 565954
rect 24294 565634 24914 565718
rect 24294 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 24914 565634
rect 24294 529954 24914 565398
rect 24294 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 24914 529954
rect 24294 529634 24914 529718
rect 24294 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 24914 529634
rect 24294 493954 24914 529398
rect 24294 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 24914 493954
rect 24294 493634 24914 493718
rect 24294 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 24914 493634
rect 24294 457954 24914 493398
rect 24294 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 24914 457954
rect 24294 457634 24914 457718
rect 24294 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 24914 457634
rect 24294 421954 24914 457398
rect 24294 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 24914 421954
rect 24294 421634 24914 421718
rect 24294 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 24914 421634
rect 24294 385954 24914 421398
rect 24294 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 24914 385954
rect 24294 385634 24914 385718
rect 24294 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 24914 385634
rect 24294 349954 24914 385398
rect 24294 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 24914 349954
rect 24294 349634 24914 349718
rect 24294 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 24914 349634
rect 24294 313954 24914 349398
rect 24294 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 24914 313954
rect 24294 313634 24914 313718
rect 24294 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 24914 313634
rect 24294 277954 24914 313398
rect 24294 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 24914 277954
rect 24294 277634 24914 277718
rect 24294 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 24914 277634
rect 24294 241954 24914 277398
rect 24294 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 24914 241954
rect 24294 241634 24914 241718
rect 24294 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 24914 241634
rect 24294 205954 24914 241398
rect 24294 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 24914 205954
rect 24294 205634 24914 205718
rect 24294 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 24914 205634
rect 24294 169954 24914 205398
rect 24294 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 24914 169954
rect 24294 169634 24914 169718
rect 24294 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 24914 169634
rect 24294 133954 24914 169398
rect 24294 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 24914 133954
rect 24294 133634 24914 133718
rect 24294 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 24914 133634
rect 24294 97954 24914 133398
rect 24294 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 24914 97954
rect 24294 97634 24914 97718
rect 24294 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 24914 97634
rect 24294 61954 24914 97398
rect 24294 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 24914 61954
rect 24294 61634 24914 61718
rect 24294 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 24914 61634
rect 24294 25954 24914 61398
rect 24294 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 24914 25954
rect 24294 25634 24914 25718
rect 24294 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 24914 25634
rect 24294 -5146 24914 25398
rect 24294 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 24914 -5146
rect 24294 -5466 24914 -5382
rect 24294 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 24914 -5466
rect 24294 -7654 24914 -5702
rect 28794 710598 29414 711590
rect 28794 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 29414 710598
rect 28794 710278 29414 710362
rect 28794 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 29414 710278
rect 28794 678454 29414 710042
rect 28794 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 29414 678454
rect 28794 678134 29414 678218
rect 28794 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 29414 678134
rect 28794 642454 29414 677898
rect 28794 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 29414 642454
rect 28794 642134 29414 642218
rect 28794 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 29414 642134
rect 28794 606454 29414 641898
rect 28794 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 29414 606454
rect 28794 606134 29414 606218
rect 28794 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 29414 606134
rect 28794 570454 29414 605898
rect 28794 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 29414 570454
rect 28794 570134 29414 570218
rect 28794 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 29414 570134
rect 28794 534454 29414 569898
rect 28794 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 29414 534454
rect 28794 534134 29414 534218
rect 28794 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 29414 534134
rect 28794 498454 29414 533898
rect 28794 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 29414 498454
rect 28794 498134 29414 498218
rect 28794 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 29414 498134
rect 28794 462454 29414 497898
rect 28794 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 29414 462454
rect 28794 462134 29414 462218
rect 28794 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 29414 462134
rect 28794 426454 29414 461898
rect 28794 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 29414 426454
rect 28794 426134 29414 426218
rect 28794 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 29414 426134
rect 28794 390454 29414 425898
rect 28794 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 29414 390454
rect 28794 390134 29414 390218
rect 28794 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 29414 390134
rect 28794 354454 29414 389898
rect 28794 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 29414 354454
rect 28794 354134 29414 354218
rect 28794 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 29414 354134
rect 28794 318454 29414 353898
rect 28794 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 29414 318454
rect 28794 318134 29414 318218
rect 28794 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 29414 318134
rect 28794 282454 29414 317898
rect 28794 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 29414 282454
rect 28794 282134 29414 282218
rect 28794 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 29414 282134
rect 28794 246454 29414 281898
rect 28794 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 29414 246454
rect 28794 246134 29414 246218
rect 28794 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 29414 246134
rect 28794 210454 29414 245898
rect 28794 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 29414 210454
rect 28794 210134 29414 210218
rect 28794 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 29414 210134
rect 28794 174454 29414 209898
rect 28794 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 29414 174454
rect 28794 174134 29414 174218
rect 28794 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 29414 174134
rect 28794 138454 29414 173898
rect 28794 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 29414 138454
rect 28794 138134 29414 138218
rect 28794 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 29414 138134
rect 28794 102454 29414 137898
rect 28794 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 29414 102454
rect 28794 102134 29414 102218
rect 28794 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 29414 102134
rect 28794 66454 29414 101898
rect 28794 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 29414 66454
rect 28794 66134 29414 66218
rect 28794 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 29414 66134
rect 28794 30454 29414 65898
rect 28794 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 29414 30454
rect 28794 30134 29414 30218
rect 28794 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 29414 30134
rect 28794 -6106 29414 29898
rect 28794 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 29414 -6106
rect 28794 -6426 29414 -6342
rect 28794 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 29414 -6426
rect 28794 -7654 29414 -6662
rect 33294 711558 33914 711590
rect 33294 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 33914 711558
rect 33294 711238 33914 711322
rect 33294 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 33914 711238
rect 33294 682954 33914 711002
rect 33294 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 33914 682954
rect 33294 682634 33914 682718
rect 33294 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 33914 682634
rect 33294 646954 33914 682398
rect 33294 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 33914 646954
rect 33294 646634 33914 646718
rect 33294 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 33914 646634
rect 33294 610954 33914 646398
rect 33294 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 33914 610954
rect 33294 610634 33914 610718
rect 33294 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 33914 610634
rect 33294 574954 33914 610398
rect 33294 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 33914 574954
rect 33294 574634 33914 574718
rect 33294 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 33914 574634
rect 33294 538954 33914 574398
rect 33294 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 33914 538954
rect 33294 538634 33914 538718
rect 33294 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 33914 538634
rect 33294 502954 33914 538398
rect 33294 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 33914 502954
rect 33294 502634 33914 502718
rect 33294 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 33914 502634
rect 33294 466954 33914 502398
rect 33294 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 33914 466954
rect 33294 466634 33914 466718
rect 33294 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 33914 466634
rect 33294 430954 33914 466398
rect 33294 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 33914 430954
rect 33294 430634 33914 430718
rect 33294 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 33914 430634
rect 33294 394954 33914 430398
rect 33294 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 33914 394954
rect 33294 394634 33914 394718
rect 33294 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 33914 394634
rect 33294 358954 33914 394398
rect 33294 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 33914 358954
rect 33294 358634 33914 358718
rect 33294 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 33914 358634
rect 33294 322954 33914 358398
rect 33294 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 33914 322954
rect 33294 322634 33914 322718
rect 33294 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 33914 322634
rect 33294 286954 33914 322398
rect 33294 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 33914 286954
rect 33294 286634 33914 286718
rect 33294 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 33914 286634
rect 33294 250954 33914 286398
rect 33294 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 33914 250954
rect 33294 250634 33914 250718
rect 33294 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 33914 250634
rect 33294 214954 33914 250398
rect 33294 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 33914 214954
rect 33294 214634 33914 214718
rect 33294 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 33914 214634
rect 33294 178954 33914 214398
rect 33294 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 33914 178954
rect 33294 178634 33914 178718
rect 33294 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 33914 178634
rect 33294 142954 33914 178398
rect 33294 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 33914 142954
rect 33294 142634 33914 142718
rect 33294 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 33914 142634
rect 33294 106954 33914 142398
rect 33294 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 33914 106954
rect 33294 106634 33914 106718
rect 33294 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 33914 106634
rect 33294 70954 33914 106398
rect 33294 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 33914 70954
rect 33294 70634 33914 70718
rect 33294 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 33914 70634
rect 33294 34954 33914 70398
rect 33294 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 33914 34954
rect 33294 34634 33914 34718
rect 33294 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 33914 34634
rect 33294 -7066 33914 34398
rect 33294 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 33914 -7066
rect 33294 -7386 33914 -7302
rect 33294 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 33914 -7386
rect 33294 -7654 33914 -7622
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 42294 705798 42914 711590
rect 42294 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 42914 705798
rect 42294 705478 42914 705562
rect 42294 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 42914 705478
rect 42294 691954 42914 705242
rect 42294 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 42914 691954
rect 42294 691634 42914 691718
rect 42294 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 42914 691634
rect 42294 655954 42914 691398
rect 42294 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 42914 655954
rect 42294 655634 42914 655718
rect 42294 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 42914 655634
rect 42294 619954 42914 655398
rect 42294 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 42914 619954
rect 42294 619634 42914 619718
rect 42294 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 42914 619634
rect 42294 583954 42914 619398
rect 42294 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 42914 583954
rect 42294 583634 42914 583718
rect 42294 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 42914 583634
rect 42294 547954 42914 583398
rect 42294 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 42914 547954
rect 42294 547634 42914 547718
rect 42294 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 42914 547634
rect 42294 511954 42914 547398
rect 42294 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 42914 511954
rect 42294 511634 42914 511718
rect 42294 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 42914 511634
rect 42294 475954 42914 511398
rect 42294 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 42914 475954
rect 42294 475634 42914 475718
rect 42294 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 42914 475634
rect 42294 439954 42914 475398
rect 42294 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 42914 439954
rect 42294 439634 42914 439718
rect 42294 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 42914 439634
rect 42294 403954 42914 439398
rect 42294 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 42914 403954
rect 42294 403634 42914 403718
rect 42294 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 42914 403634
rect 42294 367954 42914 403398
rect 42294 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 42914 367954
rect 42294 367634 42914 367718
rect 42294 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 42914 367634
rect 42294 331954 42914 367398
rect 42294 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 42914 331954
rect 42294 331634 42914 331718
rect 42294 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 42914 331634
rect 42294 295954 42914 331398
rect 42294 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 42914 295954
rect 42294 295634 42914 295718
rect 42294 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 42914 295634
rect 42294 259954 42914 295398
rect 42294 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 42914 259954
rect 42294 259634 42914 259718
rect 42294 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 42914 259634
rect 42294 223954 42914 259398
rect 46794 706758 47414 711590
rect 46794 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 47414 706758
rect 46794 706438 47414 706522
rect 46794 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 47414 706438
rect 46794 696454 47414 706202
rect 46794 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 47414 696454
rect 46794 696134 47414 696218
rect 46794 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 47414 696134
rect 46794 660454 47414 695898
rect 46794 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 47414 660454
rect 46794 660134 47414 660218
rect 46794 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 47414 660134
rect 46794 624454 47414 659898
rect 46794 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 47414 624454
rect 46794 624134 47414 624218
rect 46794 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 47414 624134
rect 46794 588454 47414 623898
rect 46794 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 47414 588454
rect 46794 588134 47414 588218
rect 46794 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 47414 588134
rect 46794 552454 47414 587898
rect 46794 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 47414 552454
rect 46794 552134 47414 552218
rect 46794 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 47414 552134
rect 46794 516454 47414 551898
rect 46794 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 47414 516454
rect 46794 516134 47414 516218
rect 46794 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 47414 516134
rect 46794 480454 47414 515898
rect 46794 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 47414 480454
rect 46794 480134 47414 480218
rect 46794 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 47414 480134
rect 46794 444454 47414 479898
rect 46794 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 47414 444454
rect 46794 444134 47414 444218
rect 46794 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 47414 444134
rect 46794 408454 47414 443898
rect 46794 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 47414 408454
rect 46794 408134 47414 408218
rect 46794 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 47414 408134
rect 46794 372454 47414 407898
rect 46794 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 47414 372454
rect 46794 372134 47414 372218
rect 46794 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 47414 372134
rect 46794 336454 47414 371898
rect 46794 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 47414 336454
rect 46794 336134 47414 336218
rect 46794 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 47414 336134
rect 46794 300454 47414 335898
rect 46794 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 47414 300454
rect 46794 300134 47414 300218
rect 46794 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 47414 300134
rect 46794 264454 47414 299898
rect 46794 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 47414 264454
rect 46794 264134 47414 264218
rect 46794 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 47414 264134
rect 46794 244084 47414 263898
rect 51294 707718 51914 711590
rect 51294 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 51914 707718
rect 51294 707398 51914 707482
rect 51294 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 51914 707398
rect 51294 700954 51914 707162
rect 51294 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 51914 700954
rect 51294 700634 51914 700718
rect 51294 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 51914 700634
rect 51294 664954 51914 700398
rect 51294 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 51914 664954
rect 51294 664634 51914 664718
rect 51294 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 51914 664634
rect 51294 628954 51914 664398
rect 51294 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 51914 628954
rect 51294 628634 51914 628718
rect 51294 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 51914 628634
rect 51294 592954 51914 628398
rect 51294 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 51914 592954
rect 51294 592634 51914 592718
rect 51294 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 51914 592634
rect 51294 556954 51914 592398
rect 51294 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 51914 556954
rect 51294 556634 51914 556718
rect 51294 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 51914 556634
rect 51294 520954 51914 556398
rect 51294 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 51914 520954
rect 51294 520634 51914 520718
rect 51294 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 51914 520634
rect 51294 484954 51914 520398
rect 51294 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 51914 484954
rect 51294 484634 51914 484718
rect 51294 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 51914 484634
rect 51294 448954 51914 484398
rect 51294 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 51914 448954
rect 51294 448634 51914 448718
rect 51294 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 51914 448634
rect 51294 412954 51914 448398
rect 51294 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 51914 412954
rect 51294 412634 51914 412718
rect 51294 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 51914 412634
rect 51294 376954 51914 412398
rect 51294 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 51914 376954
rect 51294 376634 51914 376718
rect 51294 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 51914 376634
rect 51294 340954 51914 376398
rect 51294 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 51914 340954
rect 51294 340634 51914 340718
rect 51294 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 51914 340634
rect 51294 304954 51914 340398
rect 51294 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 51914 304954
rect 51294 304634 51914 304718
rect 51294 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 51914 304634
rect 51294 268954 51914 304398
rect 51294 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 51914 268954
rect 51294 268634 51914 268718
rect 51294 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 51914 268634
rect 51294 244084 51914 268398
rect 55794 708678 56414 711590
rect 55794 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 56414 708678
rect 55794 708358 56414 708442
rect 55794 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 56414 708358
rect 55794 669454 56414 708122
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 244084 56414 272898
rect 60294 709638 60914 711590
rect 60294 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 60914 709638
rect 60294 709318 60914 709402
rect 60294 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 60914 709318
rect 60294 673954 60914 709082
rect 60294 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 60914 673954
rect 60294 673634 60914 673718
rect 60294 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 60914 673634
rect 60294 637954 60914 673398
rect 60294 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 60914 637954
rect 60294 637634 60914 637718
rect 60294 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 60914 637634
rect 60294 601954 60914 637398
rect 60294 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 60914 601954
rect 60294 601634 60914 601718
rect 60294 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 60914 601634
rect 60294 565954 60914 601398
rect 60294 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 60914 565954
rect 60294 565634 60914 565718
rect 60294 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 60914 565634
rect 60294 529954 60914 565398
rect 60294 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 60914 529954
rect 60294 529634 60914 529718
rect 60294 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 60914 529634
rect 60294 493954 60914 529398
rect 60294 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 60914 493954
rect 60294 493634 60914 493718
rect 60294 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 60914 493634
rect 60294 457954 60914 493398
rect 60294 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 60914 457954
rect 60294 457634 60914 457718
rect 60294 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 60914 457634
rect 60294 421954 60914 457398
rect 60294 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 60914 421954
rect 60294 421634 60914 421718
rect 60294 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 60914 421634
rect 60294 385954 60914 421398
rect 60294 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 60914 385954
rect 60294 385634 60914 385718
rect 60294 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 60914 385634
rect 60294 349954 60914 385398
rect 60294 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 60914 349954
rect 60294 349634 60914 349718
rect 60294 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 60914 349634
rect 60294 313954 60914 349398
rect 60294 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 60914 313954
rect 60294 313634 60914 313718
rect 60294 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 60914 313634
rect 60294 277954 60914 313398
rect 60294 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 60914 277954
rect 60294 277634 60914 277718
rect 60294 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 60914 277634
rect 60294 244084 60914 277398
rect 64794 710598 65414 711590
rect 64794 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 65414 710598
rect 64794 710278 65414 710362
rect 64794 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 65414 710278
rect 64794 678454 65414 710042
rect 64794 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 65414 678454
rect 64794 678134 65414 678218
rect 64794 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 65414 678134
rect 64794 642454 65414 677898
rect 64794 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 65414 642454
rect 64794 642134 65414 642218
rect 64794 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 65414 642134
rect 64794 606454 65414 641898
rect 64794 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 65414 606454
rect 64794 606134 65414 606218
rect 64794 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 65414 606134
rect 64794 570454 65414 605898
rect 64794 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 65414 570454
rect 64794 570134 65414 570218
rect 64794 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 65414 570134
rect 64794 534454 65414 569898
rect 64794 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 65414 534454
rect 64794 534134 65414 534218
rect 64794 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 65414 534134
rect 64794 498454 65414 533898
rect 64794 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 65414 498454
rect 64794 498134 65414 498218
rect 64794 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 65414 498134
rect 64794 462454 65414 497898
rect 64794 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 65414 462454
rect 64794 462134 65414 462218
rect 64794 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 65414 462134
rect 64794 426454 65414 461898
rect 64794 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 65414 426454
rect 64794 426134 65414 426218
rect 64794 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 65414 426134
rect 64794 390454 65414 425898
rect 64794 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 65414 390454
rect 64794 390134 65414 390218
rect 64794 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 65414 390134
rect 64794 354454 65414 389898
rect 64794 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 65414 354454
rect 64794 354134 65414 354218
rect 64794 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 65414 354134
rect 64794 318454 65414 353898
rect 64794 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 65414 318454
rect 64794 318134 65414 318218
rect 64794 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 65414 318134
rect 64794 282454 65414 317898
rect 64794 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 65414 282454
rect 64794 282134 65414 282218
rect 64794 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 65414 282134
rect 64794 246454 65414 281898
rect 64794 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 65414 246454
rect 64794 246134 65414 246218
rect 64794 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 65414 246134
rect 64794 244084 65414 245898
rect 69294 711558 69914 711590
rect 69294 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 69914 711558
rect 69294 711238 69914 711322
rect 69294 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 69914 711238
rect 69294 682954 69914 711002
rect 69294 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 69914 682954
rect 69294 682634 69914 682718
rect 69294 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 69914 682634
rect 69294 646954 69914 682398
rect 69294 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 69914 646954
rect 69294 646634 69914 646718
rect 69294 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 69914 646634
rect 69294 610954 69914 646398
rect 69294 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 69914 610954
rect 69294 610634 69914 610718
rect 69294 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 69914 610634
rect 69294 574954 69914 610398
rect 69294 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 69914 574954
rect 69294 574634 69914 574718
rect 69294 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 69914 574634
rect 69294 538954 69914 574398
rect 69294 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 69914 538954
rect 69294 538634 69914 538718
rect 69294 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 69914 538634
rect 69294 502954 69914 538398
rect 69294 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 69914 502954
rect 69294 502634 69914 502718
rect 69294 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 69914 502634
rect 69294 466954 69914 502398
rect 69294 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 69914 466954
rect 69294 466634 69914 466718
rect 69294 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 69914 466634
rect 69294 430954 69914 466398
rect 69294 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 69914 430954
rect 69294 430634 69914 430718
rect 69294 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 69914 430634
rect 69294 394954 69914 430398
rect 69294 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 69914 394954
rect 69294 394634 69914 394718
rect 69294 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 69914 394634
rect 69294 358954 69914 394398
rect 69294 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 69914 358954
rect 69294 358634 69914 358718
rect 69294 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 69914 358634
rect 69294 322954 69914 358398
rect 69294 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 69914 322954
rect 69294 322634 69914 322718
rect 69294 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 69914 322634
rect 69294 286954 69914 322398
rect 69294 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 69914 286954
rect 69294 286634 69914 286718
rect 69294 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 69914 286634
rect 69294 250954 69914 286398
rect 69294 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 69914 250954
rect 69294 250634 69914 250718
rect 69294 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 69914 250634
rect 69294 244084 69914 250398
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 244084 74414 254898
rect 78294 705798 78914 711590
rect 78294 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 78914 705798
rect 78294 705478 78914 705562
rect 78294 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 78914 705478
rect 78294 691954 78914 705242
rect 78294 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 78914 691954
rect 78294 691634 78914 691718
rect 78294 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 78914 691634
rect 78294 655954 78914 691398
rect 78294 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 78914 655954
rect 78294 655634 78914 655718
rect 78294 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 78914 655634
rect 78294 619954 78914 655398
rect 78294 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 78914 619954
rect 78294 619634 78914 619718
rect 78294 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 78914 619634
rect 78294 583954 78914 619398
rect 78294 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 78914 583954
rect 78294 583634 78914 583718
rect 78294 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 78914 583634
rect 78294 547954 78914 583398
rect 78294 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 78914 547954
rect 78294 547634 78914 547718
rect 78294 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 78914 547634
rect 78294 511954 78914 547398
rect 78294 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 78914 511954
rect 78294 511634 78914 511718
rect 78294 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 78914 511634
rect 78294 475954 78914 511398
rect 78294 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 78914 475954
rect 78294 475634 78914 475718
rect 78294 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 78914 475634
rect 78294 439954 78914 475398
rect 78294 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 78914 439954
rect 78294 439634 78914 439718
rect 78294 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 78914 439634
rect 78294 403954 78914 439398
rect 78294 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 78914 403954
rect 78294 403634 78914 403718
rect 78294 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 78914 403634
rect 78294 367954 78914 403398
rect 78294 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 78914 367954
rect 78294 367634 78914 367718
rect 78294 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 78914 367634
rect 78294 331954 78914 367398
rect 78294 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 78914 331954
rect 78294 331634 78914 331718
rect 78294 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 78914 331634
rect 78294 295954 78914 331398
rect 78294 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 78914 295954
rect 78294 295634 78914 295718
rect 78294 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 78914 295634
rect 78294 259954 78914 295398
rect 78294 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 78914 259954
rect 78294 259634 78914 259718
rect 78294 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 78914 259634
rect 78294 244084 78914 259398
rect 82794 706758 83414 711590
rect 82794 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 83414 706758
rect 82794 706438 83414 706522
rect 82794 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 83414 706438
rect 82794 696454 83414 706202
rect 82794 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 83414 696454
rect 82794 696134 83414 696218
rect 82794 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 83414 696134
rect 82794 660454 83414 695898
rect 82794 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 83414 660454
rect 82794 660134 83414 660218
rect 82794 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 83414 660134
rect 82794 624454 83414 659898
rect 82794 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 83414 624454
rect 82794 624134 83414 624218
rect 82794 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 83414 624134
rect 82794 588454 83414 623898
rect 82794 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 83414 588454
rect 82794 588134 83414 588218
rect 82794 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 83414 588134
rect 82794 552454 83414 587898
rect 82794 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 83414 552454
rect 82794 552134 83414 552218
rect 82794 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 83414 552134
rect 82794 516454 83414 551898
rect 82794 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 83414 516454
rect 82794 516134 83414 516218
rect 82794 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 83414 516134
rect 82794 480454 83414 515898
rect 82794 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 83414 480454
rect 82794 480134 83414 480218
rect 82794 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 83414 480134
rect 82794 444454 83414 479898
rect 82794 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 83414 444454
rect 82794 444134 83414 444218
rect 82794 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 83414 444134
rect 82794 408454 83414 443898
rect 82794 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 83414 408454
rect 82794 408134 83414 408218
rect 82794 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 83414 408134
rect 82794 372454 83414 407898
rect 82794 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 83414 372454
rect 82794 372134 83414 372218
rect 82794 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 83414 372134
rect 82794 336454 83414 371898
rect 82794 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 83414 336454
rect 82794 336134 83414 336218
rect 82794 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 83414 336134
rect 82794 300454 83414 335898
rect 82794 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 83414 300454
rect 82794 300134 83414 300218
rect 82794 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 83414 300134
rect 82794 264454 83414 299898
rect 82794 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 83414 264454
rect 82794 264134 83414 264218
rect 82794 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 83414 264134
rect 82794 244084 83414 263898
rect 87294 707718 87914 711590
rect 87294 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 87914 707718
rect 87294 707398 87914 707482
rect 87294 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 87914 707398
rect 87294 700954 87914 707162
rect 87294 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 87914 700954
rect 87294 700634 87914 700718
rect 87294 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 87914 700634
rect 87294 664954 87914 700398
rect 87294 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 87914 664954
rect 87294 664634 87914 664718
rect 87294 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 87914 664634
rect 87294 628954 87914 664398
rect 87294 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 87914 628954
rect 87294 628634 87914 628718
rect 87294 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 87914 628634
rect 87294 592954 87914 628398
rect 87294 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 87914 592954
rect 87294 592634 87914 592718
rect 87294 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 87914 592634
rect 87294 556954 87914 592398
rect 87294 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 87914 556954
rect 87294 556634 87914 556718
rect 87294 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 87914 556634
rect 87294 520954 87914 556398
rect 87294 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 87914 520954
rect 87294 520634 87914 520718
rect 87294 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 87914 520634
rect 87294 484954 87914 520398
rect 87294 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 87914 484954
rect 87294 484634 87914 484718
rect 87294 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 87914 484634
rect 87294 448954 87914 484398
rect 87294 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 87914 448954
rect 87294 448634 87914 448718
rect 87294 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 87914 448634
rect 87294 412954 87914 448398
rect 87294 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 87914 412954
rect 87294 412634 87914 412718
rect 87294 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 87914 412634
rect 87294 376954 87914 412398
rect 87294 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 87914 376954
rect 87294 376634 87914 376718
rect 87294 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 87914 376634
rect 87294 340954 87914 376398
rect 87294 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 87914 340954
rect 87294 340634 87914 340718
rect 87294 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 87914 340634
rect 87294 304954 87914 340398
rect 87294 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 87914 304954
rect 87294 304634 87914 304718
rect 87294 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 87914 304634
rect 87294 268954 87914 304398
rect 87294 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 87914 268954
rect 87294 268634 87914 268718
rect 87294 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 87914 268634
rect 87294 244084 87914 268398
rect 91794 708678 92414 711590
rect 91794 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 92414 708678
rect 91794 708358 92414 708442
rect 91794 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 92414 708358
rect 91794 669454 92414 708122
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 273454 92414 308898
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 244084 92414 272898
rect 96294 709638 96914 711590
rect 96294 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 96914 709638
rect 96294 709318 96914 709402
rect 96294 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 96914 709318
rect 96294 673954 96914 709082
rect 96294 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 96914 673954
rect 96294 673634 96914 673718
rect 96294 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 96914 673634
rect 96294 637954 96914 673398
rect 96294 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 96914 637954
rect 96294 637634 96914 637718
rect 96294 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 96914 637634
rect 96294 601954 96914 637398
rect 96294 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 96914 601954
rect 96294 601634 96914 601718
rect 96294 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 96914 601634
rect 96294 565954 96914 601398
rect 96294 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 96914 565954
rect 96294 565634 96914 565718
rect 96294 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 96914 565634
rect 96294 529954 96914 565398
rect 96294 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 96914 529954
rect 96294 529634 96914 529718
rect 96294 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 96914 529634
rect 96294 493954 96914 529398
rect 96294 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 96914 493954
rect 96294 493634 96914 493718
rect 96294 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 96914 493634
rect 96294 457954 96914 493398
rect 96294 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 96914 457954
rect 96294 457634 96914 457718
rect 96294 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 96914 457634
rect 96294 421954 96914 457398
rect 96294 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 96914 421954
rect 96294 421634 96914 421718
rect 96294 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 96914 421634
rect 96294 385954 96914 421398
rect 96294 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 96914 385954
rect 96294 385634 96914 385718
rect 96294 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 96914 385634
rect 96294 349954 96914 385398
rect 96294 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 96914 349954
rect 96294 349634 96914 349718
rect 96294 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 96914 349634
rect 96294 313954 96914 349398
rect 96294 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 96914 313954
rect 96294 313634 96914 313718
rect 96294 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 96914 313634
rect 96294 277954 96914 313398
rect 96294 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 96914 277954
rect 96294 277634 96914 277718
rect 96294 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 96914 277634
rect 96294 244084 96914 277398
rect 100794 710598 101414 711590
rect 100794 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 101414 710598
rect 100794 710278 101414 710362
rect 100794 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 101414 710278
rect 100794 678454 101414 710042
rect 100794 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 101414 678454
rect 100794 678134 101414 678218
rect 100794 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 101414 678134
rect 100794 642454 101414 677898
rect 100794 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 101414 642454
rect 100794 642134 101414 642218
rect 100794 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 101414 642134
rect 100794 606454 101414 641898
rect 100794 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 101414 606454
rect 100794 606134 101414 606218
rect 100794 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 101414 606134
rect 100794 570454 101414 605898
rect 100794 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 101414 570454
rect 100794 570134 101414 570218
rect 100794 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 101414 570134
rect 100794 534454 101414 569898
rect 100794 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 101414 534454
rect 100794 534134 101414 534218
rect 100794 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 101414 534134
rect 100794 498454 101414 533898
rect 100794 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 101414 498454
rect 100794 498134 101414 498218
rect 100794 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 101414 498134
rect 100794 462454 101414 497898
rect 100794 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 101414 462454
rect 100794 462134 101414 462218
rect 100794 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 101414 462134
rect 100794 426454 101414 461898
rect 100794 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 101414 426454
rect 100794 426134 101414 426218
rect 100794 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 101414 426134
rect 100794 390454 101414 425898
rect 100794 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 101414 390454
rect 100794 390134 101414 390218
rect 100794 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 101414 390134
rect 100794 354454 101414 389898
rect 100794 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 101414 354454
rect 100794 354134 101414 354218
rect 100794 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 101414 354134
rect 100794 318454 101414 353898
rect 100794 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 101414 318454
rect 100794 318134 101414 318218
rect 100794 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 101414 318134
rect 100794 282454 101414 317898
rect 100794 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 101414 282454
rect 100794 282134 101414 282218
rect 100794 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 101414 282134
rect 100794 246454 101414 281898
rect 100794 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 101414 246454
rect 100794 246134 101414 246218
rect 100794 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 101414 246134
rect 100794 244084 101414 245898
rect 105294 711558 105914 711590
rect 105294 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 105914 711558
rect 105294 711238 105914 711322
rect 105294 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 105914 711238
rect 105294 682954 105914 711002
rect 105294 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 105914 682954
rect 105294 682634 105914 682718
rect 105294 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 105914 682634
rect 105294 646954 105914 682398
rect 105294 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 105914 646954
rect 105294 646634 105914 646718
rect 105294 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 105914 646634
rect 105294 610954 105914 646398
rect 105294 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 105914 610954
rect 105294 610634 105914 610718
rect 105294 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 105914 610634
rect 105294 574954 105914 610398
rect 105294 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 105914 574954
rect 105294 574634 105914 574718
rect 105294 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 105914 574634
rect 105294 538954 105914 574398
rect 105294 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 105914 538954
rect 105294 538634 105914 538718
rect 105294 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 105914 538634
rect 105294 502954 105914 538398
rect 105294 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 105914 502954
rect 105294 502634 105914 502718
rect 105294 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 105914 502634
rect 105294 466954 105914 502398
rect 105294 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 105914 466954
rect 105294 466634 105914 466718
rect 105294 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 105914 466634
rect 105294 430954 105914 466398
rect 105294 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 105914 430954
rect 105294 430634 105914 430718
rect 105294 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 105914 430634
rect 105294 394954 105914 430398
rect 105294 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 105914 394954
rect 105294 394634 105914 394718
rect 105294 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 105914 394634
rect 105294 358954 105914 394398
rect 105294 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 105914 358954
rect 105294 358634 105914 358718
rect 105294 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 105914 358634
rect 105294 322954 105914 358398
rect 105294 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 105914 322954
rect 105294 322634 105914 322718
rect 105294 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 105914 322634
rect 105294 286954 105914 322398
rect 105294 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 105914 286954
rect 105294 286634 105914 286718
rect 105294 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 105914 286634
rect 105294 250954 105914 286398
rect 105294 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 105914 250954
rect 105294 250634 105914 250718
rect 105294 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 105914 250634
rect 105294 244084 105914 250398
rect 109794 704838 110414 711590
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 244084 110414 254898
rect 114294 705798 114914 711590
rect 114294 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 114914 705798
rect 114294 705478 114914 705562
rect 114294 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 114914 705478
rect 114294 691954 114914 705242
rect 114294 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 114914 691954
rect 114294 691634 114914 691718
rect 114294 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 114914 691634
rect 114294 655954 114914 691398
rect 114294 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 114914 655954
rect 114294 655634 114914 655718
rect 114294 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 114914 655634
rect 114294 619954 114914 655398
rect 114294 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 114914 619954
rect 114294 619634 114914 619718
rect 114294 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 114914 619634
rect 114294 583954 114914 619398
rect 114294 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 114914 583954
rect 114294 583634 114914 583718
rect 114294 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 114914 583634
rect 114294 547954 114914 583398
rect 114294 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 114914 547954
rect 114294 547634 114914 547718
rect 114294 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 114914 547634
rect 114294 511954 114914 547398
rect 114294 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 114914 511954
rect 114294 511634 114914 511718
rect 114294 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 114914 511634
rect 114294 475954 114914 511398
rect 114294 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 114914 475954
rect 114294 475634 114914 475718
rect 114294 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 114914 475634
rect 114294 439954 114914 475398
rect 114294 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 114914 439954
rect 114294 439634 114914 439718
rect 114294 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 114914 439634
rect 114294 403954 114914 439398
rect 114294 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 114914 403954
rect 114294 403634 114914 403718
rect 114294 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 114914 403634
rect 114294 367954 114914 403398
rect 114294 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 114914 367954
rect 114294 367634 114914 367718
rect 114294 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 114914 367634
rect 114294 331954 114914 367398
rect 114294 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 114914 331954
rect 114294 331634 114914 331718
rect 114294 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 114914 331634
rect 114294 295954 114914 331398
rect 114294 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 114914 295954
rect 114294 295634 114914 295718
rect 114294 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 114914 295634
rect 114294 259954 114914 295398
rect 114294 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 114914 259954
rect 114294 259634 114914 259718
rect 114294 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 114914 259634
rect 114294 244084 114914 259398
rect 118794 706758 119414 711590
rect 118794 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 119414 706758
rect 118794 706438 119414 706522
rect 118794 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 119414 706438
rect 118794 696454 119414 706202
rect 118794 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 119414 696454
rect 118794 696134 119414 696218
rect 118794 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 119414 696134
rect 118794 660454 119414 695898
rect 118794 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 119414 660454
rect 118794 660134 119414 660218
rect 118794 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 119414 660134
rect 118794 624454 119414 659898
rect 118794 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 119414 624454
rect 118794 624134 119414 624218
rect 118794 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 119414 624134
rect 118794 588454 119414 623898
rect 118794 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 119414 588454
rect 118794 588134 119414 588218
rect 118794 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 119414 588134
rect 118794 552454 119414 587898
rect 118794 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 119414 552454
rect 118794 552134 119414 552218
rect 118794 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 119414 552134
rect 118794 516454 119414 551898
rect 118794 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 119414 516454
rect 118794 516134 119414 516218
rect 118794 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 119414 516134
rect 118794 480454 119414 515898
rect 118794 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 119414 480454
rect 118794 480134 119414 480218
rect 118794 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 119414 480134
rect 118794 444454 119414 479898
rect 118794 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 119414 444454
rect 118794 444134 119414 444218
rect 118794 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 119414 444134
rect 118794 408454 119414 443898
rect 118794 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 119414 408454
rect 118794 408134 119414 408218
rect 118794 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 119414 408134
rect 118794 372454 119414 407898
rect 118794 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 119414 372454
rect 118794 372134 119414 372218
rect 118794 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 119414 372134
rect 118794 336454 119414 371898
rect 118794 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 119414 336454
rect 118794 336134 119414 336218
rect 118794 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 119414 336134
rect 118794 300454 119414 335898
rect 118794 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 119414 300454
rect 118794 300134 119414 300218
rect 118794 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 119414 300134
rect 118794 264454 119414 299898
rect 118794 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 119414 264454
rect 118794 264134 119414 264218
rect 118794 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 119414 264134
rect 118794 244084 119414 263898
rect 123294 707718 123914 711590
rect 123294 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 123914 707718
rect 123294 707398 123914 707482
rect 123294 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 123914 707398
rect 123294 700954 123914 707162
rect 123294 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 123914 700954
rect 123294 700634 123914 700718
rect 123294 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 123914 700634
rect 123294 664954 123914 700398
rect 123294 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 123914 664954
rect 123294 664634 123914 664718
rect 123294 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 123914 664634
rect 123294 628954 123914 664398
rect 123294 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 123914 628954
rect 123294 628634 123914 628718
rect 123294 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 123914 628634
rect 123294 592954 123914 628398
rect 123294 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 123914 592954
rect 123294 592634 123914 592718
rect 123294 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 123914 592634
rect 123294 556954 123914 592398
rect 123294 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 123914 556954
rect 123294 556634 123914 556718
rect 123294 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 123914 556634
rect 123294 520954 123914 556398
rect 123294 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 123914 520954
rect 123294 520634 123914 520718
rect 123294 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 123914 520634
rect 123294 484954 123914 520398
rect 123294 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 123914 484954
rect 123294 484634 123914 484718
rect 123294 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 123914 484634
rect 123294 448954 123914 484398
rect 123294 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 123914 448954
rect 123294 448634 123914 448718
rect 123294 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 123914 448634
rect 123294 412954 123914 448398
rect 123294 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 123914 412954
rect 123294 412634 123914 412718
rect 123294 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 123914 412634
rect 123294 376954 123914 412398
rect 123294 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 123914 376954
rect 123294 376634 123914 376718
rect 123294 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 123914 376634
rect 123294 340954 123914 376398
rect 123294 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 123914 340954
rect 123294 340634 123914 340718
rect 123294 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 123914 340634
rect 123294 304954 123914 340398
rect 123294 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 123914 304954
rect 123294 304634 123914 304718
rect 123294 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 123914 304634
rect 123294 268954 123914 304398
rect 123294 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 123914 268954
rect 123294 268634 123914 268718
rect 123294 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 123914 268634
rect 123294 244084 123914 268398
rect 127794 708678 128414 711590
rect 127794 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 128414 708678
rect 127794 708358 128414 708442
rect 127794 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 128414 708358
rect 127794 669454 128414 708122
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 244084 128414 272898
rect 132294 709638 132914 711590
rect 132294 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 132914 709638
rect 132294 709318 132914 709402
rect 132294 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 132914 709318
rect 132294 673954 132914 709082
rect 132294 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 132914 673954
rect 132294 673634 132914 673718
rect 132294 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 132914 673634
rect 132294 637954 132914 673398
rect 132294 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 132914 637954
rect 132294 637634 132914 637718
rect 132294 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 132914 637634
rect 132294 601954 132914 637398
rect 132294 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 132914 601954
rect 132294 601634 132914 601718
rect 132294 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 132914 601634
rect 132294 565954 132914 601398
rect 132294 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 132914 565954
rect 132294 565634 132914 565718
rect 132294 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 132914 565634
rect 132294 529954 132914 565398
rect 132294 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 132914 529954
rect 132294 529634 132914 529718
rect 132294 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 132914 529634
rect 132294 493954 132914 529398
rect 132294 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 132914 493954
rect 132294 493634 132914 493718
rect 132294 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 132914 493634
rect 132294 457954 132914 493398
rect 132294 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 132914 457954
rect 132294 457634 132914 457718
rect 132294 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 132914 457634
rect 132294 421954 132914 457398
rect 132294 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 132914 421954
rect 132294 421634 132914 421718
rect 132294 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 132914 421634
rect 132294 385954 132914 421398
rect 132294 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 132914 385954
rect 132294 385634 132914 385718
rect 132294 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 132914 385634
rect 132294 349954 132914 385398
rect 132294 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 132914 349954
rect 132294 349634 132914 349718
rect 132294 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 132914 349634
rect 132294 313954 132914 349398
rect 132294 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 132914 313954
rect 132294 313634 132914 313718
rect 132294 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 132914 313634
rect 132294 277954 132914 313398
rect 132294 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 132914 277954
rect 132294 277634 132914 277718
rect 132294 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 132914 277634
rect 132294 244084 132914 277398
rect 136794 710598 137414 711590
rect 136794 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 137414 710598
rect 136794 710278 137414 710362
rect 136794 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 137414 710278
rect 136794 678454 137414 710042
rect 136794 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 137414 678454
rect 136794 678134 137414 678218
rect 136794 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 137414 678134
rect 136794 642454 137414 677898
rect 136794 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 137414 642454
rect 136794 642134 137414 642218
rect 136794 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 137414 642134
rect 136794 606454 137414 641898
rect 136794 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 137414 606454
rect 136794 606134 137414 606218
rect 136794 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 137414 606134
rect 136794 570454 137414 605898
rect 136794 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 137414 570454
rect 136794 570134 137414 570218
rect 136794 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 137414 570134
rect 136794 534454 137414 569898
rect 136794 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 137414 534454
rect 136794 534134 137414 534218
rect 136794 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 137414 534134
rect 136794 498454 137414 533898
rect 136794 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 137414 498454
rect 136794 498134 137414 498218
rect 136794 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 137414 498134
rect 136794 462454 137414 497898
rect 136794 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 137414 462454
rect 136794 462134 137414 462218
rect 136794 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 137414 462134
rect 136794 426454 137414 461898
rect 136794 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 137414 426454
rect 136794 426134 137414 426218
rect 136794 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 137414 426134
rect 136794 390454 137414 425898
rect 136794 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 137414 390454
rect 136794 390134 137414 390218
rect 136794 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 137414 390134
rect 136794 354454 137414 389898
rect 136794 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 137414 354454
rect 136794 354134 137414 354218
rect 136794 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 137414 354134
rect 136794 318454 137414 353898
rect 136794 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 137414 318454
rect 136794 318134 137414 318218
rect 136794 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 137414 318134
rect 136794 282454 137414 317898
rect 136794 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 137414 282454
rect 136794 282134 137414 282218
rect 136794 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 137414 282134
rect 136794 246454 137414 281898
rect 136794 246218 136826 246454
rect 137062 246218 137146 246454
rect 137382 246218 137414 246454
rect 136794 246134 137414 246218
rect 136794 245898 136826 246134
rect 137062 245898 137146 246134
rect 137382 245898 137414 246134
rect 136794 244084 137414 245898
rect 141294 711558 141914 711590
rect 141294 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 141914 711558
rect 141294 711238 141914 711322
rect 141294 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 141914 711238
rect 141294 682954 141914 711002
rect 141294 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 141914 682954
rect 141294 682634 141914 682718
rect 141294 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 141914 682634
rect 141294 646954 141914 682398
rect 141294 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 141914 646954
rect 141294 646634 141914 646718
rect 141294 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 141914 646634
rect 141294 610954 141914 646398
rect 141294 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 141914 610954
rect 141294 610634 141914 610718
rect 141294 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 141914 610634
rect 141294 574954 141914 610398
rect 141294 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 141914 574954
rect 141294 574634 141914 574718
rect 141294 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 141914 574634
rect 141294 538954 141914 574398
rect 141294 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 141914 538954
rect 141294 538634 141914 538718
rect 141294 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 141914 538634
rect 141294 502954 141914 538398
rect 141294 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 141914 502954
rect 141294 502634 141914 502718
rect 141294 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 141914 502634
rect 141294 466954 141914 502398
rect 141294 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 141914 466954
rect 141294 466634 141914 466718
rect 141294 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 141914 466634
rect 141294 430954 141914 466398
rect 141294 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 141914 430954
rect 141294 430634 141914 430718
rect 141294 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 141914 430634
rect 141294 394954 141914 430398
rect 141294 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 141914 394954
rect 141294 394634 141914 394718
rect 141294 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 141914 394634
rect 141294 358954 141914 394398
rect 141294 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 141914 358954
rect 141294 358634 141914 358718
rect 141294 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 141914 358634
rect 141294 322954 141914 358398
rect 141294 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 141914 322954
rect 141294 322634 141914 322718
rect 141294 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 141914 322634
rect 141294 286954 141914 322398
rect 141294 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 141914 286954
rect 141294 286634 141914 286718
rect 141294 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 141914 286634
rect 141294 250954 141914 286398
rect 141294 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 141914 250954
rect 141294 250634 141914 250718
rect 141294 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 141914 250634
rect 141294 244084 141914 250398
rect 145794 704838 146414 711590
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 244084 146414 254898
rect 150294 705798 150914 711590
rect 150294 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 150914 705798
rect 150294 705478 150914 705562
rect 150294 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 150914 705478
rect 150294 691954 150914 705242
rect 150294 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 150914 691954
rect 150294 691634 150914 691718
rect 150294 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 150914 691634
rect 150294 655954 150914 691398
rect 150294 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 150914 655954
rect 150294 655634 150914 655718
rect 150294 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 150914 655634
rect 150294 619954 150914 655398
rect 150294 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 150914 619954
rect 150294 619634 150914 619718
rect 150294 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 150914 619634
rect 150294 583954 150914 619398
rect 150294 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 150914 583954
rect 150294 583634 150914 583718
rect 150294 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 150914 583634
rect 150294 547954 150914 583398
rect 150294 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 150914 547954
rect 150294 547634 150914 547718
rect 150294 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 150914 547634
rect 150294 511954 150914 547398
rect 150294 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 150914 511954
rect 150294 511634 150914 511718
rect 150294 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 150914 511634
rect 150294 475954 150914 511398
rect 150294 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 150914 475954
rect 150294 475634 150914 475718
rect 150294 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 150914 475634
rect 150294 439954 150914 475398
rect 150294 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 150914 439954
rect 150294 439634 150914 439718
rect 150294 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 150914 439634
rect 150294 403954 150914 439398
rect 150294 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 150914 403954
rect 150294 403634 150914 403718
rect 150294 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 150914 403634
rect 150294 367954 150914 403398
rect 150294 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 150914 367954
rect 150294 367634 150914 367718
rect 150294 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 150914 367634
rect 150294 331954 150914 367398
rect 150294 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 150914 331954
rect 150294 331634 150914 331718
rect 150294 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 150914 331634
rect 150294 295954 150914 331398
rect 150294 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 150914 295954
rect 150294 295634 150914 295718
rect 150294 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 150914 295634
rect 150294 259954 150914 295398
rect 150294 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 150914 259954
rect 150294 259634 150914 259718
rect 150294 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 150914 259634
rect 150294 244084 150914 259398
rect 154794 706758 155414 711590
rect 154794 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 155414 706758
rect 154794 706438 155414 706522
rect 154794 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 155414 706438
rect 154794 696454 155414 706202
rect 154794 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 155414 696454
rect 154794 696134 155414 696218
rect 154794 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 155414 696134
rect 154794 660454 155414 695898
rect 154794 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 155414 660454
rect 154794 660134 155414 660218
rect 154794 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 155414 660134
rect 154794 624454 155414 659898
rect 154794 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 155414 624454
rect 154794 624134 155414 624218
rect 154794 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 155414 624134
rect 154794 588454 155414 623898
rect 154794 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 155414 588454
rect 154794 588134 155414 588218
rect 154794 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 155414 588134
rect 154794 552454 155414 587898
rect 154794 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 155414 552454
rect 154794 552134 155414 552218
rect 154794 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 155414 552134
rect 154794 516454 155414 551898
rect 154794 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 155414 516454
rect 154794 516134 155414 516218
rect 154794 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 155414 516134
rect 154794 480454 155414 515898
rect 154794 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 155414 480454
rect 154794 480134 155414 480218
rect 154794 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 155414 480134
rect 154794 444454 155414 479898
rect 154794 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 155414 444454
rect 154794 444134 155414 444218
rect 154794 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 155414 444134
rect 154794 408454 155414 443898
rect 154794 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 155414 408454
rect 154794 408134 155414 408218
rect 154794 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 155414 408134
rect 154794 372454 155414 407898
rect 154794 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 155414 372454
rect 154794 372134 155414 372218
rect 154794 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 155414 372134
rect 154794 336454 155414 371898
rect 154794 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 155414 336454
rect 154794 336134 155414 336218
rect 154794 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 155414 336134
rect 154794 300454 155414 335898
rect 154794 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 155414 300454
rect 154794 300134 155414 300218
rect 154794 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 155414 300134
rect 154794 264454 155414 299898
rect 154794 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 155414 264454
rect 154794 264134 155414 264218
rect 154794 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 155414 264134
rect 154794 244084 155414 263898
rect 159294 707718 159914 711590
rect 159294 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 159914 707718
rect 159294 707398 159914 707482
rect 159294 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 159914 707398
rect 159294 700954 159914 707162
rect 159294 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 159914 700954
rect 159294 700634 159914 700718
rect 159294 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 159914 700634
rect 159294 664954 159914 700398
rect 159294 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 159914 664954
rect 159294 664634 159914 664718
rect 159294 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 159914 664634
rect 159294 628954 159914 664398
rect 159294 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 159914 628954
rect 159294 628634 159914 628718
rect 159294 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 159914 628634
rect 159294 592954 159914 628398
rect 159294 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 159914 592954
rect 159294 592634 159914 592718
rect 159294 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 159914 592634
rect 159294 556954 159914 592398
rect 159294 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 159914 556954
rect 159294 556634 159914 556718
rect 159294 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 159914 556634
rect 159294 520954 159914 556398
rect 159294 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 159914 520954
rect 159294 520634 159914 520718
rect 159294 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 159914 520634
rect 159294 484954 159914 520398
rect 159294 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 159914 484954
rect 159294 484634 159914 484718
rect 159294 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 159914 484634
rect 159294 448954 159914 484398
rect 159294 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 159914 448954
rect 159294 448634 159914 448718
rect 159294 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 159914 448634
rect 159294 412954 159914 448398
rect 159294 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 159914 412954
rect 159294 412634 159914 412718
rect 159294 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 159914 412634
rect 159294 376954 159914 412398
rect 159294 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 159914 376954
rect 159294 376634 159914 376718
rect 159294 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 159914 376634
rect 159294 340954 159914 376398
rect 159294 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 159914 340954
rect 159294 340634 159914 340718
rect 159294 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 159914 340634
rect 159294 304954 159914 340398
rect 159294 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 159914 304954
rect 159294 304634 159914 304718
rect 159294 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 159914 304634
rect 159294 268954 159914 304398
rect 159294 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 159914 268954
rect 159294 268634 159914 268718
rect 159294 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 159914 268634
rect 159294 244084 159914 268398
rect 163794 708678 164414 711590
rect 163794 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 164414 708678
rect 163794 708358 164414 708442
rect 163794 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 164414 708358
rect 163794 669454 164414 708122
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 244084 164414 272898
rect 168294 709638 168914 711590
rect 168294 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 168914 709638
rect 168294 709318 168914 709402
rect 168294 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 168914 709318
rect 168294 673954 168914 709082
rect 168294 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 168914 673954
rect 168294 673634 168914 673718
rect 168294 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 168914 673634
rect 168294 637954 168914 673398
rect 168294 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 168914 637954
rect 168294 637634 168914 637718
rect 168294 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 168914 637634
rect 168294 601954 168914 637398
rect 168294 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 168914 601954
rect 168294 601634 168914 601718
rect 168294 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 168914 601634
rect 168294 565954 168914 601398
rect 168294 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 168914 565954
rect 168294 565634 168914 565718
rect 168294 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 168914 565634
rect 168294 529954 168914 565398
rect 168294 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 168914 529954
rect 168294 529634 168914 529718
rect 168294 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 168914 529634
rect 168294 493954 168914 529398
rect 168294 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 168914 493954
rect 168294 493634 168914 493718
rect 168294 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 168914 493634
rect 168294 457954 168914 493398
rect 168294 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 168914 457954
rect 168294 457634 168914 457718
rect 168294 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 168914 457634
rect 168294 421954 168914 457398
rect 168294 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 168914 421954
rect 168294 421634 168914 421718
rect 168294 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 168914 421634
rect 168294 385954 168914 421398
rect 168294 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 168914 385954
rect 168294 385634 168914 385718
rect 168294 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 168914 385634
rect 168294 349954 168914 385398
rect 168294 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 168914 349954
rect 168294 349634 168914 349718
rect 168294 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 168914 349634
rect 168294 313954 168914 349398
rect 168294 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 168914 313954
rect 168294 313634 168914 313718
rect 168294 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 168914 313634
rect 168294 277954 168914 313398
rect 168294 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 168914 277954
rect 168294 277634 168914 277718
rect 168294 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 168914 277634
rect 168294 244084 168914 277398
rect 172794 710598 173414 711590
rect 172794 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 173414 710598
rect 172794 710278 173414 710362
rect 172794 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 173414 710278
rect 172794 678454 173414 710042
rect 172794 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 173414 678454
rect 172794 678134 173414 678218
rect 172794 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 173414 678134
rect 172794 642454 173414 677898
rect 172794 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 173414 642454
rect 172794 642134 173414 642218
rect 172794 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 173414 642134
rect 172794 606454 173414 641898
rect 172794 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 173414 606454
rect 172794 606134 173414 606218
rect 172794 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 173414 606134
rect 172794 570454 173414 605898
rect 172794 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 173414 570454
rect 172794 570134 173414 570218
rect 172794 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 173414 570134
rect 172794 534454 173414 569898
rect 172794 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 173414 534454
rect 172794 534134 173414 534218
rect 172794 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 173414 534134
rect 172794 498454 173414 533898
rect 172794 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 173414 498454
rect 172794 498134 173414 498218
rect 172794 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 173414 498134
rect 172794 462454 173414 497898
rect 172794 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 173414 462454
rect 172794 462134 173414 462218
rect 172794 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 173414 462134
rect 172794 426454 173414 461898
rect 172794 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 173414 426454
rect 172794 426134 173414 426218
rect 172794 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 173414 426134
rect 172794 390454 173414 425898
rect 172794 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 173414 390454
rect 172794 390134 173414 390218
rect 172794 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 173414 390134
rect 172794 354454 173414 389898
rect 172794 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 173414 354454
rect 172794 354134 173414 354218
rect 172794 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 173414 354134
rect 172794 318454 173414 353898
rect 172794 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 173414 318454
rect 172794 318134 173414 318218
rect 172794 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 173414 318134
rect 172794 282454 173414 317898
rect 172794 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 173414 282454
rect 172794 282134 173414 282218
rect 172794 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 173414 282134
rect 172794 246454 173414 281898
rect 172794 246218 172826 246454
rect 173062 246218 173146 246454
rect 173382 246218 173414 246454
rect 172794 246134 173414 246218
rect 172794 245898 172826 246134
rect 173062 245898 173146 246134
rect 173382 245898 173414 246134
rect 172794 244084 173414 245898
rect 177294 711558 177914 711590
rect 177294 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 177914 711558
rect 177294 711238 177914 711322
rect 177294 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 177914 711238
rect 177294 682954 177914 711002
rect 177294 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 177914 682954
rect 177294 682634 177914 682718
rect 177294 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 177914 682634
rect 177294 646954 177914 682398
rect 177294 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 177914 646954
rect 177294 646634 177914 646718
rect 177294 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 177914 646634
rect 177294 610954 177914 646398
rect 177294 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 177914 610954
rect 177294 610634 177914 610718
rect 177294 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 177914 610634
rect 177294 574954 177914 610398
rect 177294 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 177914 574954
rect 177294 574634 177914 574718
rect 177294 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 177914 574634
rect 177294 538954 177914 574398
rect 177294 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 177914 538954
rect 177294 538634 177914 538718
rect 177294 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 177914 538634
rect 177294 502954 177914 538398
rect 177294 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 177914 502954
rect 177294 502634 177914 502718
rect 177294 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 177914 502634
rect 177294 466954 177914 502398
rect 177294 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 177914 466954
rect 177294 466634 177914 466718
rect 177294 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 177914 466634
rect 177294 430954 177914 466398
rect 177294 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 177914 430954
rect 177294 430634 177914 430718
rect 177294 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 177914 430634
rect 177294 394954 177914 430398
rect 177294 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 177914 394954
rect 177294 394634 177914 394718
rect 177294 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 177914 394634
rect 177294 358954 177914 394398
rect 177294 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 177914 358954
rect 177294 358634 177914 358718
rect 177294 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 177914 358634
rect 177294 322954 177914 358398
rect 177294 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 177914 322954
rect 177294 322634 177914 322718
rect 177294 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 177914 322634
rect 177294 286954 177914 322398
rect 177294 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 177914 286954
rect 177294 286634 177914 286718
rect 177294 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 177914 286634
rect 177294 250954 177914 286398
rect 177294 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 177914 250954
rect 177294 250634 177914 250718
rect 177294 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 177914 250634
rect 177294 244084 177914 250398
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 244084 182414 254898
rect 186294 705798 186914 711590
rect 186294 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 186914 705798
rect 186294 705478 186914 705562
rect 186294 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 186914 705478
rect 186294 691954 186914 705242
rect 186294 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 186914 691954
rect 186294 691634 186914 691718
rect 186294 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 186914 691634
rect 186294 655954 186914 691398
rect 186294 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 186914 655954
rect 186294 655634 186914 655718
rect 186294 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 186914 655634
rect 186294 619954 186914 655398
rect 186294 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 186914 619954
rect 186294 619634 186914 619718
rect 186294 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 186914 619634
rect 186294 583954 186914 619398
rect 186294 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 186914 583954
rect 186294 583634 186914 583718
rect 186294 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 186914 583634
rect 186294 547954 186914 583398
rect 186294 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 186914 547954
rect 186294 547634 186914 547718
rect 186294 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 186914 547634
rect 186294 511954 186914 547398
rect 186294 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 186914 511954
rect 186294 511634 186914 511718
rect 186294 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 186914 511634
rect 186294 475954 186914 511398
rect 186294 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 186914 475954
rect 186294 475634 186914 475718
rect 186294 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 186914 475634
rect 186294 439954 186914 475398
rect 186294 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 186914 439954
rect 186294 439634 186914 439718
rect 186294 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 186914 439634
rect 186294 403954 186914 439398
rect 186294 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 186914 403954
rect 186294 403634 186914 403718
rect 186294 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 186914 403634
rect 186294 367954 186914 403398
rect 186294 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 186914 367954
rect 186294 367634 186914 367718
rect 186294 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 186914 367634
rect 186294 331954 186914 367398
rect 186294 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 186914 331954
rect 186294 331634 186914 331718
rect 186294 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 186914 331634
rect 186294 295954 186914 331398
rect 186294 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 186914 295954
rect 186294 295634 186914 295718
rect 186294 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 186914 295634
rect 186294 259954 186914 295398
rect 186294 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 186914 259954
rect 186294 259634 186914 259718
rect 186294 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 186914 259634
rect 186294 244084 186914 259398
rect 190794 706758 191414 711590
rect 190794 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 191414 706758
rect 190794 706438 191414 706522
rect 190794 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 191414 706438
rect 190794 696454 191414 706202
rect 190794 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 191414 696454
rect 190794 696134 191414 696218
rect 190794 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 191414 696134
rect 190794 660454 191414 695898
rect 190794 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 191414 660454
rect 190794 660134 191414 660218
rect 190794 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 191414 660134
rect 190794 624454 191414 659898
rect 190794 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 191414 624454
rect 190794 624134 191414 624218
rect 190794 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 191414 624134
rect 190794 588454 191414 623898
rect 190794 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 191414 588454
rect 190794 588134 191414 588218
rect 190794 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 191414 588134
rect 190794 552454 191414 587898
rect 190794 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 191414 552454
rect 190794 552134 191414 552218
rect 190794 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 191414 552134
rect 190794 516454 191414 551898
rect 190794 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 191414 516454
rect 190794 516134 191414 516218
rect 190794 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 191414 516134
rect 190794 480454 191414 515898
rect 190794 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 191414 480454
rect 190794 480134 191414 480218
rect 190794 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 191414 480134
rect 190794 444454 191414 479898
rect 190794 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 191414 444454
rect 190794 444134 191414 444218
rect 190794 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 191414 444134
rect 190794 408454 191414 443898
rect 190794 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 191414 408454
rect 190794 408134 191414 408218
rect 190794 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 191414 408134
rect 190794 372454 191414 407898
rect 190794 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 191414 372454
rect 190794 372134 191414 372218
rect 190794 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 191414 372134
rect 190794 336454 191414 371898
rect 190794 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 191414 336454
rect 190794 336134 191414 336218
rect 190794 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 191414 336134
rect 190794 300454 191414 335898
rect 190794 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 191414 300454
rect 190794 300134 191414 300218
rect 190794 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 191414 300134
rect 190794 264454 191414 299898
rect 190794 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 191414 264454
rect 190794 264134 191414 264218
rect 190794 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 191414 264134
rect 190794 244084 191414 263898
rect 195294 707718 195914 711590
rect 195294 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 195914 707718
rect 195294 707398 195914 707482
rect 195294 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 195914 707398
rect 195294 700954 195914 707162
rect 195294 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 195914 700954
rect 195294 700634 195914 700718
rect 195294 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 195914 700634
rect 195294 664954 195914 700398
rect 195294 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 195914 664954
rect 195294 664634 195914 664718
rect 195294 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 195914 664634
rect 195294 628954 195914 664398
rect 195294 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 195914 628954
rect 195294 628634 195914 628718
rect 195294 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 195914 628634
rect 195294 592954 195914 628398
rect 195294 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 195914 592954
rect 195294 592634 195914 592718
rect 195294 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 195914 592634
rect 195294 556954 195914 592398
rect 195294 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 195914 556954
rect 195294 556634 195914 556718
rect 195294 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 195914 556634
rect 195294 520954 195914 556398
rect 195294 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 195914 520954
rect 195294 520634 195914 520718
rect 195294 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 195914 520634
rect 195294 484954 195914 520398
rect 195294 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 195914 484954
rect 195294 484634 195914 484718
rect 195294 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 195914 484634
rect 195294 448954 195914 484398
rect 195294 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 195914 448954
rect 195294 448634 195914 448718
rect 195294 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 195914 448634
rect 195294 412954 195914 448398
rect 195294 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 195914 412954
rect 195294 412634 195914 412718
rect 195294 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 195914 412634
rect 195294 376954 195914 412398
rect 195294 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 195914 376954
rect 195294 376634 195914 376718
rect 195294 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 195914 376634
rect 195294 340954 195914 376398
rect 195294 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 195914 340954
rect 195294 340634 195914 340718
rect 195294 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 195914 340634
rect 195294 304954 195914 340398
rect 195294 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 195914 304954
rect 195294 304634 195914 304718
rect 195294 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 195914 304634
rect 195294 268954 195914 304398
rect 195294 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 195914 268954
rect 195294 268634 195914 268718
rect 195294 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 195914 268634
rect 195294 244084 195914 268398
rect 199794 708678 200414 711590
rect 199794 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 200414 708678
rect 199794 708358 200414 708442
rect 199794 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 200414 708358
rect 199794 669454 200414 708122
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199794 244084 200414 272898
rect 204294 709638 204914 711590
rect 204294 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 204914 709638
rect 204294 709318 204914 709402
rect 204294 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 204914 709318
rect 204294 673954 204914 709082
rect 204294 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 204914 673954
rect 204294 673634 204914 673718
rect 204294 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 204914 673634
rect 204294 637954 204914 673398
rect 204294 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 204914 637954
rect 204294 637634 204914 637718
rect 204294 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 204914 637634
rect 204294 601954 204914 637398
rect 204294 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 204914 601954
rect 204294 601634 204914 601718
rect 204294 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 204914 601634
rect 204294 565954 204914 601398
rect 204294 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 204914 565954
rect 204294 565634 204914 565718
rect 204294 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 204914 565634
rect 204294 529954 204914 565398
rect 204294 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 204914 529954
rect 204294 529634 204914 529718
rect 204294 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 204914 529634
rect 204294 493954 204914 529398
rect 204294 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 204914 493954
rect 204294 493634 204914 493718
rect 204294 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 204914 493634
rect 204294 457954 204914 493398
rect 204294 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 204914 457954
rect 204294 457634 204914 457718
rect 204294 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 204914 457634
rect 204294 421954 204914 457398
rect 204294 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 204914 421954
rect 204294 421634 204914 421718
rect 204294 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 204914 421634
rect 204294 385954 204914 421398
rect 204294 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 204914 385954
rect 204294 385634 204914 385718
rect 204294 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 204914 385634
rect 204294 349954 204914 385398
rect 204294 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 204914 349954
rect 204294 349634 204914 349718
rect 204294 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 204914 349634
rect 204294 313954 204914 349398
rect 204294 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 204914 313954
rect 204294 313634 204914 313718
rect 204294 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 204914 313634
rect 204294 277954 204914 313398
rect 204294 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 204914 277954
rect 204294 277634 204914 277718
rect 204294 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 204914 277634
rect 204294 244084 204914 277398
rect 208794 710598 209414 711590
rect 208794 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 209414 710598
rect 208794 710278 209414 710362
rect 208794 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 209414 710278
rect 208794 678454 209414 710042
rect 208794 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 209414 678454
rect 208794 678134 209414 678218
rect 208794 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 209414 678134
rect 208794 642454 209414 677898
rect 208794 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 209414 642454
rect 208794 642134 209414 642218
rect 208794 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 209414 642134
rect 208794 606454 209414 641898
rect 208794 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 209414 606454
rect 208794 606134 209414 606218
rect 208794 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 209414 606134
rect 208794 570454 209414 605898
rect 208794 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 209414 570454
rect 208794 570134 209414 570218
rect 208794 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 209414 570134
rect 208794 534454 209414 569898
rect 208794 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 209414 534454
rect 208794 534134 209414 534218
rect 208794 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 209414 534134
rect 208794 498454 209414 533898
rect 208794 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 209414 498454
rect 208794 498134 209414 498218
rect 208794 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 209414 498134
rect 208794 462454 209414 497898
rect 208794 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 209414 462454
rect 208794 462134 209414 462218
rect 208794 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 209414 462134
rect 208794 426454 209414 461898
rect 208794 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 209414 426454
rect 208794 426134 209414 426218
rect 208794 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 209414 426134
rect 208794 390454 209414 425898
rect 208794 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 209414 390454
rect 208794 390134 209414 390218
rect 208794 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 209414 390134
rect 208794 354454 209414 389898
rect 208794 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 209414 354454
rect 208794 354134 209414 354218
rect 208794 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 209414 354134
rect 208794 318454 209414 353898
rect 208794 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 209414 318454
rect 208794 318134 209414 318218
rect 208794 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 209414 318134
rect 208794 282454 209414 317898
rect 208794 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 209414 282454
rect 208794 282134 209414 282218
rect 208794 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 209414 282134
rect 208794 246454 209414 281898
rect 208794 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 209414 246454
rect 208794 246134 209414 246218
rect 208794 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 209414 246134
rect 208794 244084 209414 245898
rect 213294 711558 213914 711590
rect 213294 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 213914 711558
rect 213294 711238 213914 711322
rect 213294 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 213914 711238
rect 213294 682954 213914 711002
rect 213294 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 213914 682954
rect 213294 682634 213914 682718
rect 213294 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 213914 682634
rect 213294 646954 213914 682398
rect 213294 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 213914 646954
rect 213294 646634 213914 646718
rect 213294 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 213914 646634
rect 213294 610954 213914 646398
rect 213294 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 213914 610954
rect 213294 610634 213914 610718
rect 213294 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 213914 610634
rect 213294 574954 213914 610398
rect 213294 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 213914 574954
rect 213294 574634 213914 574718
rect 213294 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 213914 574634
rect 213294 538954 213914 574398
rect 213294 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 213914 538954
rect 213294 538634 213914 538718
rect 213294 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 213914 538634
rect 213294 502954 213914 538398
rect 213294 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 213914 502954
rect 213294 502634 213914 502718
rect 213294 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 213914 502634
rect 213294 466954 213914 502398
rect 213294 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 213914 466954
rect 213294 466634 213914 466718
rect 213294 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 213914 466634
rect 213294 430954 213914 466398
rect 213294 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 213914 430954
rect 213294 430634 213914 430718
rect 213294 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 213914 430634
rect 213294 394954 213914 430398
rect 213294 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 213914 394954
rect 213294 394634 213914 394718
rect 213294 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 213914 394634
rect 213294 358954 213914 394398
rect 213294 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 213914 358954
rect 213294 358634 213914 358718
rect 213294 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 213914 358634
rect 213294 322954 213914 358398
rect 213294 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 213914 322954
rect 213294 322634 213914 322718
rect 213294 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 213914 322634
rect 213294 286954 213914 322398
rect 213294 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 213914 286954
rect 213294 286634 213914 286718
rect 213294 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 213914 286634
rect 213294 250954 213914 286398
rect 213294 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 213914 250954
rect 213294 250634 213914 250718
rect 213294 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 213914 250634
rect 213294 244084 213914 250398
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 244084 218414 254898
rect 222294 705798 222914 711590
rect 222294 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 222914 705798
rect 222294 705478 222914 705562
rect 222294 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 222914 705478
rect 222294 691954 222914 705242
rect 222294 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 222914 691954
rect 222294 691634 222914 691718
rect 222294 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 222914 691634
rect 222294 655954 222914 691398
rect 222294 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 222914 655954
rect 222294 655634 222914 655718
rect 222294 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 222914 655634
rect 222294 619954 222914 655398
rect 222294 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 222914 619954
rect 222294 619634 222914 619718
rect 222294 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 222914 619634
rect 222294 583954 222914 619398
rect 222294 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 222914 583954
rect 222294 583634 222914 583718
rect 222294 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 222914 583634
rect 222294 547954 222914 583398
rect 222294 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 222914 547954
rect 222294 547634 222914 547718
rect 222294 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 222914 547634
rect 222294 511954 222914 547398
rect 222294 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 222914 511954
rect 222294 511634 222914 511718
rect 222294 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 222914 511634
rect 222294 475954 222914 511398
rect 222294 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 222914 475954
rect 222294 475634 222914 475718
rect 222294 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 222914 475634
rect 222294 439954 222914 475398
rect 222294 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 222914 439954
rect 222294 439634 222914 439718
rect 222294 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 222914 439634
rect 222294 403954 222914 439398
rect 222294 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 222914 403954
rect 222294 403634 222914 403718
rect 222294 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 222914 403634
rect 222294 367954 222914 403398
rect 222294 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 222914 367954
rect 222294 367634 222914 367718
rect 222294 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 222914 367634
rect 222294 331954 222914 367398
rect 222294 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 222914 331954
rect 222294 331634 222914 331718
rect 222294 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 222914 331634
rect 222294 295954 222914 331398
rect 222294 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 222914 295954
rect 222294 295634 222914 295718
rect 222294 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 222914 295634
rect 222294 259954 222914 295398
rect 222294 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 222914 259954
rect 222294 259634 222914 259718
rect 222294 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 222914 259634
rect 222294 244084 222914 259398
rect 226794 706758 227414 711590
rect 226794 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 227414 706758
rect 226794 706438 227414 706522
rect 226794 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 227414 706438
rect 226794 696454 227414 706202
rect 226794 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 227414 696454
rect 226794 696134 227414 696218
rect 226794 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 227414 696134
rect 226794 660454 227414 695898
rect 226794 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 227414 660454
rect 226794 660134 227414 660218
rect 226794 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 227414 660134
rect 226794 624454 227414 659898
rect 226794 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 227414 624454
rect 226794 624134 227414 624218
rect 226794 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 227414 624134
rect 226794 588454 227414 623898
rect 226794 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 227414 588454
rect 226794 588134 227414 588218
rect 226794 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 227414 588134
rect 226794 552454 227414 587898
rect 226794 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 227414 552454
rect 226794 552134 227414 552218
rect 226794 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 227414 552134
rect 226794 516454 227414 551898
rect 226794 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 227414 516454
rect 226794 516134 227414 516218
rect 226794 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 227414 516134
rect 226794 480454 227414 515898
rect 226794 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 227414 480454
rect 226794 480134 227414 480218
rect 226794 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 227414 480134
rect 226794 444454 227414 479898
rect 226794 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 227414 444454
rect 226794 444134 227414 444218
rect 226794 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 227414 444134
rect 226794 408454 227414 443898
rect 226794 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 227414 408454
rect 226794 408134 227414 408218
rect 226794 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 227414 408134
rect 226794 372454 227414 407898
rect 226794 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 227414 372454
rect 226794 372134 227414 372218
rect 226794 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 227414 372134
rect 226794 336454 227414 371898
rect 226794 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 227414 336454
rect 226794 336134 227414 336218
rect 226794 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 227414 336134
rect 226794 300454 227414 335898
rect 226794 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 227414 300454
rect 226794 300134 227414 300218
rect 226794 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 227414 300134
rect 226794 264454 227414 299898
rect 226794 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 227414 264454
rect 226794 264134 227414 264218
rect 226794 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 227414 264134
rect 226794 244084 227414 263898
rect 231294 707718 231914 711590
rect 231294 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 231914 707718
rect 231294 707398 231914 707482
rect 231294 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 231914 707398
rect 231294 700954 231914 707162
rect 231294 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 231914 700954
rect 231294 700634 231914 700718
rect 231294 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 231914 700634
rect 231294 664954 231914 700398
rect 231294 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 231914 664954
rect 231294 664634 231914 664718
rect 231294 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 231914 664634
rect 231294 628954 231914 664398
rect 231294 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 231914 628954
rect 231294 628634 231914 628718
rect 231294 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 231914 628634
rect 231294 592954 231914 628398
rect 231294 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 231914 592954
rect 231294 592634 231914 592718
rect 231294 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 231914 592634
rect 231294 556954 231914 592398
rect 231294 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 231914 556954
rect 231294 556634 231914 556718
rect 231294 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 231914 556634
rect 231294 520954 231914 556398
rect 231294 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 231914 520954
rect 231294 520634 231914 520718
rect 231294 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 231914 520634
rect 231294 484954 231914 520398
rect 231294 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 231914 484954
rect 231294 484634 231914 484718
rect 231294 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 231914 484634
rect 231294 448954 231914 484398
rect 231294 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 231914 448954
rect 231294 448634 231914 448718
rect 231294 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 231914 448634
rect 231294 412954 231914 448398
rect 231294 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 231914 412954
rect 231294 412634 231914 412718
rect 231294 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 231914 412634
rect 231294 376954 231914 412398
rect 231294 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 231914 376954
rect 231294 376634 231914 376718
rect 231294 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 231914 376634
rect 231294 340954 231914 376398
rect 231294 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 231914 340954
rect 231294 340634 231914 340718
rect 231294 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 231914 340634
rect 231294 304954 231914 340398
rect 231294 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 231914 304954
rect 231294 304634 231914 304718
rect 231294 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 231914 304634
rect 231294 268954 231914 304398
rect 231294 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 231914 268954
rect 231294 268634 231914 268718
rect 231294 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 231914 268634
rect 231294 244084 231914 268398
rect 235794 708678 236414 711590
rect 235794 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 236414 708678
rect 235794 708358 236414 708442
rect 235794 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 236414 708358
rect 235794 669454 236414 708122
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381454 236414 416898
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 273454 236414 308898
rect 235794 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 236414 273454
rect 235794 273134 236414 273218
rect 235794 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 236414 273134
rect 235794 244084 236414 272898
rect 240294 709638 240914 711590
rect 240294 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 240914 709638
rect 240294 709318 240914 709402
rect 240294 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 240914 709318
rect 240294 673954 240914 709082
rect 240294 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 240914 673954
rect 240294 673634 240914 673718
rect 240294 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 240914 673634
rect 240294 637954 240914 673398
rect 240294 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 240914 637954
rect 240294 637634 240914 637718
rect 240294 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 240914 637634
rect 240294 601954 240914 637398
rect 240294 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 240914 601954
rect 240294 601634 240914 601718
rect 240294 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 240914 601634
rect 240294 565954 240914 601398
rect 240294 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 240914 565954
rect 240294 565634 240914 565718
rect 240294 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 240914 565634
rect 240294 529954 240914 565398
rect 240294 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 240914 529954
rect 240294 529634 240914 529718
rect 240294 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 240914 529634
rect 240294 493954 240914 529398
rect 240294 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 240914 493954
rect 240294 493634 240914 493718
rect 240294 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 240914 493634
rect 240294 457954 240914 493398
rect 240294 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 240914 457954
rect 240294 457634 240914 457718
rect 240294 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 240914 457634
rect 240294 421954 240914 457398
rect 240294 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 240914 421954
rect 240294 421634 240914 421718
rect 240294 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 240914 421634
rect 240294 385954 240914 421398
rect 240294 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 240914 385954
rect 240294 385634 240914 385718
rect 240294 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 240914 385634
rect 240294 349954 240914 385398
rect 240294 349718 240326 349954
rect 240562 349718 240646 349954
rect 240882 349718 240914 349954
rect 240294 349634 240914 349718
rect 240294 349398 240326 349634
rect 240562 349398 240646 349634
rect 240882 349398 240914 349634
rect 240294 313954 240914 349398
rect 240294 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 240914 313954
rect 240294 313634 240914 313718
rect 240294 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 240914 313634
rect 240294 277954 240914 313398
rect 240294 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 240914 277954
rect 240294 277634 240914 277718
rect 240294 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 240914 277634
rect 240294 244084 240914 277398
rect 244794 710598 245414 711590
rect 244794 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 245414 710598
rect 244794 710278 245414 710362
rect 244794 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 245414 710278
rect 244794 678454 245414 710042
rect 244794 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 245414 678454
rect 244794 678134 245414 678218
rect 244794 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 245414 678134
rect 244794 642454 245414 677898
rect 244794 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 245414 642454
rect 244794 642134 245414 642218
rect 244794 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 245414 642134
rect 244794 606454 245414 641898
rect 244794 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 245414 606454
rect 244794 606134 245414 606218
rect 244794 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 245414 606134
rect 244794 570454 245414 605898
rect 244794 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 245414 570454
rect 244794 570134 245414 570218
rect 244794 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 245414 570134
rect 244794 534454 245414 569898
rect 244794 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 245414 534454
rect 244794 534134 245414 534218
rect 244794 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 245414 534134
rect 244794 498454 245414 533898
rect 244794 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 245414 498454
rect 244794 498134 245414 498218
rect 244794 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 245414 498134
rect 244794 462454 245414 497898
rect 244794 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 245414 462454
rect 244794 462134 245414 462218
rect 244794 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 245414 462134
rect 244794 426454 245414 461898
rect 244794 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 245414 426454
rect 244794 426134 245414 426218
rect 244794 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 245414 426134
rect 244794 390454 245414 425898
rect 244794 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 245414 390454
rect 244794 390134 245414 390218
rect 244794 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 245414 390134
rect 244794 354454 245414 389898
rect 244794 354218 244826 354454
rect 245062 354218 245146 354454
rect 245382 354218 245414 354454
rect 244794 354134 245414 354218
rect 244794 353898 244826 354134
rect 245062 353898 245146 354134
rect 245382 353898 245414 354134
rect 244794 318454 245414 353898
rect 244794 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 245414 318454
rect 244794 318134 245414 318218
rect 244794 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 245414 318134
rect 244794 282454 245414 317898
rect 244794 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 245414 282454
rect 244794 282134 245414 282218
rect 244794 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 245414 282134
rect 244794 246454 245414 281898
rect 244794 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 245414 246454
rect 244794 246134 245414 246218
rect 244794 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 245414 246134
rect 244794 244084 245414 245898
rect 249294 711558 249914 711590
rect 249294 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 249914 711558
rect 249294 711238 249914 711322
rect 249294 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 249914 711238
rect 249294 682954 249914 711002
rect 249294 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 249914 682954
rect 249294 682634 249914 682718
rect 249294 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 249914 682634
rect 249294 646954 249914 682398
rect 249294 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 249914 646954
rect 249294 646634 249914 646718
rect 249294 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 249914 646634
rect 249294 610954 249914 646398
rect 249294 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 249914 610954
rect 249294 610634 249914 610718
rect 249294 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 249914 610634
rect 249294 574954 249914 610398
rect 249294 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 249914 574954
rect 249294 574634 249914 574718
rect 249294 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 249914 574634
rect 249294 538954 249914 574398
rect 249294 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 249914 538954
rect 249294 538634 249914 538718
rect 249294 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 249914 538634
rect 249294 502954 249914 538398
rect 249294 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 249914 502954
rect 249294 502634 249914 502718
rect 249294 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 249914 502634
rect 249294 466954 249914 502398
rect 249294 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 249914 466954
rect 249294 466634 249914 466718
rect 249294 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 249914 466634
rect 249294 430954 249914 466398
rect 249294 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 249914 430954
rect 249294 430634 249914 430718
rect 249294 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 249914 430634
rect 249294 394954 249914 430398
rect 249294 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 249914 394954
rect 249294 394634 249914 394718
rect 249294 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 249914 394634
rect 249294 358954 249914 394398
rect 249294 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 249914 358954
rect 249294 358634 249914 358718
rect 249294 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 249914 358634
rect 249294 322954 249914 358398
rect 249294 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 249914 322954
rect 249294 322634 249914 322718
rect 249294 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 249914 322634
rect 249294 286954 249914 322398
rect 249294 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 249914 286954
rect 249294 286634 249914 286718
rect 249294 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 249914 286634
rect 249294 250954 249914 286398
rect 249294 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 249914 250954
rect 249294 250634 249914 250718
rect 249294 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 249914 250634
rect 249294 244084 249914 250398
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 291454 254414 326898
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 244084 254414 254898
rect 258294 705798 258914 711590
rect 258294 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 258914 705798
rect 258294 705478 258914 705562
rect 258294 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 258914 705478
rect 258294 691954 258914 705242
rect 258294 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 258914 691954
rect 258294 691634 258914 691718
rect 258294 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 258914 691634
rect 258294 655954 258914 691398
rect 258294 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 258914 655954
rect 258294 655634 258914 655718
rect 258294 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 258914 655634
rect 258294 619954 258914 655398
rect 258294 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 258914 619954
rect 258294 619634 258914 619718
rect 258294 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 258914 619634
rect 258294 583954 258914 619398
rect 258294 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 258914 583954
rect 258294 583634 258914 583718
rect 258294 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 258914 583634
rect 258294 547954 258914 583398
rect 258294 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 258914 547954
rect 258294 547634 258914 547718
rect 258294 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 258914 547634
rect 258294 511954 258914 547398
rect 258294 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 258914 511954
rect 258294 511634 258914 511718
rect 258294 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 258914 511634
rect 258294 475954 258914 511398
rect 258294 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 258914 475954
rect 258294 475634 258914 475718
rect 258294 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 258914 475634
rect 258294 439954 258914 475398
rect 258294 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 258914 439954
rect 258294 439634 258914 439718
rect 258294 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 258914 439634
rect 258294 403954 258914 439398
rect 258294 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 258914 403954
rect 258294 403634 258914 403718
rect 258294 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 258914 403634
rect 258294 367954 258914 403398
rect 258294 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 258914 367954
rect 258294 367634 258914 367718
rect 258294 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 258914 367634
rect 258294 331954 258914 367398
rect 258294 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 258914 331954
rect 258294 331634 258914 331718
rect 258294 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 258914 331634
rect 258294 295954 258914 331398
rect 258294 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 258914 295954
rect 258294 295634 258914 295718
rect 258294 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 258914 295634
rect 258294 259954 258914 295398
rect 258294 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 258914 259954
rect 258294 259634 258914 259718
rect 258294 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 258914 259634
rect 258294 244084 258914 259398
rect 262794 706758 263414 711590
rect 262794 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 263414 706758
rect 262794 706438 263414 706522
rect 262794 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 263414 706438
rect 262794 696454 263414 706202
rect 262794 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 263414 696454
rect 262794 696134 263414 696218
rect 262794 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 263414 696134
rect 262794 660454 263414 695898
rect 262794 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 263414 660454
rect 262794 660134 263414 660218
rect 262794 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 263414 660134
rect 262794 624454 263414 659898
rect 262794 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 263414 624454
rect 262794 624134 263414 624218
rect 262794 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 263414 624134
rect 262794 588454 263414 623898
rect 262794 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 263414 588454
rect 262794 588134 263414 588218
rect 262794 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 263414 588134
rect 262794 552454 263414 587898
rect 262794 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 263414 552454
rect 262794 552134 263414 552218
rect 262794 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 263414 552134
rect 262794 516454 263414 551898
rect 262794 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 263414 516454
rect 262794 516134 263414 516218
rect 262794 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 263414 516134
rect 262794 480454 263414 515898
rect 262794 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 263414 480454
rect 262794 480134 263414 480218
rect 262794 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 263414 480134
rect 262794 444454 263414 479898
rect 262794 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 263414 444454
rect 262794 444134 263414 444218
rect 262794 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 263414 444134
rect 262794 408454 263414 443898
rect 262794 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 263414 408454
rect 262794 408134 263414 408218
rect 262794 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 263414 408134
rect 262794 372454 263414 407898
rect 262794 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 263414 372454
rect 262794 372134 263414 372218
rect 262794 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 263414 372134
rect 262794 336454 263414 371898
rect 262794 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 263414 336454
rect 262794 336134 263414 336218
rect 262794 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 263414 336134
rect 262794 300454 263414 335898
rect 262794 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 263414 300454
rect 262794 300134 263414 300218
rect 262794 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 263414 300134
rect 262794 264454 263414 299898
rect 262794 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 263414 264454
rect 262794 264134 263414 264218
rect 262794 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 263414 264134
rect 262794 244084 263414 263898
rect 267294 707718 267914 711590
rect 267294 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 267914 707718
rect 267294 707398 267914 707482
rect 267294 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 267914 707398
rect 267294 700954 267914 707162
rect 267294 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 267914 700954
rect 267294 700634 267914 700718
rect 267294 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 267914 700634
rect 267294 664954 267914 700398
rect 267294 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 267914 664954
rect 267294 664634 267914 664718
rect 267294 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 267914 664634
rect 267294 628954 267914 664398
rect 267294 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 267914 628954
rect 267294 628634 267914 628718
rect 267294 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 267914 628634
rect 267294 592954 267914 628398
rect 267294 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 267914 592954
rect 267294 592634 267914 592718
rect 267294 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 267914 592634
rect 267294 556954 267914 592398
rect 267294 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 267914 556954
rect 267294 556634 267914 556718
rect 267294 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 267914 556634
rect 267294 520954 267914 556398
rect 267294 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 267914 520954
rect 267294 520634 267914 520718
rect 267294 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 267914 520634
rect 267294 484954 267914 520398
rect 267294 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 267914 484954
rect 267294 484634 267914 484718
rect 267294 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 267914 484634
rect 267294 448954 267914 484398
rect 267294 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 267914 448954
rect 267294 448634 267914 448718
rect 267294 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 267914 448634
rect 267294 412954 267914 448398
rect 267294 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 267914 412954
rect 267294 412634 267914 412718
rect 267294 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 267914 412634
rect 267294 376954 267914 412398
rect 267294 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 267914 376954
rect 267294 376634 267914 376718
rect 267294 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 267914 376634
rect 267294 340954 267914 376398
rect 267294 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 267914 340954
rect 267294 340634 267914 340718
rect 267294 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 267914 340634
rect 267294 304954 267914 340398
rect 267294 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 267914 304954
rect 267294 304634 267914 304718
rect 267294 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 267914 304634
rect 267294 268954 267914 304398
rect 267294 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 267914 268954
rect 267294 268634 267914 268718
rect 267294 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 267914 268634
rect 267294 244084 267914 268398
rect 271794 708678 272414 711590
rect 271794 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 272414 708678
rect 271794 708358 272414 708442
rect 271794 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 272414 708358
rect 271794 669454 272414 708122
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 345454 272414 380898
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 273454 272414 308898
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 244084 272414 272898
rect 276294 709638 276914 711590
rect 276294 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 276914 709638
rect 276294 709318 276914 709402
rect 276294 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 276914 709318
rect 276294 673954 276914 709082
rect 276294 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 276914 673954
rect 276294 673634 276914 673718
rect 276294 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 276914 673634
rect 276294 637954 276914 673398
rect 276294 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 276914 637954
rect 276294 637634 276914 637718
rect 276294 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 276914 637634
rect 276294 601954 276914 637398
rect 276294 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 276914 601954
rect 276294 601634 276914 601718
rect 276294 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 276914 601634
rect 276294 565954 276914 601398
rect 276294 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 276914 565954
rect 276294 565634 276914 565718
rect 276294 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 276914 565634
rect 276294 529954 276914 565398
rect 276294 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 276914 529954
rect 276294 529634 276914 529718
rect 276294 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 276914 529634
rect 276294 493954 276914 529398
rect 276294 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 276914 493954
rect 276294 493634 276914 493718
rect 276294 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 276914 493634
rect 276294 457954 276914 493398
rect 276294 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 276914 457954
rect 276294 457634 276914 457718
rect 276294 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 276914 457634
rect 276294 421954 276914 457398
rect 276294 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 276914 421954
rect 276294 421634 276914 421718
rect 276294 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 276914 421634
rect 276294 385954 276914 421398
rect 276294 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 276914 385954
rect 276294 385634 276914 385718
rect 276294 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 276914 385634
rect 276294 349954 276914 385398
rect 276294 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 276914 349954
rect 276294 349634 276914 349718
rect 276294 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 276914 349634
rect 276294 313954 276914 349398
rect 276294 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 276914 313954
rect 276294 313634 276914 313718
rect 276294 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 276914 313634
rect 276294 277954 276914 313398
rect 276294 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 276914 277954
rect 276294 277634 276914 277718
rect 276294 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 276914 277634
rect 276294 244084 276914 277398
rect 280794 710598 281414 711590
rect 280794 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 281414 710598
rect 280794 710278 281414 710362
rect 280794 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 281414 710278
rect 280794 678454 281414 710042
rect 280794 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 281414 678454
rect 280794 678134 281414 678218
rect 280794 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 281414 678134
rect 280794 642454 281414 677898
rect 280794 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 281414 642454
rect 280794 642134 281414 642218
rect 280794 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 281414 642134
rect 280794 606454 281414 641898
rect 280794 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 281414 606454
rect 280794 606134 281414 606218
rect 280794 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 281414 606134
rect 280794 570454 281414 605898
rect 280794 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 281414 570454
rect 280794 570134 281414 570218
rect 280794 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 281414 570134
rect 280794 534454 281414 569898
rect 280794 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 281414 534454
rect 280794 534134 281414 534218
rect 280794 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 281414 534134
rect 280794 498454 281414 533898
rect 280794 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 281414 498454
rect 280794 498134 281414 498218
rect 280794 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 281414 498134
rect 280794 462454 281414 497898
rect 280794 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 281414 462454
rect 280794 462134 281414 462218
rect 280794 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 281414 462134
rect 280794 426454 281414 461898
rect 280794 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 281414 426454
rect 280794 426134 281414 426218
rect 280794 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 281414 426134
rect 280794 390454 281414 425898
rect 280794 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 281414 390454
rect 280794 390134 281414 390218
rect 280794 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 281414 390134
rect 280794 354454 281414 389898
rect 280794 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 281414 354454
rect 280794 354134 281414 354218
rect 280794 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 281414 354134
rect 280794 318454 281414 353898
rect 280794 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 281414 318454
rect 280794 318134 281414 318218
rect 280794 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 281414 318134
rect 280794 282454 281414 317898
rect 280794 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 281414 282454
rect 280794 282134 281414 282218
rect 280794 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 281414 282134
rect 280794 246454 281414 281898
rect 280794 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 281414 246454
rect 280794 246134 281414 246218
rect 280794 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 281414 246134
rect 280794 244084 281414 245898
rect 285294 711558 285914 711590
rect 285294 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 285914 711558
rect 285294 711238 285914 711322
rect 285294 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 285914 711238
rect 285294 682954 285914 711002
rect 285294 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 285914 682954
rect 285294 682634 285914 682718
rect 285294 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 285914 682634
rect 285294 646954 285914 682398
rect 285294 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 285914 646954
rect 285294 646634 285914 646718
rect 285294 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 285914 646634
rect 285294 610954 285914 646398
rect 285294 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 285914 610954
rect 285294 610634 285914 610718
rect 285294 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 285914 610634
rect 285294 574954 285914 610398
rect 285294 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 285914 574954
rect 285294 574634 285914 574718
rect 285294 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 285914 574634
rect 285294 538954 285914 574398
rect 285294 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 285914 538954
rect 285294 538634 285914 538718
rect 285294 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 285914 538634
rect 285294 502954 285914 538398
rect 285294 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 285914 502954
rect 285294 502634 285914 502718
rect 285294 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 285914 502634
rect 285294 466954 285914 502398
rect 285294 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 285914 466954
rect 285294 466634 285914 466718
rect 285294 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 285914 466634
rect 285294 430954 285914 466398
rect 285294 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 285914 430954
rect 285294 430634 285914 430718
rect 285294 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 285914 430634
rect 285294 394954 285914 430398
rect 285294 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 285914 394954
rect 285294 394634 285914 394718
rect 285294 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 285914 394634
rect 285294 358954 285914 394398
rect 285294 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 285914 358954
rect 285294 358634 285914 358718
rect 285294 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 285914 358634
rect 285294 322954 285914 358398
rect 285294 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 285914 322954
rect 285294 322634 285914 322718
rect 285294 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 285914 322634
rect 285294 286954 285914 322398
rect 285294 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 285914 286954
rect 285294 286634 285914 286718
rect 285294 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 285914 286634
rect 285294 250954 285914 286398
rect 285294 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 285914 250954
rect 285294 250634 285914 250718
rect 285294 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 285914 250634
rect 285294 244084 285914 250398
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 244084 290414 254898
rect 294294 705798 294914 711590
rect 294294 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 294914 705798
rect 294294 705478 294914 705562
rect 294294 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 294914 705478
rect 294294 691954 294914 705242
rect 294294 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 294914 691954
rect 294294 691634 294914 691718
rect 294294 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 294914 691634
rect 294294 655954 294914 691398
rect 294294 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 294914 655954
rect 294294 655634 294914 655718
rect 294294 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 294914 655634
rect 294294 619954 294914 655398
rect 294294 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 294914 619954
rect 294294 619634 294914 619718
rect 294294 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 294914 619634
rect 294294 583954 294914 619398
rect 294294 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 294914 583954
rect 294294 583634 294914 583718
rect 294294 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 294914 583634
rect 294294 547954 294914 583398
rect 294294 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 294914 547954
rect 294294 547634 294914 547718
rect 294294 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 294914 547634
rect 294294 511954 294914 547398
rect 294294 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 294914 511954
rect 294294 511634 294914 511718
rect 294294 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 294914 511634
rect 294294 475954 294914 511398
rect 294294 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 294914 475954
rect 294294 475634 294914 475718
rect 294294 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 294914 475634
rect 294294 439954 294914 475398
rect 294294 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 294914 439954
rect 294294 439634 294914 439718
rect 294294 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 294914 439634
rect 294294 403954 294914 439398
rect 294294 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 294914 403954
rect 294294 403634 294914 403718
rect 294294 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 294914 403634
rect 294294 367954 294914 403398
rect 294294 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 294914 367954
rect 294294 367634 294914 367718
rect 294294 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 294914 367634
rect 294294 331954 294914 367398
rect 294294 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 294914 331954
rect 294294 331634 294914 331718
rect 294294 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 294914 331634
rect 294294 295954 294914 331398
rect 294294 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 294914 295954
rect 294294 295634 294914 295718
rect 294294 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 294914 295634
rect 294294 259954 294914 295398
rect 294294 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 294914 259954
rect 294294 259634 294914 259718
rect 294294 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 294914 259634
rect 294294 244084 294914 259398
rect 298794 706758 299414 711590
rect 298794 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 299414 706758
rect 298794 706438 299414 706522
rect 298794 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 299414 706438
rect 298794 696454 299414 706202
rect 298794 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 299414 696454
rect 298794 696134 299414 696218
rect 298794 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 299414 696134
rect 298794 660454 299414 695898
rect 298794 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 299414 660454
rect 298794 660134 299414 660218
rect 298794 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 299414 660134
rect 298794 624454 299414 659898
rect 298794 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 299414 624454
rect 298794 624134 299414 624218
rect 298794 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 299414 624134
rect 298794 588454 299414 623898
rect 298794 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 299414 588454
rect 298794 588134 299414 588218
rect 298794 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 299414 588134
rect 298794 552454 299414 587898
rect 298794 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 299414 552454
rect 298794 552134 299414 552218
rect 298794 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 299414 552134
rect 298794 516454 299414 551898
rect 298794 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 299414 516454
rect 298794 516134 299414 516218
rect 298794 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 299414 516134
rect 298794 480454 299414 515898
rect 298794 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 299414 480454
rect 298794 480134 299414 480218
rect 298794 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 299414 480134
rect 298794 444454 299414 479898
rect 298794 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 299414 444454
rect 298794 444134 299414 444218
rect 298794 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 299414 444134
rect 298794 408454 299414 443898
rect 298794 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 299414 408454
rect 298794 408134 299414 408218
rect 298794 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 299414 408134
rect 298794 372454 299414 407898
rect 298794 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 299414 372454
rect 298794 372134 299414 372218
rect 298794 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 299414 372134
rect 298794 336454 299414 371898
rect 298794 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 299414 336454
rect 298794 336134 299414 336218
rect 298794 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 299414 336134
rect 298794 300454 299414 335898
rect 298794 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 299414 300454
rect 298794 300134 299414 300218
rect 298794 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 299414 300134
rect 298794 264454 299414 299898
rect 298794 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 299414 264454
rect 298794 264134 299414 264218
rect 298794 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 299414 264134
rect 298794 244084 299414 263898
rect 303294 707718 303914 711590
rect 303294 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 303914 707718
rect 303294 707398 303914 707482
rect 303294 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 303914 707398
rect 303294 700954 303914 707162
rect 303294 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 303914 700954
rect 303294 700634 303914 700718
rect 303294 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 303914 700634
rect 303294 664954 303914 700398
rect 303294 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 303914 664954
rect 303294 664634 303914 664718
rect 303294 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 303914 664634
rect 303294 628954 303914 664398
rect 303294 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 303914 628954
rect 303294 628634 303914 628718
rect 303294 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 303914 628634
rect 303294 592954 303914 628398
rect 303294 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 303914 592954
rect 303294 592634 303914 592718
rect 303294 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 303914 592634
rect 303294 556954 303914 592398
rect 303294 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 303914 556954
rect 303294 556634 303914 556718
rect 303294 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 303914 556634
rect 303294 520954 303914 556398
rect 303294 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 303914 520954
rect 303294 520634 303914 520718
rect 303294 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 303914 520634
rect 303294 484954 303914 520398
rect 303294 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 303914 484954
rect 303294 484634 303914 484718
rect 303294 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 303914 484634
rect 303294 448954 303914 484398
rect 303294 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 303914 448954
rect 303294 448634 303914 448718
rect 303294 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 303914 448634
rect 303294 412954 303914 448398
rect 303294 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 303914 412954
rect 303294 412634 303914 412718
rect 303294 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 303914 412634
rect 303294 376954 303914 412398
rect 303294 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 303914 376954
rect 303294 376634 303914 376718
rect 303294 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 303914 376634
rect 303294 340954 303914 376398
rect 303294 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 303914 340954
rect 303294 340634 303914 340718
rect 303294 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 303914 340634
rect 303294 304954 303914 340398
rect 303294 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 303914 304954
rect 303294 304634 303914 304718
rect 303294 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 303914 304634
rect 303294 268954 303914 304398
rect 303294 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 303914 268954
rect 303294 268634 303914 268718
rect 303294 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 303914 268634
rect 303294 244084 303914 268398
rect 307794 708678 308414 711590
rect 307794 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 308414 708678
rect 307794 708358 308414 708442
rect 307794 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 308414 708358
rect 307794 669454 308414 708122
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 244084 308414 272898
rect 312294 709638 312914 711590
rect 312294 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 312914 709638
rect 312294 709318 312914 709402
rect 312294 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 312914 709318
rect 312294 673954 312914 709082
rect 312294 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 312914 673954
rect 312294 673634 312914 673718
rect 312294 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 312914 673634
rect 312294 637954 312914 673398
rect 312294 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 312914 637954
rect 312294 637634 312914 637718
rect 312294 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 312914 637634
rect 312294 601954 312914 637398
rect 312294 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 312914 601954
rect 312294 601634 312914 601718
rect 312294 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 312914 601634
rect 312294 565954 312914 601398
rect 312294 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 312914 565954
rect 312294 565634 312914 565718
rect 312294 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 312914 565634
rect 312294 529954 312914 565398
rect 312294 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 312914 529954
rect 312294 529634 312914 529718
rect 312294 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 312914 529634
rect 312294 493954 312914 529398
rect 312294 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 312914 493954
rect 312294 493634 312914 493718
rect 312294 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 312914 493634
rect 312294 457954 312914 493398
rect 312294 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 312914 457954
rect 312294 457634 312914 457718
rect 312294 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 312914 457634
rect 312294 421954 312914 457398
rect 312294 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 312914 421954
rect 312294 421634 312914 421718
rect 312294 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 312914 421634
rect 312294 385954 312914 421398
rect 312294 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 312914 385954
rect 312294 385634 312914 385718
rect 312294 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 312914 385634
rect 312294 349954 312914 385398
rect 312294 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 312914 349954
rect 312294 349634 312914 349718
rect 312294 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 312914 349634
rect 312294 313954 312914 349398
rect 312294 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 312914 313954
rect 312294 313634 312914 313718
rect 312294 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 312914 313634
rect 312294 277954 312914 313398
rect 312294 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 312914 277954
rect 312294 277634 312914 277718
rect 312294 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 312914 277634
rect 312294 244084 312914 277398
rect 316794 710598 317414 711590
rect 316794 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 317414 710598
rect 316794 710278 317414 710362
rect 316794 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 317414 710278
rect 316794 678454 317414 710042
rect 316794 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 317414 678454
rect 316794 678134 317414 678218
rect 316794 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 317414 678134
rect 316794 642454 317414 677898
rect 316794 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 317414 642454
rect 316794 642134 317414 642218
rect 316794 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 317414 642134
rect 316794 606454 317414 641898
rect 316794 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 317414 606454
rect 316794 606134 317414 606218
rect 316794 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 317414 606134
rect 316794 570454 317414 605898
rect 316794 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 317414 570454
rect 316794 570134 317414 570218
rect 316794 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 317414 570134
rect 316794 534454 317414 569898
rect 316794 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 317414 534454
rect 316794 534134 317414 534218
rect 316794 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 317414 534134
rect 316794 498454 317414 533898
rect 316794 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 317414 498454
rect 316794 498134 317414 498218
rect 316794 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 317414 498134
rect 316794 462454 317414 497898
rect 316794 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 317414 462454
rect 316794 462134 317414 462218
rect 316794 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 317414 462134
rect 316794 426454 317414 461898
rect 316794 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 317414 426454
rect 316794 426134 317414 426218
rect 316794 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 317414 426134
rect 316794 390454 317414 425898
rect 316794 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 317414 390454
rect 316794 390134 317414 390218
rect 316794 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 317414 390134
rect 316794 354454 317414 389898
rect 316794 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 317414 354454
rect 316794 354134 317414 354218
rect 316794 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 317414 354134
rect 316794 318454 317414 353898
rect 316794 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 317414 318454
rect 316794 318134 317414 318218
rect 316794 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 317414 318134
rect 316794 282454 317414 317898
rect 316794 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 317414 282454
rect 316794 282134 317414 282218
rect 316794 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 317414 282134
rect 316794 246454 317414 281898
rect 316794 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 317414 246454
rect 316794 246134 317414 246218
rect 316794 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 317414 246134
rect 316794 244084 317414 245898
rect 321294 711558 321914 711590
rect 321294 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 321914 711558
rect 321294 711238 321914 711322
rect 321294 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 321914 711238
rect 321294 682954 321914 711002
rect 321294 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 321914 682954
rect 321294 682634 321914 682718
rect 321294 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 321914 682634
rect 321294 646954 321914 682398
rect 321294 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 321914 646954
rect 321294 646634 321914 646718
rect 321294 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 321914 646634
rect 321294 610954 321914 646398
rect 321294 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 321914 610954
rect 321294 610634 321914 610718
rect 321294 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 321914 610634
rect 321294 574954 321914 610398
rect 321294 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 321914 574954
rect 321294 574634 321914 574718
rect 321294 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 321914 574634
rect 321294 538954 321914 574398
rect 321294 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 321914 538954
rect 321294 538634 321914 538718
rect 321294 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 321914 538634
rect 321294 502954 321914 538398
rect 321294 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 321914 502954
rect 321294 502634 321914 502718
rect 321294 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 321914 502634
rect 321294 466954 321914 502398
rect 321294 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 321914 466954
rect 321294 466634 321914 466718
rect 321294 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 321914 466634
rect 321294 430954 321914 466398
rect 321294 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 321914 430954
rect 321294 430634 321914 430718
rect 321294 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 321914 430634
rect 321294 394954 321914 430398
rect 321294 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 321914 394954
rect 321294 394634 321914 394718
rect 321294 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 321914 394634
rect 321294 358954 321914 394398
rect 321294 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 321914 358954
rect 321294 358634 321914 358718
rect 321294 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 321914 358634
rect 321294 322954 321914 358398
rect 321294 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 321914 322954
rect 321294 322634 321914 322718
rect 321294 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 321914 322634
rect 321294 286954 321914 322398
rect 321294 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 321914 286954
rect 321294 286634 321914 286718
rect 321294 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 321914 286634
rect 321294 250954 321914 286398
rect 321294 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 321914 250954
rect 321294 250634 321914 250718
rect 321294 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 321914 250634
rect 321294 244084 321914 250398
rect 325794 704838 326414 711590
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 244084 326414 254898
rect 330294 705798 330914 711590
rect 330294 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 330914 705798
rect 330294 705478 330914 705562
rect 330294 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 330914 705478
rect 330294 691954 330914 705242
rect 330294 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 330914 691954
rect 330294 691634 330914 691718
rect 330294 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 330914 691634
rect 330294 655954 330914 691398
rect 330294 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 330914 655954
rect 330294 655634 330914 655718
rect 330294 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 330914 655634
rect 330294 619954 330914 655398
rect 330294 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 330914 619954
rect 330294 619634 330914 619718
rect 330294 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 330914 619634
rect 330294 583954 330914 619398
rect 330294 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 330914 583954
rect 330294 583634 330914 583718
rect 330294 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 330914 583634
rect 330294 547954 330914 583398
rect 330294 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 330914 547954
rect 330294 547634 330914 547718
rect 330294 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 330914 547634
rect 330294 511954 330914 547398
rect 330294 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 330914 511954
rect 330294 511634 330914 511718
rect 330294 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 330914 511634
rect 330294 475954 330914 511398
rect 330294 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 330914 475954
rect 330294 475634 330914 475718
rect 330294 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 330914 475634
rect 330294 439954 330914 475398
rect 330294 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 330914 439954
rect 330294 439634 330914 439718
rect 330294 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 330914 439634
rect 330294 403954 330914 439398
rect 330294 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 330914 403954
rect 330294 403634 330914 403718
rect 330294 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 330914 403634
rect 330294 367954 330914 403398
rect 330294 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 330914 367954
rect 330294 367634 330914 367718
rect 330294 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 330914 367634
rect 330294 331954 330914 367398
rect 330294 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 330914 331954
rect 330294 331634 330914 331718
rect 330294 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 330914 331634
rect 330294 295954 330914 331398
rect 330294 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 330914 295954
rect 330294 295634 330914 295718
rect 330294 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 330914 295634
rect 330294 259954 330914 295398
rect 330294 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 330914 259954
rect 330294 259634 330914 259718
rect 330294 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 330914 259634
rect 330294 244084 330914 259398
rect 334794 706758 335414 711590
rect 334794 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 335414 706758
rect 334794 706438 335414 706522
rect 334794 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 335414 706438
rect 334794 696454 335414 706202
rect 334794 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 335414 696454
rect 334794 696134 335414 696218
rect 334794 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 335414 696134
rect 334794 660454 335414 695898
rect 334794 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 335414 660454
rect 334794 660134 335414 660218
rect 334794 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 335414 660134
rect 334794 624454 335414 659898
rect 334794 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 335414 624454
rect 334794 624134 335414 624218
rect 334794 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 335414 624134
rect 334794 588454 335414 623898
rect 334794 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 335414 588454
rect 334794 588134 335414 588218
rect 334794 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 335414 588134
rect 334794 552454 335414 587898
rect 334794 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 335414 552454
rect 334794 552134 335414 552218
rect 334794 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 335414 552134
rect 334794 516454 335414 551898
rect 334794 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 335414 516454
rect 334794 516134 335414 516218
rect 334794 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 335414 516134
rect 334794 480454 335414 515898
rect 334794 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 335414 480454
rect 334794 480134 335414 480218
rect 334794 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 335414 480134
rect 334794 444454 335414 479898
rect 334794 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 335414 444454
rect 334794 444134 335414 444218
rect 334794 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 335414 444134
rect 334794 408454 335414 443898
rect 334794 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 335414 408454
rect 334794 408134 335414 408218
rect 334794 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 335414 408134
rect 334794 372454 335414 407898
rect 334794 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 335414 372454
rect 334794 372134 335414 372218
rect 334794 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 335414 372134
rect 334794 336454 335414 371898
rect 334794 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 335414 336454
rect 334794 336134 335414 336218
rect 334794 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 335414 336134
rect 334794 300454 335414 335898
rect 334794 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 335414 300454
rect 334794 300134 335414 300218
rect 334794 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 335414 300134
rect 334794 264454 335414 299898
rect 334794 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 335414 264454
rect 334794 264134 335414 264218
rect 334794 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 335414 264134
rect 334794 244084 335414 263898
rect 339294 707718 339914 711590
rect 339294 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 339914 707718
rect 339294 707398 339914 707482
rect 339294 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 339914 707398
rect 339294 700954 339914 707162
rect 339294 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 339914 700954
rect 339294 700634 339914 700718
rect 339294 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 339914 700634
rect 339294 664954 339914 700398
rect 339294 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 339914 664954
rect 339294 664634 339914 664718
rect 339294 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 339914 664634
rect 339294 628954 339914 664398
rect 339294 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 339914 628954
rect 339294 628634 339914 628718
rect 339294 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 339914 628634
rect 339294 592954 339914 628398
rect 339294 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 339914 592954
rect 339294 592634 339914 592718
rect 339294 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 339914 592634
rect 339294 556954 339914 592398
rect 339294 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 339914 556954
rect 339294 556634 339914 556718
rect 339294 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 339914 556634
rect 339294 520954 339914 556398
rect 339294 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 339914 520954
rect 339294 520634 339914 520718
rect 339294 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 339914 520634
rect 339294 484954 339914 520398
rect 339294 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 339914 484954
rect 339294 484634 339914 484718
rect 339294 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 339914 484634
rect 339294 448954 339914 484398
rect 339294 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 339914 448954
rect 339294 448634 339914 448718
rect 339294 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 339914 448634
rect 339294 412954 339914 448398
rect 339294 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 339914 412954
rect 339294 412634 339914 412718
rect 339294 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 339914 412634
rect 339294 376954 339914 412398
rect 339294 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 339914 376954
rect 339294 376634 339914 376718
rect 339294 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 339914 376634
rect 339294 340954 339914 376398
rect 339294 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 339914 340954
rect 339294 340634 339914 340718
rect 339294 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 339914 340634
rect 339294 304954 339914 340398
rect 339294 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 339914 304954
rect 339294 304634 339914 304718
rect 339294 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 339914 304634
rect 339294 268954 339914 304398
rect 339294 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 339914 268954
rect 339294 268634 339914 268718
rect 339294 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 339914 268634
rect 339294 244084 339914 268398
rect 343794 708678 344414 711590
rect 343794 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 344414 708678
rect 343794 708358 344414 708442
rect 343794 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 344414 708358
rect 343794 669454 344414 708122
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 244084 344414 272898
rect 348294 709638 348914 711590
rect 348294 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 348914 709638
rect 348294 709318 348914 709402
rect 348294 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 348914 709318
rect 348294 673954 348914 709082
rect 348294 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 348914 673954
rect 348294 673634 348914 673718
rect 348294 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 348914 673634
rect 348294 637954 348914 673398
rect 348294 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 348914 637954
rect 348294 637634 348914 637718
rect 348294 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 348914 637634
rect 348294 601954 348914 637398
rect 348294 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 348914 601954
rect 348294 601634 348914 601718
rect 348294 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 348914 601634
rect 348294 565954 348914 601398
rect 348294 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 348914 565954
rect 348294 565634 348914 565718
rect 348294 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 348914 565634
rect 348294 529954 348914 565398
rect 348294 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 348914 529954
rect 348294 529634 348914 529718
rect 348294 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 348914 529634
rect 348294 493954 348914 529398
rect 348294 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 348914 493954
rect 348294 493634 348914 493718
rect 348294 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 348914 493634
rect 348294 457954 348914 493398
rect 348294 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 348914 457954
rect 348294 457634 348914 457718
rect 348294 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 348914 457634
rect 348294 421954 348914 457398
rect 348294 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 348914 421954
rect 348294 421634 348914 421718
rect 348294 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 348914 421634
rect 348294 385954 348914 421398
rect 348294 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 348914 385954
rect 348294 385634 348914 385718
rect 348294 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 348914 385634
rect 348294 349954 348914 385398
rect 348294 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 348914 349954
rect 348294 349634 348914 349718
rect 348294 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 348914 349634
rect 348294 313954 348914 349398
rect 348294 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 348914 313954
rect 348294 313634 348914 313718
rect 348294 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 348914 313634
rect 348294 277954 348914 313398
rect 348294 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 348914 277954
rect 348294 277634 348914 277718
rect 348294 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 348914 277634
rect 348294 244084 348914 277398
rect 352794 710598 353414 711590
rect 352794 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 353414 710598
rect 352794 710278 353414 710362
rect 352794 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 353414 710278
rect 352794 678454 353414 710042
rect 352794 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 353414 678454
rect 352794 678134 353414 678218
rect 352794 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 353414 678134
rect 352794 642454 353414 677898
rect 352794 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 353414 642454
rect 352794 642134 353414 642218
rect 352794 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 353414 642134
rect 352794 606454 353414 641898
rect 352794 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 353414 606454
rect 352794 606134 353414 606218
rect 352794 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 353414 606134
rect 352794 570454 353414 605898
rect 352794 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 353414 570454
rect 352794 570134 353414 570218
rect 352794 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 353414 570134
rect 352794 534454 353414 569898
rect 352794 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 353414 534454
rect 352794 534134 353414 534218
rect 352794 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 353414 534134
rect 352794 498454 353414 533898
rect 352794 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 353414 498454
rect 352794 498134 353414 498218
rect 352794 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 353414 498134
rect 352794 462454 353414 497898
rect 352794 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 353414 462454
rect 352794 462134 353414 462218
rect 352794 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 353414 462134
rect 352794 426454 353414 461898
rect 352794 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 353414 426454
rect 352794 426134 353414 426218
rect 352794 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 353414 426134
rect 352794 390454 353414 425898
rect 352794 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 353414 390454
rect 352794 390134 353414 390218
rect 352794 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 353414 390134
rect 352794 354454 353414 389898
rect 352794 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 353414 354454
rect 352794 354134 353414 354218
rect 352794 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 353414 354134
rect 352794 318454 353414 353898
rect 352794 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 353414 318454
rect 352794 318134 353414 318218
rect 352794 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 353414 318134
rect 352794 282454 353414 317898
rect 352794 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 353414 282454
rect 352794 282134 353414 282218
rect 352794 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 353414 282134
rect 352794 246454 353414 281898
rect 352794 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 353414 246454
rect 352794 246134 353414 246218
rect 352794 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 353414 246134
rect 352794 244084 353414 245898
rect 357294 711558 357914 711590
rect 357294 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 357914 711558
rect 357294 711238 357914 711322
rect 357294 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 357914 711238
rect 357294 682954 357914 711002
rect 357294 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 357914 682954
rect 357294 682634 357914 682718
rect 357294 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 357914 682634
rect 357294 646954 357914 682398
rect 357294 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 357914 646954
rect 357294 646634 357914 646718
rect 357294 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 357914 646634
rect 357294 610954 357914 646398
rect 357294 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 357914 610954
rect 357294 610634 357914 610718
rect 357294 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 357914 610634
rect 357294 574954 357914 610398
rect 357294 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 357914 574954
rect 357294 574634 357914 574718
rect 357294 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 357914 574634
rect 357294 538954 357914 574398
rect 357294 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 357914 538954
rect 357294 538634 357914 538718
rect 357294 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 357914 538634
rect 357294 502954 357914 538398
rect 357294 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 357914 502954
rect 357294 502634 357914 502718
rect 357294 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 357914 502634
rect 357294 466954 357914 502398
rect 357294 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 357914 466954
rect 357294 466634 357914 466718
rect 357294 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 357914 466634
rect 357294 430954 357914 466398
rect 357294 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 357914 430954
rect 357294 430634 357914 430718
rect 357294 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 357914 430634
rect 357294 394954 357914 430398
rect 357294 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 357914 394954
rect 357294 394634 357914 394718
rect 357294 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 357914 394634
rect 357294 358954 357914 394398
rect 357294 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 357914 358954
rect 357294 358634 357914 358718
rect 357294 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 357914 358634
rect 357294 322954 357914 358398
rect 357294 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 357914 322954
rect 357294 322634 357914 322718
rect 357294 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 357914 322634
rect 357294 286954 357914 322398
rect 357294 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 357914 286954
rect 357294 286634 357914 286718
rect 357294 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 357914 286634
rect 357294 250954 357914 286398
rect 357294 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 357914 250954
rect 357294 250634 357914 250718
rect 357294 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 357914 250634
rect 357294 244084 357914 250398
rect 361794 704838 362414 711590
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 244084 362414 254898
rect 366294 705798 366914 711590
rect 366294 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 366914 705798
rect 366294 705478 366914 705562
rect 366294 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 366914 705478
rect 366294 691954 366914 705242
rect 366294 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 366914 691954
rect 366294 691634 366914 691718
rect 366294 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 366914 691634
rect 366294 655954 366914 691398
rect 366294 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 366914 655954
rect 366294 655634 366914 655718
rect 366294 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 366914 655634
rect 366294 619954 366914 655398
rect 366294 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 366914 619954
rect 366294 619634 366914 619718
rect 366294 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 366914 619634
rect 366294 583954 366914 619398
rect 366294 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 366914 583954
rect 366294 583634 366914 583718
rect 366294 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 366914 583634
rect 366294 547954 366914 583398
rect 366294 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 366914 547954
rect 366294 547634 366914 547718
rect 366294 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 366914 547634
rect 366294 511954 366914 547398
rect 366294 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 366914 511954
rect 366294 511634 366914 511718
rect 366294 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 366914 511634
rect 366294 475954 366914 511398
rect 366294 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 366914 475954
rect 366294 475634 366914 475718
rect 366294 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 366914 475634
rect 366294 439954 366914 475398
rect 366294 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 366914 439954
rect 366294 439634 366914 439718
rect 366294 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 366914 439634
rect 366294 403954 366914 439398
rect 366294 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 366914 403954
rect 366294 403634 366914 403718
rect 366294 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 366914 403634
rect 366294 367954 366914 403398
rect 366294 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 366914 367954
rect 366294 367634 366914 367718
rect 366294 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 366914 367634
rect 366294 331954 366914 367398
rect 366294 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 366914 331954
rect 366294 331634 366914 331718
rect 366294 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 366914 331634
rect 366294 295954 366914 331398
rect 366294 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 366914 295954
rect 366294 295634 366914 295718
rect 366294 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 366914 295634
rect 366294 259954 366914 295398
rect 366294 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 366914 259954
rect 366294 259634 366914 259718
rect 366294 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 366914 259634
rect 366294 244084 366914 259398
rect 370794 706758 371414 711590
rect 370794 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 371414 706758
rect 370794 706438 371414 706522
rect 370794 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 371414 706438
rect 370794 696454 371414 706202
rect 370794 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 371414 696454
rect 370794 696134 371414 696218
rect 370794 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 371414 696134
rect 370794 660454 371414 695898
rect 370794 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 371414 660454
rect 370794 660134 371414 660218
rect 370794 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 371414 660134
rect 370794 624454 371414 659898
rect 370794 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 371414 624454
rect 370794 624134 371414 624218
rect 370794 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 371414 624134
rect 370794 588454 371414 623898
rect 370794 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 371414 588454
rect 370794 588134 371414 588218
rect 370794 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 371414 588134
rect 370794 552454 371414 587898
rect 370794 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 371414 552454
rect 370794 552134 371414 552218
rect 370794 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 371414 552134
rect 370794 516454 371414 551898
rect 370794 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 371414 516454
rect 370794 516134 371414 516218
rect 370794 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 371414 516134
rect 370794 480454 371414 515898
rect 370794 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 371414 480454
rect 370794 480134 371414 480218
rect 370794 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 371414 480134
rect 370794 444454 371414 479898
rect 370794 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 371414 444454
rect 370794 444134 371414 444218
rect 370794 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 371414 444134
rect 370794 408454 371414 443898
rect 370794 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 371414 408454
rect 370794 408134 371414 408218
rect 370794 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 371414 408134
rect 370794 372454 371414 407898
rect 370794 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 371414 372454
rect 370794 372134 371414 372218
rect 370794 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 371414 372134
rect 370794 336454 371414 371898
rect 370794 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 371414 336454
rect 370794 336134 371414 336218
rect 370794 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 371414 336134
rect 370794 300454 371414 335898
rect 370794 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 371414 300454
rect 370794 300134 371414 300218
rect 370794 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 371414 300134
rect 370794 264454 371414 299898
rect 370794 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 371414 264454
rect 370794 264134 371414 264218
rect 370794 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 371414 264134
rect 370794 244084 371414 263898
rect 375294 707718 375914 711590
rect 375294 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 375914 707718
rect 375294 707398 375914 707482
rect 375294 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 375914 707398
rect 375294 700954 375914 707162
rect 375294 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 375914 700954
rect 375294 700634 375914 700718
rect 375294 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 375914 700634
rect 375294 664954 375914 700398
rect 375294 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 375914 664954
rect 375294 664634 375914 664718
rect 375294 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 375914 664634
rect 375294 628954 375914 664398
rect 375294 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 375914 628954
rect 375294 628634 375914 628718
rect 375294 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 375914 628634
rect 375294 592954 375914 628398
rect 375294 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 375914 592954
rect 375294 592634 375914 592718
rect 375294 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 375914 592634
rect 375294 556954 375914 592398
rect 375294 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 375914 556954
rect 375294 556634 375914 556718
rect 375294 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 375914 556634
rect 375294 520954 375914 556398
rect 375294 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 375914 520954
rect 375294 520634 375914 520718
rect 375294 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 375914 520634
rect 375294 484954 375914 520398
rect 375294 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 375914 484954
rect 375294 484634 375914 484718
rect 375294 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 375914 484634
rect 375294 448954 375914 484398
rect 375294 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 375914 448954
rect 375294 448634 375914 448718
rect 375294 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 375914 448634
rect 375294 412954 375914 448398
rect 375294 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 375914 412954
rect 375294 412634 375914 412718
rect 375294 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 375914 412634
rect 375294 376954 375914 412398
rect 375294 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 375914 376954
rect 375294 376634 375914 376718
rect 375294 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 375914 376634
rect 375294 340954 375914 376398
rect 375294 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 375914 340954
rect 375294 340634 375914 340718
rect 375294 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 375914 340634
rect 375294 304954 375914 340398
rect 375294 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 375914 304954
rect 375294 304634 375914 304718
rect 375294 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 375914 304634
rect 375294 268954 375914 304398
rect 375294 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 375914 268954
rect 375294 268634 375914 268718
rect 375294 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 375914 268634
rect 375294 244084 375914 268398
rect 379794 708678 380414 711590
rect 379794 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 380414 708678
rect 379794 708358 380414 708442
rect 379794 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 380414 708358
rect 379794 669454 380414 708122
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 244084 380414 272898
rect 384294 709638 384914 711590
rect 384294 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 384914 709638
rect 384294 709318 384914 709402
rect 384294 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 384914 709318
rect 384294 673954 384914 709082
rect 384294 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 384914 673954
rect 384294 673634 384914 673718
rect 384294 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 384914 673634
rect 384294 637954 384914 673398
rect 384294 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 384914 637954
rect 384294 637634 384914 637718
rect 384294 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 384914 637634
rect 384294 601954 384914 637398
rect 384294 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 384914 601954
rect 384294 601634 384914 601718
rect 384294 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 384914 601634
rect 384294 565954 384914 601398
rect 384294 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 384914 565954
rect 384294 565634 384914 565718
rect 384294 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 384914 565634
rect 384294 529954 384914 565398
rect 384294 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 384914 529954
rect 384294 529634 384914 529718
rect 384294 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 384914 529634
rect 384294 493954 384914 529398
rect 384294 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 384914 493954
rect 384294 493634 384914 493718
rect 384294 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 384914 493634
rect 384294 457954 384914 493398
rect 384294 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 384914 457954
rect 384294 457634 384914 457718
rect 384294 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 384914 457634
rect 384294 421954 384914 457398
rect 384294 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 384914 421954
rect 384294 421634 384914 421718
rect 384294 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 384914 421634
rect 384294 385954 384914 421398
rect 384294 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 384914 385954
rect 384294 385634 384914 385718
rect 384294 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 384914 385634
rect 384294 349954 384914 385398
rect 384294 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 384914 349954
rect 384294 349634 384914 349718
rect 384294 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 384914 349634
rect 384294 313954 384914 349398
rect 384294 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 384914 313954
rect 384294 313634 384914 313718
rect 384294 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 384914 313634
rect 384294 277954 384914 313398
rect 384294 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 384914 277954
rect 384294 277634 384914 277718
rect 384294 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 384914 277634
rect 384294 244084 384914 277398
rect 388794 710598 389414 711590
rect 388794 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 389414 710598
rect 388794 710278 389414 710362
rect 388794 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 389414 710278
rect 388794 678454 389414 710042
rect 388794 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 389414 678454
rect 388794 678134 389414 678218
rect 388794 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 389414 678134
rect 388794 642454 389414 677898
rect 388794 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 389414 642454
rect 388794 642134 389414 642218
rect 388794 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 389414 642134
rect 388794 606454 389414 641898
rect 388794 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 389414 606454
rect 388794 606134 389414 606218
rect 388794 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 389414 606134
rect 388794 570454 389414 605898
rect 388794 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 389414 570454
rect 388794 570134 389414 570218
rect 388794 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 389414 570134
rect 388794 534454 389414 569898
rect 388794 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 389414 534454
rect 388794 534134 389414 534218
rect 388794 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 389414 534134
rect 388794 498454 389414 533898
rect 388794 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 389414 498454
rect 388794 498134 389414 498218
rect 388794 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 389414 498134
rect 388794 462454 389414 497898
rect 388794 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 389414 462454
rect 388794 462134 389414 462218
rect 388794 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 389414 462134
rect 388794 426454 389414 461898
rect 388794 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 389414 426454
rect 388794 426134 389414 426218
rect 388794 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 389414 426134
rect 388794 390454 389414 425898
rect 388794 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 389414 390454
rect 388794 390134 389414 390218
rect 388794 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 389414 390134
rect 388794 354454 389414 389898
rect 388794 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 389414 354454
rect 388794 354134 389414 354218
rect 388794 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 389414 354134
rect 388794 318454 389414 353898
rect 388794 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 389414 318454
rect 388794 318134 389414 318218
rect 388794 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 389414 318134
rect 388794 282454 389414 317898
rect 388794 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 389414 282454
rect 388794 282134 389414 282218
rect 388794 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 389414 282134
rect 388794 246454 389414 281898
rect 388794 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 389414 246454
rect 388794 246134 389414 246218
rect 388794 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 389414 246134
rect 388794 244084 389414 245898
rect 393294 711558 393914 711590
rect 393294 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 393914 711558
rect 393294 711238 393914 711322
rect 393294 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 393914 711238
rect 393294 682954 393914 711002
rect 393294 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 393914 682954
rect 393294 682634 393914 682718
rect 393294 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 393914 682634
rect 393294 646954 393914 682398
rect 393294 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 393914 646954
rect 393294 646634 393914 646718
rect 393294 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 393914 646634
rect 393294 610954 393914 646398
rect 393294 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 393914 610954
rect 393294 610634 393914 610718
rect 393294 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 393914 610634
rect 393294 574954 393914 610398
rect 393294 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 393914 574954
rect 393294 574634 393914 574718
rect 393294 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 393914 574634
rect 393294 538954 393914 574398
rect 393294 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 393914 538954
rect 393294 538634 393914 538718
rect 393294 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 393914 538634
rect 393294 502954 393914 538398
rect 393294 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 393914 502954
rect 393294 502634 393914 502718
rect 393294 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 393914 502634
rect 393294 466954 393914 502398
rect 393294 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 393914 466954
rect 393294 466634 393914 466718
rect 393294 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 393914 466634
rect 393294 430954 393914 466398
rect 393294 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 393914 430954
rect 393294 430634 393914 430718
rect 393294 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 393914 430634
rect 393294 394954 393914 430398
rect 393294 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 393914 394954
rect 393294 394634 393914 394718
rect 393294 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 393914 394634
rect 393294 358954 393914 394398
rect 393294 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 393914 358954
rect 393294 358634 393914 358718
rect 393294 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 393914 358634
rect 393294 322954 393914 358398
rect 393294 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 393914 322954
rect 393294 322634 393914 322718
rect 393294 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 393914 322634
rect 393294 286954 393914 322398
rect 393294 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 393914 286954
rect 393294 286634 393914 286718
rect 393294 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 393914 286634
rect 393294 250954 393914 286398
rect 393294 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 393914 250954
rect 393294 250634 393914 250718
rect 393294 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 393914 250634
rect 393294 244084 393914 250398
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 244084 398414 254898
rect 402294 705798 402914 711590
rect 402294 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 402914 705798
rect 402294 705478 402914 705562
rect 402294 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 402914 705478
rect 402294 691954 402914 705242
rect 402294 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 402914 691954
rect 402294 691634 402914 691718
rect 402294 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 402914 691634
rect 402294 655954 402914 691398
rect 402294 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 402914 655954
rect 402294 655634 402914 655718
rect 402294 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 402914 655634
rect 402294 619954 402914 655398
rect 402294 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 402914 619954
rect 402294 619634 402914 619718
rect 402294 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 402914 619634
rect 402294 583954 402914 619398
rect 402294 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 402914 583954
rect 402294 583634 402914 583718
rect 402294 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 402914 583634
rect 402294 547954 402914 583398
rect 402294 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 402914 547954
rect 402294 547634 402914 547718
rect 402294 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 402914 547634
rect 402294 511954 402914 547398
rect 402294 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 402914 511954
rect 402294 511634 402914 511718
rect 402294 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 402914 511634
rect 402294 475954 402914 511398
rect 402294 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 402914 475954
rect 402294 475634 402914 475718
rect 402294 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 402914 475634
rect 402294 439954 402914 475398
rect 402294 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 402914 439954
rect 402294 439634 402914 439718
rect 402294 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 402914 439634
rect 402294 403954 402914 439398
rect 402294 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 402914 403954
rect 402294 403634 402914 403718
rect 402294 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 402914 403634
rect 402294 367954 402914 403398
rect 402294 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 402914 367954
rect 402294 367634 402914 367718
rect 402294 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 402914 367634
rect 402294 331954 402914 367398
rect 402294 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 402914 331954
rect 402294 331634 402914 331718
rect 402294 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 402914 331634
rect 402294 295954 402914 331398
rect 402294 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 402914 295954
rect 402294 295634 402914 295718
rect 402294 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 402914 295634
rect 402294 259954 402914 295398
rect 402294 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 402914 259954
rect 402294 259634 402914 259718
rect 402294 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 402914 259634
rect 402294 244084 402914 259398
rect 406794 706758 407414 711590
rect 406794 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 407414 706758
rect 406794 706438 407414 706522
rect 406794 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 407414 706438
rect 406794 696454 407414 706202
rect 406794 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 407414 696454
rect 406794 696134 407414 696218
rect 406794 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 407414 696134
rect 406794 660454 407414 695898
rect 406794 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 407414 660454
rect 406794 660134 407414 660218
rect 406794 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 407414 660134
rect 406794 624454 407414 659898
rect 406794 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 407414 624454
rect 406794 624134 407414 624218
rect 406794 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 407414 624134
rect 406794 588454 407414 623898
rect 406794 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 407414 588454
rect 406794 588134 407414 588218
rect 406794 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 407414 588134
rect 406794 552454 407414 587898
rect 406794 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 407414 552454
rect 406794 552134 407414 552218
rect 406794 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 407414 552134
rect 406794 516454 407414 551898
rect 406794 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 407414 516454
rect 406794 516134 407414 516218
rect 406794 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 407414 516134
rect 406794 480454 407414 515898
rect 406794 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 407414 480454
rect 406794 480134 407414 480218
rect 406794 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 407414 480134
rect 406794 444454 407414 479898
rect 406794 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 407414 444454
rect 406794 444134 407414 444218
rect 406794 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 407414 444134
rect 406794 408454 407414 443898
rect 406794 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 407414 408454
rect 406794 408134 407414 408218
rect 406794 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 407414 408134
rect 406794 372454 407414 407898
rect 406794 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 407414 372454
rect 406794 372134 407414 372218
rect 406794 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 407414 372134
rect 406794 336454 407414 371898
rect 406794 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 407414 336454
rect 406794 336134 407414 336218
rect 406794 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 407414 336134
rect 406794 300454 407414 335898
rect 406794 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 407414 300454
rect 406794 300134 407414 300218
rect 406794 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 407414 300134
rect 406794 264454 407414 299898
rect 406794 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 407414 264454
rect 406794 264134 407414 264218
rect 406794 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 407414 264134
rect 71300 241953 77300 241984
rect 71300 241717 71462 241953
rect 71698 241717 71782 241953
rect 72018 241717 72102 241953
rect 72338 241717 72422 241953
rect 72658 241717 72742 241953
rect 72978 241717 73062 241953
rect 73298 241717 73382 241953
rect 73618 241717 73702 241953
rect 73938 241717 74022 241953
rect 74258 241717 74342 241953
rect 74578 241717 74662 241953
rect 74898 241717 74982 241953
rect 75218 241717 75302 241953
rect 75538 241717 75622 241953
rect 75858 241717 75942 241953
rect 76178 241717 76262 241953
rect 76498 241717 76582 241953
rect 76818 241717 76902 241953
rect 77138 241717 77300 241953
rect 71300 241633 77300 241717
rect 71300 241397 71462 241633
rect 71698 241397 71782 241633
rect 72018 241397 72102 241633
rect 72338 241397 72422 241633
rect 72658 241397 72742 241633
rect 72978 241397 73062 241633
rect 73298 241397 73382 241633
rect 73618 241397 73702 241633
rect 73938 241397 74022 241633
rect 74258 241397 74342 241633
rect 74578 241397 74662 241633
rect 74898 241397 74982 241633
rect 75218 241397 75302 241633
rect 75538 241397 75622 241633
rect 75858 241397 75942 241633
rect 76178 241397 76262 241633
rect 76498 241397 76582 241633
rect 76818 241397 76902 241633
rect 77138 241397 77300 241633
rect 71300 241366 77300 241397
rect 46000 237453 50794 237484
rect 46000 237217 46039 237453
rect 46275 237217 46359 237453
rect 46595 237217 46679 237453
rect 46915 237217 46999 237453
rect 47235 237217 47319 237453
rect 47555 237217 47639 237453
rect 47875 237217 47959 237453
rect 48195 237217 48279 237453
rect 48515 237217 48599 237453
rect 48835 237217 48919 237453
rect 49155 237217 49239 237453
rect 49475 237217 49559 237453
rect 49795 237217 49879 237453
rect 50115 237217 50199 237453
rect 50435 237217 50519 237453
rect 50755 237217 50794 237453
rect 46000 237133 50794 237217
rect 46000 236897 46039 237133
rect 46275 236897 46359 237133
rect 46595 236897 46679 237133
rect 46915 236897 46999 237133
rect 47235 236897 47319 237133
rect 47555 236897 47639 237133
rect 47875 236897 47959 237133
rect 48195 236897 48279 237133
rect 48515 236897 48599 237133
rect 48835 236897 48919 237133
rect 49155 236897 49239 237133
rect 49475 236897 49559 237133
rect 49795 236897 49879 237133
rect 50115 236897 50199 237133
rect 50435 236897 50519 237133
rect 50755 236897 50794 237133
rect 46000 236866 50794 236897
rect 42294 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 42914 223954
rect 42294 223634 42914 223718
rect 42294 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 42914 223634
rect 42294 187954 42914 223398
rect 42294 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 42914 187954
rect 42294 187634 42914 187718
rect 42294 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 42914 187634
rect 42294 151954 42914 187398
rect 42294 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 42914 151954
rect 42294 151634 42914 151718
rect 42294 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 42914 151634
rect 42294 115954 42914 151398
rect 42294 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 42914 115954
rect 42294 115634 42914 115718
rect 42294 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 42914 115634
rect 42294 79954 42914 115398
rect 42294 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 42914 79954
rect 42294 79634 42914 79718
rect 42294 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 42914 79634
rect 42294 43954 42914 79398
rect 42294 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 42914 43954
rect 42294 43634 42914 43718
rect 42294 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 42914 43634
rect 42294 7954 42914 43398
rect 42294 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 42914 7954
rect 42294 7634 42914 7718
rect 42294 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 42914 7634
rect 42294 -1306 42914 7398
rect 42294 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 42914 -1306
rect 42294 -1626 42914 -1542
rect 42294 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 42914 -1626
rect 42294 -7654 42914 -1862
rect 46794 228453 47414 228484
rect 46794 228217 46826 228453
rect 47062 228217 47146 228453
rect 47382 228217 47414 228453
rect 46794 228133 47414 228217
rect 46794 227897 46826 228133
rect 47062 227897 47146 228133
rect 47382 227897 47414 228133
rect 46794 192454 47414 227897
rect 46794 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 47414 192454
rect 46794 192134 47414 192218
rect 46794 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 47414 192134
rect 46794 156454 47414 191898
rect 46794 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 47414 156454
rect 46794 156134 47414 156218
rect 46794 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 47414 156134
rect 46794 120454 47414 155898
rect 46794 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 47414 120454
rect 46794 120134 47414 120218
rect 46794 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 47414 120134
rect 46794 84454 47414 119898
rect 46794 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 47414 84454
rect 46794 84134 47414 84218
rect 46794 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 47414 84134
rect 46794 48454 47414 83898
rect 46794 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 47414 48454
rect 46794 48134 47414 48218
rect 46794 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 47414 48134
rect 46794 12454 47414 47898
rect 46794 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 47414 12454
rect 46794 12134 47414 12218
rect 46794 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 47414 12134
rect 46794 -2266 47414 11898
rect 46794 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 47414 -2266
rect 46794 -2586 47414 -2502
rect 46794 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 47414 -2586
rect 46794 -7654 47414 -2822
rect 51294 196954 51914 228484
rect 51294 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 51914 196954
rect 51294 196634 51914 196718
rect 51294 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 51914 196634
rect 51294 160954 51914 196398
rect 51294 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 51914 160954
rect 51294 160634 51914 160718
rect 51294 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 51914 160634
rect 51294 124954 51914 160398
rect 51294 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 51914 124954
rect 51294 124634 51914 124718
rect 51294 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 51914 124634
rect 51294 88954 51914 124398
rect 51294 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 51914 88954
rect 51294 88634 51914 88718
rect 51294 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 51914 88634
rect 51294 52954 51914 88398
rect 51294 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 51914 52954
rect 51294 52634 51914 52718
rect 51294 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 51914 52634
rect 51294 16954 51914 52398
rect 51294 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 51914 16954
rect 51294 16634 51914 16718
rect 51294 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 51914 16634
rect 51294 -3226 51914 16398
rect 51294 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 51914 -3226
rect 51294 -3546 51914 -3462
rect 51294 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 51914 -3546
rect 51294 -7654 51914 -3782
rect 55794 201454 56414 228484
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -4186 56414 20898
rect 55794 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 56414 -4186
rect 55794 -4506 56414 -4422
rect 55794 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 56414 -4506
rect 55794 -7654 56414 -4742
rect 60294 205954 60914 228484
rect 60294 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 60914 205954
rect 60294 205634 60914 205718
rect 60294 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 60914 205634
rect 60294 169954 60914 205398
rect 60294 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 60914 169954
rect 60294 169634 60914 169718
rect 60294 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 60914 169634
rect 60294 133954 60914 169398
rect 60294 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 60914 133954
rect 60294 133634 60914 133718
rect 60294 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 60914 133634
rect 60294 97954 60914 133398
rect 60294 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 60914 97954
rect 60294 97634 60914 97718
rect 60294 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 60914 97634
rect 60294 61954 60914 97398
rect 60294 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 60914 61954
rect 60294 61634 60914 61718
rect 60294 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 60914 61634
rect 60294 25954 60914 61398
rect 60294 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 60914 25954
rect 60294 25634 60914 25718
rect 60294 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 60914 25634
rect 60294 -5146 60914 25398
rect 60294 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 60914 -5146
rect 60294 -5466 60914 -5382
rect 60294 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 60914 -5466
rect 60294 -7654 60914 -5702
rect 64794 210454 65414 228484
rect 64794 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 65414 210454
rect 64794 210134 65414 210218
rect 64794 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 65414 210134
rect 64794 174454 65414 209898
rect 64794 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 65414 174454
rect 64794 174134 65414 174218
rect 64794 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 65414 174134
rect 64794 138454 65414 173898
rect 64794 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 65414 138454
rect 64794 138134 65414 138218
rect 64794 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 65414 138134
rect 64794 102454 65414 137898
rect 64794 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 65414 102454
rect 64794 102134 65414 102218
rect 64794 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 65414 102134
rect 64794 66454 65414 101898
rect 64794 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 65414 66454
rect 64794 66134 65414 66218
rect 64794 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 65414 66134
rect 64794 30454 65414 65898
rect 64794 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 65414 30454
rect 64794 30134 65414 30218
rect 64794 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 65414 30134
rect 64794 -6106 65414 29898
rect 64794 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 65414 -6106
rect 64794 -6426 65414 -6342
rect 64794 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 65414 -6426
rect 64794 -7654 65414 -6662
rect 69294 214954 69914 228484
rect 69294 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 69914 214954
rect 69294 214634 69914 214718
rect 69294 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 69914 214634
rect 69294 178954 69914 214398
rect 69294 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 69914 178954
rect 69294 178634 69914 178718
rect 69294 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 69914 178634
rect 69294 142954 69914 178398
rect 69294 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 69914 142954
rect 69294 142634 69914 142718
rect 69294 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 69914 142634
rect 69294 106954 69914 142398
rect 69294 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 69914 106954
rect 69294 106634 69914 106718
rect 69294 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 69914 106634
rect 69294 70954 69914 106398
rect 69294 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 69914 70954
rect 69294 70634 69914 70718
rect 69294 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 69914 70634
rect 69294 34954 69914 70398
rect 69294 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 69914 34954
rect 69294 34634 69914 34718
rect 69294 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 69914 34634
rect 69294 -7066 69914 34398
rect 69294 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 69914 -7066
rect 69294 -7386 69914 -7302
rect 69294 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 69914 -7386
rect 69294 -7654 69914 -7622
rect 73794 219454 74414 228484
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 78294 223954 78914 228484
rect 78294 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 78914 223954
rect 78294 223634 78914 223718
rect 78294 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 78914 223634
rect 78294 187954 78914 223398
rect 78294 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 78914 187954
rect 78294 187634 78914 187718
rect 78294 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 78914 187634
rect 78294 151954 78914 187398
rect 78294 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 78914 151954
rect 78294 151634 78914 151718
rect 78294 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 78914 151634
rect 78294 115954 78914 151398
rect 78294 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 78914 115954
rect 78294 115634 78914 115718
rect 78294 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 78914 115634
rect 78294 79954 78914 115398
rect 78294 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 78914 79954
rect 78294 79634 78914 79718
rect 78294 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 78914 79634
rect 78294 43954 78914 79398
rect 78294 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 78914 43954
rect 78294 43634 78914 43718
rect 78294 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 78914 43634
rect 78294 7954 78914 43398
rect 78294 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 78914 7954
rect 78294 7634 78914 7718
rect 78294 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 78914 7634
rect 78294 -1306 78914 7398
rect 78294 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 78914 -1306
rect 78294 -1626 78914 -1542
rect 78294 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 78914 -1626
rect 78294 -7654 78914 -1862
rect 82794 228453 83414 228484
rect 82794 228217 82826 228453
rect 83062 228217 83146 228453
rect 83382 228217 83414 228453
rect 82794 228133 83414 228217
rect 82794 227897 82826 228133
rect 83062 227897 83146 228133
rect 83382 227897 83414 228133
rect 82794 192454 83414 227897
rect 82794 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 83414 192454
rect 82794 192134 83414 192218
rect 82794 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 83414 192134
rect 82794 156454 83414 191898
rect 82794 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 83414 156454
rect 82794 156134 83414 156218
rect 82794 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 83414 156134
rect 82794 120454 83414 155898
rect 82794 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 83414 120454
rect 82794 120134 83414 120218
rect 82794 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 83414 120134
rect 82794 84454 83414 119898
rect 82794 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 83414 84454
rect 82794 84134 83414 84218
rect 82794 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 83414 84134
rect 82794 48454 83414 83898
rect 82794 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 83414 48454
rect 82794 48134 83414 48218
rect 82794 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 83414 48134
rect 82794 12454 83414 47898
rect 82794 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 83414 12454
rect 82794 12134 83414 12218
rect 82794 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 83414 12134
rect 82794 -2266 83414 11898
rect 82794 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 83414 -2266
rect 82794 -2586 83414 -2502
rect 82794 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 83414 -2586
rect 82794 -7654 83414 -2822
rect 87294 196954 87914 228484
rect 87294 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 87914 196954
rect 87294 196634 87914 196718
rect 87294 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 87914 196634
rect 87294 160954 87914 196398
rect 87294 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 87914 160954
rect 87294 160634 87914 160718
rect 87294 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 87914 160634
rect 87294 124954 87914 160398
rect 87294 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 87914 124954
rect 87294 124634 87914 124718
rect 87294 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 87914 124634
rect 87294 88954 87914 124398
rect 87294 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 87914 88954
rect 87294 88634 87914 88718
rect 87294 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 87914 88634
rect 87294 52954 87914 88398
rect 87294 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 87914 52954
rect 87294 52634 87914 52718
rect 87294 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 87914 52634
rect 87294 16954 87914 52398
rect 87294 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 87914 16954
rect 87294 16634 87914 16718
rect 87294 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 87914 16634
rect 87294 -3226 87914 16398
rect 87294 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 87914 -3226
rect 87294 -3546 87914 -3462
rect 87294 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 87914 -3546
rect 87294 -7654 87914 -3782
rect 91794 201454 92414 228484
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 129454 92414 164898
rect 91794 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 92414 129454
rect 91794 129134 92414 129218
rect 91794 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 92414 129134
rect 91794 93454 92414 128898
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 91794 57454 92414 92898
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -4186 92414 20898
rect 91794 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 92414 -4186
rect 91794 -4506 92414 -4422
rect 91794 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 92414 -4506
rect 91794 -7654 92414 -4742
rect 96294 205954 96914 228484
rect 96294 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 96914 205954
rect 96294 205634 96914 205718
rect 96294 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 96914 205634
rect 96294 169954 96914 205398
rect 96294 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 96914 169954
rect 96294 169634 96914 169718
rect 96294 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 96914 169634
rect 96294 133954 96914 169398
rect 96294 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 96914 133954
rect 96294 133634 96914 133718
rect 96294 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 96914 133634
rect 96294 97954 96914 133398
rect 96294 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 96914 97954
rect 96294 97634 96914 97718
rect 96294 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 96914 97634
rect 96294 61954 96914 97398
rect 96294 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 96914 61954
rect 96294 61634 96914 61718
rect 96294 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 96914 61634
rect 96294 25954 96914 61398
rect 96294 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 96914 25954
rect 96294 25634 96914 25718
rect 96294 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 96914 25634
rect 96294 -5146 96914 25398
rect 96294 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 96914 -5146
rect 96294 -5466 96914 -5382
rect 96294 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 96914 -5466
rect 96294 -7654 96914 -5702
rect 100794 210454 101414 228484
rect 100794 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 101414 210454
rect 100794 210134 101414 210218
rect 100794 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 101414 210134
rect 100794 174454 101414 209898
rect 100794 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 101414 174454
rect 100794 174134 101414 174218
rect 100794 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 101414 174134
rect 100794 138454 101414 173898
rect 100794 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 101414 138454
rect 100794 138134 101414 138218
rect 100794 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 101414 138134
rect 100794 102454 101414 137898
rect 100794 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 101414 102454
rect 100794 102134 101414 102218
rect 100794 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 101414 102134
rect 100794 66454 101414 101898
rect 100794 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 101414 66454
rect 100794 66134 101414 66218
rect 100794 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 101414 66134
rect 100794 30454 101414 65898
rect 100794 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 101414 30454
rect 100794 30134 101414 30218
rect 100794 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 101414 30134
rect 100794 -6106 101414 29898
rect 100794 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 101414 -6106
rect 100794 -6426 101414 -6342
rect 100794 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 101414 -6426
rect 100794 -7654 101414 -6662
rect 105294 214954 105914 228484
rect 105294 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 105914 214954
rect 105294 214634 105914 214718
rect 105294 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 105914 214634
rect 105294 178954 105914 214398
rect 105294 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 105914 178954
rect 105294 178634 105914 178718
rect 105294 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 105914 178634
rect 105294 142954 105914 178398
rect 105294 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 105914 142954
rect 105294 142634 105914 142718
rect 105294 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 105914 142634
rect 105294 106954 105914 142398
rect 105294 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 105914 106954
rect 105294 106634 105914 106718
rect 105294 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 105914 106634
rect 105294 70954 105914 106398
rect 105294 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 105914 70954
rect 105294 70634 105914 70718
rect 105294 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 105914 70634
rect 105294 34954 105914 70398
rect 105294 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 105914 34954
rect 105294 34634 105914 34718
rect 105294 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 105914 34634
rect 105294 -7066 105914 34398
rect 105294 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 105914 -7066
rect 105294 -7386 105914 -7302
rect 105294 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 105914 -7386
rect 105294 -7654 105914 -7622
rect 109794 219454 110414 228484
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 114294 223954 114914 228484
rect 114294 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 114914 223954
rect 114294 223634 114914 223718
rect 114294 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 114914 223634
rect 114294 187954 114914 223398
rect 114294 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 114914 187954
rect 114294 187634 114914 187718
rect 114294 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 114914 187634
rect 114294 151954 114914 187398
rect 114294 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 114914 151954
rect 114294 151634 114914 151718
rect 114294 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 114914 151634
rect 114294 115954 114914 151398
rect 118794 228453 119414 228484
rect 118794 228217 118826 228453
rect 119062 228217 119146 228453
rect 119382 228217 119414 228453
rect 118794 228133 119414 228217
rect 118794 227897 118826 228133
rect 119062 227897 119146 228133
rect 119382 227897 119414 228133
rect 118794 192454 119414 227897
rect 118794 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 119414 192454
rect 118794 192134 119414 192218
rect 118794 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 119414 192134
rect 118794 156454 119414 191898
rect 118794 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 119414 156454
rect 118794 156134 119414 156218
rect 118794 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 119414 156134
rect 118794 142000 119414 155898
rect 123294 196954 123914 228484
rect 123294 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 123914 196954
rect 123294 196634 123914 196718
rect 123294 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 123914 196634
rect 123294 160954 123914 196398
rect 123294 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 123914 160954
rect 123294 160634 123914 160718
rect 123294 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 123914 160634
rect 123294 142000 123914 160398
rect 127794 201454 128414 228484
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 127794 165454 128414 200898
rect 127794 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 128414 165454
rect 127794 165134 128414 165218
rect 127794 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 128414 165134
rect 127794 142000 128414 164898
rect 132294 205954 132914 228484
rect 132294 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205718 132914 205954
rect 132294 205634 132914 205718
rect 132294 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205398 132914 205634
rect 132294 169954 132914 205398
rect 135914 205954 165514 205986
rect 135914 205718 136036 205954
rect 136272 205718 136356 205954
rect 136592 205718 136676 205954
rect 136912 205718 136996 205954
rect 137232 205718 137316 205954
rect 137552 205718 137636 205954
rect 137872 205718 137956 205954
rect 138192 205718 138276 205954
rect 138512 205718 138596 205954
rect 138832 205718 138916 205954
rect 139152 205718 139236 205954
rect 139472 205718 139556 205954
rect 139792 205718 139876 205954
rect 140112 205718 140196 205954
rect 140432 205718 140516 205954
rect 140752 205718 140836 205954
rect 141072 205718 141156 205954
rect 141392 205718 141476 205954
rect 141712 205718 141796 205954
rect 142032 205718 142116 205954
rect 142352 205718 142436 205954
rect 142672 205718 142756 205954
rect 142992 205718 143076 205954
rect 143312 205718 143396 205954
rect 143632 205718 143716 205954
rect 143952 205718 144036 205954
rect 144272 205718 144356 205954
rect 144592 205718 144676 205954
rect 144912 205718 144996 205954
rect 145232 205718 145316 205954
rect 145552 205718 145636 205954
rect 145872 205718 145956 205954
rect 146192 205718 146276 205954
rect 146512 205718 146596 205954
rect 146832 205718 146916 205954
rect 147152 205718 147236 205954
rect 147472 205718 147556 205954
rect 147792 205718 147876 205954
rect 148112 205718 148196 205954
rect 148432 205718 148516 205954
rect 148752 205718 148836 205954
rect 149072 205718 149156 205954
rect 149392 205718 149476 205954
rect 149712 205718 149796 205954
rect 150032 205718 150116 205954
rect 150352 205718 150436 205954
rect 150672 205718 150756 205954
rect 150992 205718 151076 205954
rect 151312 205718 151396 205954
rect 151632 205718 151716 205954
rect 151952 205718 152036 205954
rect 152272 205718 152356 205954
rect 152592 205718 152676 205954
rect 152912 205718 152996 205954
rect 153232 205718 153316 205954
rect 153552 205718 153636 205954
rect 153872 205718 153956 205954
rect 154192 205718 154276 205954
rect 154512 205718 154596 205954
rect 154832 205718 154916 205954
rect 155152 205718 155236 205954
rect 155472 205718 155556 205954
rect 155792 205718 155876 205954
rect 156112 205718 156196 205954
rect 156432 205718 156516 205954
rect 156752 205718 156836 205954
rect 157072 205718 157156 205954
rect 157392 205718 157476 205954
rect 157712 205718 157796 205954
rect 158032 205718 158116 205954
rect 158352 205718 158436 205954
rect 158672 205718 158756 205954
rect 158992 205718 159076 205954
rect 159312 205718 159396 205954
rect 159632 205718 159716 205954
rect 159952 205718 160036 205954
rect 160272 205718 160356 205954
rect 160592 205718 160676 205954
rect 160912 205718 160996 205954
rect 161232 205718 161316 205954
rect 161552 205718 161636 205954
rect 161872 205718 161956 205954
rect 162192 205718 162276 205954
rect 162512 205718 162596 205954
rect 162832 205718 162916 205954
rect 163152 205718 163236 205954
rect 163472 205718 163556 205954
rect 163792 205718 163876 205954
rect 164112 205718 164196 205954
rect 164432 205718 164516 205954
rect 164752 205718 164836 205954
rect 165072 205718 165156 205954
rect 165392 205718 165514 205954
rect 135914 205634 165514 205718
rect 135914 205398 136036 205634
rect 136272 205398 136356 205634
rect 136592 205398 136676 205634
rect 136912 205398 136996 205634
rect 137232 205398 137316 205634
rect 137552 205398 137636 205634
rect 137872 205398 137956 205634
rect 138192 205398 138276 205634
rect 138512 205398 138596 205634
rect 138832 205398 138916 205634
rect 139152 205398 139236 205634
rect 139472 205398 139556 205634
rect 139792 205398 139876 205634
rect 140112 205398 140196 205634
rect 140432 205398 140516 205634
rect 140752 205398 140836 205634
rect 141072 205398 141156 205634
rect 141392 205398 141476 205634
rect 141712 205398 141796 205634
rect 142032 205398 142116 205634
rect 142352 205398 142436 205634
rect 142672 205398 142756 205634
rect 142992 205398 143076 205634
rect 143312 205398 143396 205634
rect 143632 205398 143716 205634
rect 143952 205398 144036 205634
rect 144272 205398 144356 205634
rect 144592 205398 144676 205634
rect 144912 205398 144996 205634
rect 145232 205398 145316 205634
rect 145552 205398 145636 205634
rect 145872 205398 145956 205634
rect 146192 205398 146276 205634
rect 146512 205398 146596 205634
rect 146832 205398 146916 205634
rect 147152 205398 147236 205634
rect 147472 205398 147556 205634
rect 147792 205398 147876 205634
rect 148112 205398 148196 205634
rect 148432 205398 148516 205634
rect 148752 205398 148836 205634
rect 149072 205398 149156 205634
rect 149392 205398 149476 205634
rect 149712 205398 149796 205634
rect 150032 205398 150116 205634
rect 150352 205398 150436 205634
rect 150672 205398 150756 205634
rect 150992 205398 151076 205634
rect 151312 205398 151396 205634
rect 151632 205398 151716 205634
rect 151952 205398 152036 205634
rect 152272 205398 152356 205634
rect 152592 205398 152676 205634
rect 152912 205398 152996 205634
rect 153232 205398 153316 205634
rect 153552 205398 153636 205634
rect 153872 205398 153956 205634
rect 154192 205398 154276 205634
rect 154512 205398 154596 205634
rect 154832 205398 154916 205634
rect 155152 205398 155236 205634
rect 155472 205398 155556 205634
rect 155792 205398 155876 205634
rect 156112 205398 156196 205634
rect 156432 205398 156516 205634
rect 156752 205398 156836 205634
rect 157072 205398 157156 205634
rect 157392 205398 157476 205634
rect 157712 205398 157796 205634
rect 158032 205398 158116 205634
rect 158352 205398 158436 205634
rect 158672 205398 158756 205634
rect 158992 205398 159076 205634
rect 159312 205398 159396 205634
rect 159632 205398 159716 205634
rect 159952 205398 160036 205634
rect 160272 205398 160356 205634
rect 160592 205398 160676 205634
rect 160912 205398 160996 205634
rect 161232 205398 161316 205634
rect 161552 205398 161636 205634
rect 161872 205398 161956 205634
rect 162192 205398 162276 205634
rect 162512 205398 162596 205634
rect 162832 205398 162916 205634
rect 163152 205398 163236 205634
rect 163472 205398 163556 205634
rect 163792 205398 163876 205634
rect 164112 205398 164196 205634
rect 164432 205398 164516 205634
rect 164752 205398 164836 205634
rect 165072 205398 165156 205634
rect 165392 205398 165514 205634
rect 135914 205366 165514 205398
rect 168294 205954 168914 228484
rect 168294 205718 168326 205954
rect 168562 205718 168646 205954
rect 168882 205718 168914 205954
rect 168294 205634 168914 205718
rect 168294 205398 168326 205634
rect 168562 205398 168646 205634
rect 168882 205398 168914 205634
rect 137314 201454 165514 201486
rect 137314 201218 137376 201454
rect 137612 201218 137696 201454
rect 137932 201218 138016 201454
rect 138252 201218 138336 201454
rect 138572 201218 138656 201454
rect 138892 201218 138976 201454
rect 139212 201218 139296 201454
rect 139532 201218 139616 201454
rect 139852 201218 139936 201454
rect 140172 201218 140256 201454
rect 140492 201218 140576 201454
rect 140812 201218 140896 201454
rect 141132 201218 141216 201454
rect 141452 201218 141536 201454
rect 141772 201218 141856 201454
rect 142092 201218 142176 201454
rect 142412 201218 142496 201454
rect 142732 201218 142816 201454
rect 143052 201218 143136 201454
rect 143372 201218 143456 201454
rect 143692 201218 143776 201454
rect 144012 201218 144096 201454
rect 144332 201218 144416 201454
rect 144652 201218 144736 201454
rect 144972 201218 145056 201454
rect 145292 201218 145376 201454
rect 145612 201218 145696 201454
rect 145932 201218 146016 201454
rect 146252 201218 146336 201454
rect 146572 201218 146656 201454
rect 146892 201218 146976 201454
rect 147212 201218 147296 201454
rect 147532 201218 147616 201454
rect 147852 201218 147936 201454
rect 148172 201218 148256 201454
rect 148492 201218 148576 201454
rect 148812 201218 148896 201454
rect 149132 201218 149216 201454
rect 149452 201218 149536 201454
rect 149772 201218 149856 201454
rect 150092 201218 150176 201454
rect 150412 201218 150496 201454
rect 150732 201218 150816 201454
rect 151052 201218 151136 201454
rect 151372 201218 151456 201454
rect 151692 201218 151776 201454
rect 152012 201218 152096 201454
rect 152332 201218 152416 201454
rect 152652 201218 152736 201454
rect 152972 201218 153056 201454
rect 153292 201218 153376 201454
rect 153612 201218 153696 201454
rect 153932 201218 154016 201454
rect 154252 201218 154336 201454
rect 154572 201218 154656 201454
rect 154892 201218 154976 201454
rect 155212 201218 155296 201454
rect 155532 201218 155616 201454
rect 155852 201218 155936 201454
rect 156172 201218 156256 201454
rect 156492 201218 156576 201454
rect 156812 201218 156896 201454
rect 157132 201218 157216 201454
rect 157452 201218 157536 201454
rect 157772 201218 157856 201454
rect 158092 201218 158176 201454
rect 158412 201218 158496 201454
rect 158732 201218 158816 201454
rect 159052 201218 159136 201454
rect 159372 201218 159456 201454
rect 159692 201218 159776 201454
rect 160012 201218 160096 201454
rect 160332 201218 160416 201454
rect 160652 201218 160736 201454
rect 160972 201218 161056 201454
rect 161292 201218 161376 201454
rect 161612 201218 161696 201454
rect 161932 201218 162016 201454
rect 162252 201218 162336 201454
rect 162572 201218 162656 201454
rect 162892 201218 162976 201454
rect 163212 201218 163296 201454
rect 163532 201218 163616 201454
rect 163852 201218 163936 201454
rect 164172 201218 164256 201454
rect 164492 201218 164576 201454
rect 164812 201218 164896 201454
rect 165132 201218 165216 201454
rect 165452 201218 165514 201454
rect 137314 201134 165514 201218
rect 137314 200898 137376 201134
rect 137612 200898 137696 201134
rect 137932 200898 138016 201134
rect 138252 200898 138336 201134
rect 138572 200898 138656 201134
rect 138892 200898 138976 201134
rect 139212 200898 139296 201134
rect 139532 200898 139616 201134
rect 139852 200898 139936 201134
rect 140172 200898 140256 201134
rect 140492 200898 140576 201134
rect 140812 200898 140896 201134
rect 141132 200898 141216 201134
rect 141452 200898 141536 201134
rect 141772 200898 141856 201134
rect 142092 200898 142176 201134
rect 142412 200898 142496 201134
rect 142732 200898 142816 201134
rect 143052 200898 143136 201134
rect 143372 200898 143456 201134
rect 143692 200898 143776 201134
rect 144012 200898 144096 201134
rect 144332 200898 144416 201134
rect 144652 200898 144736 201134
rect 144972 200898 145056 201134
rect 145292 200898 145376 201134
rect 145612 200898 145696 201134
rect 145932 200898 146016 201134
rect 146252 200898 146336 201134
rect 146572 200898 146656 201134
rect 146892 200898 146976 201134
rect 147212 200898 147296 201134
rect 147532 200898 147616 201134
rect 147852 200898 147936 201134
rect 148172 200898 148256 201134
rect 148492 200898 148576 201134
rect 148812 200898 148896 201134
rect 149132 200898 149216 201134
rect 149452 200898 149536 201134
rect 149772 200898 149856 201134
rect 150092 200898 150176 201134
rect 150412 200898 150496 201134
rect 150732 200898 150816 201134
rect 151052 200898 151136 201134
rect 151372 200898 151456 201134
rect 151692 200898 151776 201134
rect 152012 200898 152096 201134
rect 152332 200898 152416 201134
rect 152652 200898 152736 201134
rect 152972 200898 153056 201134
rect 153292 200898 153376 201134
rect 153612 200898 153696 201134
rect 153932 200898 154016 201134
rect 154252 200898 154336 201134
rect 154572 200898 154656 201134
rect 154892 200898 154976 201134
rect 155212 200898 155296 201134
rect 155532 200898 155616 201134
rect 155852 200898 155936 201134
rect 156172 200898 156256 201134
rect 156492 200898 156576 201134
rect 156812 200898 156896 201134
rect 157132 200898 157216 201134
rect 157452 200898 157536 201134
rect 157772 200898 157856 201134
rect 158092 200898 158176 201134
rect 158412 200898 158496 201134
rect 158732 200898 158816 201134
rect 159052 200898 159136 201134
rect 159372 200898 159456 201134
rect 159692 200898 159776 201134
rect 160012 200898 160096 201134
rect 160332 200898 160416 201134
rect 160652 200898 160736 201134
rect 160972 200898 161056 201134
rect 161292 200898 161376 201134
rect 161612 200898 161696 201134
rect 161932 200898 162016 201134
rect 162252 200898 162336 201134
rect 162572 200898 162656 201134
rect 162892 200898 162976 201134
rect 163212 200898 163296 201134
rect 163532 200898 163616 201134
rect 163852 200898 163936 201134
rect 164172 200898 164256 201134
rect 164492 200898 164576 201134
rect 164812 200898 164896 201134
rect 165132 200898 165216 201134
rect 165452 200898 165514 201134
rect 137314 200866 165514 200898
rect 144683 200700 144749 200701
rect 144683 200636 144684 200700
rect 144748 200636 144749 200700
rect 144683 200635 144749 200636
rect 144686 195669 144746 200635
rect 149835 196348 149901 196349
rect 149835 196284 149836 196348
rect 149900 196284 149901 196348
rect 149835 196283 149901 196284
rect 144683 195668 144749 195669
rect 144683 195604 144684 195668
rect 144748 195604 144749 195668
rect 144683 195603 144749 195604
rect 148731 194716 148797 194717
rect 148731 194652 148732 194716
rect 148796 194652 148797 194716
rect 148731 194651 148797 194652
rect 143579 191808 143645 191809
rect 143579 191744 143580 191808
rect 143644 191744 143645 191808
rect 143579 191743 143645 191744
rect 141739 191316 141805 191317
rect 141739 191252 141740 191316
rect 141804 191252 141805 191316
rect 141739 191251 141805 191252
rect 140635 186964 140701 186965
rect 140635 186900 140636 186964
rect 140700 186900 140701 186964
rect 140635 186899 140701 186900
rect 140451 179212 140517 179213
rect 140451 179148 140452 179212
rect 140516 179148 140517 179212
rect 140451 179147 140517 179148
rect 132294 169718 132326 169954
rect 132562 169718 132646 169954
rect 132882 169718 132914 169954
rect 132294 169634 132914 169718
rect 132294 169398 132326 169634
rect 132562 169398 132646 169634
rect 132882 169398 132914 169634
rect 132294 142000 132914 169398
rect 140454 143173 140514 179147
rect 140451 143172 140517 143173
rect 140451 143108 140452 143172
rect 140516 143108 140517 143172
rect 140451 143107 140517 143108
rect 140638 142765 140698 186899
rect 141742 166429 141802 191251
rect 141923 190636 141989 190637
rect 141923 190572 141924 190636
rect 141988 190572 141989 190636
rect 141923 190571 141989 190572
rect 141739 166428 141805 166429
rect 141739 166364 141740 166428
rect 141804 166364 141805 166428
rect 141739 166363 141805 166364
rect 141926 166293 141986 190571
rect 142659 178804 142725 178805
rect 142659 178740 142660 178804
rect 142724 178740 142725 178804
rect 142659 178739 142725 178740
rect 142662 176765 142722 178739
rect 142659 176764 142725 176765
rect 142659 176700 142660 176764
rect 142724 176700 142725 176764
rect 142659 176699 142725 176700
rect 142291 173908 142357 173909
rect 142291 173844 142292 173908
rect 142356 173844 142357 173908
rect 142291 173843 142357 173844
rect 142107 171324 142173 171325
rect 142107 171260 142108 171324
rect 142172 171260 142173 171324
rect 142107 171259 142173 171260
rect 142110 170917 142170 171259
rect 142107 170916 142173 170917
rect 142107 170852 142108 170916
rect 142172 170852 142173 170916
rect 142107 170851 142173 170852
rect 141923 166292 141989 166293
rect 141923 166228 141924 166292
rect 141988 166228 141989 166292
rect 141923 166227 141989 166228
rect 142107 162212 142173 162213
rect 142107 162210 142108 162212
rect 141926 162150 142108 162210
rect 140635 142764 140701 142765
rect 140635 142700 140636 142764
rect 140700 142700 140701 142764
rect 140635 142699 140701 142700
rect 141926 142490 141986 162150
rect 142107 162148 142108 162150
rect 142172 162148 142173 162212
rect 142107 162147 142173 162148
rect 142294 143445 142354 173843
rect 142659 173772 142725 173773
rect 142659 173708 142660 173772
rect 142724 173708 142725 173772
rect 142659 173707 142725 173708
rect 142475 173636 142541 173637
rect 142475 173572 142476 173636
rect 142540 173572 142541 173636
rect 142475 173571 142541 173572
rect 142291 143444 142357 143445
rect 142291 143380 142292 143444
rect 142356 143380 142357 143444
rect 142291 143379 142357 143380
rect 142478 143309 142538 173571
rect 142475 143308 142541 143309
rect 142475 143244 142476 143308
rect 142540 143244 142541 143308
rect 142475 143243 142541 143244
rect 142107 142492 142173 142493
rect 142107 142490 142108 142492
rect 141926 142430 142108 142490
rect 142107 142428 142108 142430
rect 142172 142428 142173 142492
rect 142107 142427 142173 142428
rect 142662 142221 142722 173707
rect 143582 142629 143642 191743
rect 148734 191045 148794 194651
rect 148731 191044 148797 191045
rect 148731 190980 148732 191044
rect 148796 190980 148797 191044
rect 148731 190979 148797 190980
rect 149838 190637 149898 196283
rect 151307 196076 151373 196077
rect 151307 196012 151308 196076
rect 151372 196012 151373 196076
rect 151307 196011 151373 196012
rect 151310 191319 151370 196011
rect 151307 191318 151373 191319
rect 151307 191254 151308 191318
rect 151372 191254 151373 191318
rect 151307 191253 151373 191254
rect 149835 190636 149901 190637
rect 149835 190572 149836 190636
rect 149900 190572 149901 190636
rect 149835 190571 149901 190572
rect 146155 180708 146221 180709
rect 146155 180644 146156 180708
rect 146220 180644 146221 180708
rect 146155 180643 146221 180644
rect 144131 173772 144197 173773
rect 144131 173708 144132 173772
rect 144196 173708 144197 173772
rect 144131 173707 144197 173708
rect 144134 143037 144194 173707
rect 144131 143036 144197 143037
rect 144131 142972 144132 143036
rect 144196 142972 144197 143036
rect 144131 142971 144197 142972
rect 146158 142901 146218 180643
rect 168294 169954 168914 205398
rect 168294 169718 168326 169954
rect 168562 169718 168646 169954
rect 168882 169718 168914 169954
rect 168294 169634 168914 169718
rect 168294 169398 168326 169634
rect 168562 169398 168646 169634
rect 168882 169398 168914 169634
rect 146155 142900 146221 142901
rect 146155 142836 146156 142900
rect 146220 142836 146221 142900
rect 146155 142835 146221 142836
rect 143579 142628 143645 142629
rect 143579 142564 143580 142628
rect 143644 142564 143645 142628
rect 143579 142563 143645 142564
rect 142659 142220 142725 142221
rect 142659 142156 142660 142220
rect 142724 142156 142725 142220
rect 142659 142155 142725 142156
rect 168294 142000 168914 169398
rect 172794 210454 173414 228484
rect 172794 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 173414 210454
rect 172794 210134 173414 210218
rect 172794 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 173414 210134
rect 172794 174454 173414 209898
rect 172794 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 173414 174454
rect 172794 174134 173414 174218
rect 172794 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 173414 174134
rect 172794 142000 173414 173898
rect 177294 214954 177914 228484
rect 177294 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 177914 214954
rect 177294 214634 177914 214718
rect 177294 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 177914 214634
rect 177294 178954 177914 214398
rect 177294 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 177914 178954
rect 177294 178634 177914 178718
rect 177294 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 177914 178634
rect 177294 142954 177914 178398
rect 177294 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 177914 142954
rect 177294 142634 177914 142718
rect 177294 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 177914 142634
rect 177294 142000 177914 142398
rect 181794 219454 182414 228484
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 142000 182414 146898
rect 186294 223954 186914 228484
rect 186294 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 186914 223954
rect 186294 223634 186914 223718
rect 186294 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 186914 223634
rect 186294 187954 186914 223398
rect 186294 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 186914 187954
rect 186294 187634 186914 187718
rect 186294 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 186914 187634
rect 186294 151954 186914 187398
rect 186294 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 186914 151954
rect 186294 151634 186914 151718
rect 186294 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 186914 151634
rect 114294 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 114914 115954
rect 114294 115634 114914 115718
rect 114294 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 114914 115634
rect 114294 79954 114914 115398
rect 139568 115954 139888 115986
rect 139568 115718 139610 115954
rect 139846 115718 139888 115954
rect 139568 115634 139888 115718
rect 139568 115398 139610 115634
rect 139846 115398 139888 115634
rect 139568 115366 139888 115398
rect 170288 115954 170608 115986
rect 170288 115718 170330 115954
rect 170566 115718 170608 115954
rect 170288 115634 170608 115718
rect 170288 115398 170330 115634
rect 170566 115398 170608 115634
rect 170288 115366 170608 115398
rect 186294 115954 186914 151398
rect 186294 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 186914 115954
rect 186294 115634 186914 115718
rect 186294 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 186914 115634
rect 124208 111454 124528 111486
rect 124208 111218 124250 111454
rect 124486 111218 124528 111454
rect 124208 111134 124528 111218
rect 124208 110898 124250 111134
rect 124486 110898 124528 111134
rect 124208 110866 124528 110898
rect 154928 111454 155248 111486
rect 154928 111218 154970 111454
rect 155206 111218 155248 111454
rect 154928 111134 155248 111218
rect 154928 110898 154970 111134
rect 155206 110898 155248 111134
rect 154928 110866 155248 110898
rect 172283 80476 172349 80477
rect 172283 80412 172284 80476
rect 172348 80412 172349 80476
rect 172283 80411 172349 80412
rect 171547 80340 171613 80341
rect 171547 80276 171548 80340
rect 171612 80276 171613 80340
rect 171547 80275 171613 80276
rect 159403 80204 159469 80205
rect 159403 80140 159404 80204
rect 159468 80140 159469 80204
rect 159403 80139 159469 80140
rect 114294 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 114914 79954
rect 125915 79932 125981 79933
rect 125915 79868 125916 79932
rect 125980 79868 125981 79932
rect 125915 79867 125981 79868
rect 127571 79932 127637 79933
rect 127571 79868 127572 79932
rect 127636 79868 127637 79932
rect 127571 79867 127637 79868
rect 128307 79932 128373 79933
rect 128307 79868 128308 79932
rect 128372 79868 128373 79932
rect 128307 79867 128373 79868
rect 128859 79932 128925 79933
rect 128859 79868 128860 79932
rect 128924 79868 128925 79932
rect 128859 79867 128925 79868
rect 129043 79932 129109 79933
rect 129043 79868 129044 79932
rect 129108 79868 129109 79932
rect 129043 79867 129109 79868
rect 129779 79932 129845 79933
rect 129779 79868 129780 79932
rect 129844 79868 129845 79932
rect 129779 79867 129845 79868
rect 130699 79932 130765 79933
rect 130699 79868 130700 79932
rect 130764 79868 130765 79932
rect 130699 79867 130765 79868
rect 131251 79932 131317 79933
rect 131251 79868 131252 79932
rect 131316 79868 131317 79932
rect 131251 79867 131317 79868
rect 131619 79932 131685 79933
rect 131619 79868 131620 79932
rect 131684 79868 131685 79932
rect 131619 79867 131685 79868
rect 131803 79932 131869 79933
rect 131803 79868 131804 79932
rect 131868 79868 131869 79932
rect 131803 79867 131869 79868
rect 133091 79932 133157 79933
rect 133091 79868 133092 79932
rect 133156 79868 133157 79932
rect 133091 79867 133157 79868
rect 133827 79932 133893 79933
rect 133827 79868 133828 79932
rect 133892 79868 133893 79932
rect 133827 79867 133893 79868
rect 135483 79932 135549 79933
rect 135483 79868 135484 79932
rect 135548 79868 135549 79932
rect 135483 79867 135549 79868
rect 135851 79932 135917 79933
rect 135851 79868 135852 79932
rect 135916 79868 135917 79932
rect 135851 79867 135917 79868
rect 137691 79932 137757 79933
rect 137691 79868 137692 79932
rect 137756 79868 137757 79932
rect 137691 79867 137757 79868
rect 138427 79932 138493 79933
rect 138427 79868 138428 79932
rect 138492 79868 138493 79932
rect 138427 79867 138493 79868
rect 140267 79932 140333 79933
rect 140267 79868 140268 79932
rect 140332 79868 140333 79932
rect 140267 79867 140333 79868
rect 141003 79932 141069 79933
rect 141003 79868 141004 79932
rect 141068 79868 141069 79932
rect 141003 79867 141069 79868
rect 142659 79932 142725 79933
rect 142659 79868 142660 79932
rect 142724 79868 142725 79932
rect 142659 79867 142725 79868
rect 143763 79932 143829 79933
rect 143763 79868 143764 79932
rect 143828 79868 143829 79932
rect 143763 79867 143829 79868
rect 144315 79932 144381 79933
rect 144315 79868 144316 79932
rect 144380 79868 144381 79932
rect 144315 79867 144381 79868
rect 145603 79932 145669 79933
rect 145603 79868 145604 79932
rect 145668 79868 145669 79932
rect 145603 79867 145669 79868
rect 146891 79932 146957 79933
rect 146891 79868 146892 79932
rect 146956 79868 146957 79932
rect 146891 79867 146957 79868
rect 147259 79932 147325 79933
rect 147259 79868 147260 79932
rect 147324 79868 147325 79932
rect 147259 79867 147325 79868
rect 148363 79932 148429 79933
rect 148363 79868 148364 79932
rect 148428 79868 148429 79932
rect 148363 79867 148429 79868
rect 148731 79932 148797 79933
rect 148731 79868 148732 79932
rect 148796 79868 148797 79932
rect 148731 79867 148797 79868
rect 149835 79932 149901 79933
rect 149835 79868 149836 79932
rect 149900 79868 149901 79932
rect 149835 79867 149901 79868
rect 151675 79932 151741 79933
rect 151675 79868 151676 79932
rect 151740 79868 151741 79932
rect 152963 79932 153029 79933
rect 152963 79930 152964 79932
rect 151675 79867 151741 79868
rect 152598 79870 152964 79930
rect 114294 79634 114914 79718
rect 114294 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 114914 79634
rect 114294 43954 114914 79398
rect 125731 78708 125797 78709
rect 125731 78644 125732 78708
rect 125796 78644 125797 78708
rect 125731 78643 125797 78644
rect 114294 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 114914 43954
rect 114294 43634 114914 43718
rect 114294 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 114914 43634
rect 114294 7954 114914 43398
rect 114294 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 114914 7954
rect 114294 7634 114914 7718
rect 114294 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 114914 7634
rect 114294 -1306 114914 7398
rect 114294 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 114914 -1306
rect 114294 -1626 114914 -1542
rect 114294 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 114914 -1626
rect 114294 -7654 114914 -1862
rect 118794 48454 119414 78000
rect 118794 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 119414 48454
rect 118794 48134 119414 48218
rect 118794 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 119414 48134
rect 118794 12454 119414 47898
rect 118794 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 119414 12454
rect 118794 12134 119414 12218
rect 118794 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 119414 12134
rect 118794 -2266 119414 11898
rect 118794 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 119414 -2266
rect 118794 -2586 119414 -2502
rect 118794 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 119414 -2586
rect 118794 -7654 119414 -2822
rect 123294 52954 123914 78000
rect 125734 72453 125794 78643
rect 125918 74493 125978 79867
rect 127387 79796 127453 79797
rect 127387 79732 127388 79796
rect 127452 79732 127453 79796
rect 127387 79731 127453 79732
rect 126099 78844 126165 78845
rect 126099 78780 126100 78844
rect 126164 78780 126165 78844
rect 126099 78779 126165 78780
rect 125915 74492 125981 74493
rect 125915 74428 125916 74492
rect 125980 74428 125981 74492
rect 125915 74427 125981 74428
rect 125731 72452 125797 72453
rect 125731 72388 125732 72452
rect 125796 72388 125797 72452
rect 125731 72387 125797 72388
rect 123294 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 123914 52954
rect 123294 52634 123914 52718
rect 123294 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 123914 52634
rect 123294 16954 123914 52398
rect 123294 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 123914 16954
rect 123294 16634 123914 16718
rect 123294 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 123914 16634
rect 123294 -3226 123914 16398
rect 126102 4861 126162 78779
rect 127203 78708 127269 78709
rect 127203 78644 127204 78708
rect 127268 78644 127269 78708
rect 127203 78643 127269 78644
rect 127206 68237 127266 78643
rect 127203 68236 127269 68237
rect 127203 68172 127204 68236
rect 127268 68172 127269 68236
rect 127203 68171 127269 68172
rect 127390 25533 127450 79731
rect 127574 78301 127634 79867
rect 127571 78300 127637 78301
rect 127571 78236 127572 78300
rect 127636 78236 127637 78300
rect 127571 78235 127637 78236
rect 128310 78165 128370 79867
rect 128307 78164 128373 78165
rect 128307 78100 128308 78164
rect 128372 78100 128373 78164
rect 128307 78099 128373 78100
rect 128491 78164 128557 78165
rect 128491 78100 128492 78164
rect 128556 78100 128557 78164
rect 128491 78099 128557 78100
rect 127794 57454 128414 78000
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127387 25532 127453 25533
rect 127387 25468 127388 25532
rect 127452 25468 127453 25532
rect 127387 25467 127453 25468
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 126099 4860 126165 4861
rect 126099 4796 126100 4860
rect 126164 4796 126165 4860
rect 126099 4795 126165 4796
rect 123294 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 123914 -3226
rect 123294 -3546 123914 -3462
rect 123294 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 123914 -3546
rect 123294 -7654 123914 -3782
rect 127794 -4186 128414 20898
rect 128494 16590 128554 78099
rect 128675 77348 128741 77349
rect 128675 77284 128676 77348
rect 128740 77284 128741 77348
rect 128675 77283 128741 77284
rect 128678 73813 128738 77283
rect 128675 73812 128741 73813
rect 128675 73748 128676 73812
rect 128740 73748 128741 73812
rect 128675 73747 128741 73748
rect 128862 72589 128922 79867
rect 129046 75989 129106 79867
rect 129043 75988 129109 75989
rect 129043 75924 129044 75988
rect 129108 75924 129109 75988
rect 129043 75923 129109 75924
rect 128859 72588 128925 72589
rect 128859 72524 128860 72588
rect 128924 72524 128925 72588
rect 128859 72523 128925 72524
rect 128494 16530 128738 16590
rect 128678 7581 128738 16530
rect 129782 8941 129842 79867
rect 130147 79660 130213 79661
rect 130147 79596 130148 79660
rect 130212 79596 130213 79660
rect 130147 79595 130213 79596
rect 130515 79660 130581 79661
rect 130515 79596 130516 79660
rect 130580 79596 130581 79660
rect 130515 79595 130581 79596
rect 129963 78844 130029 78845
rect 129963 78780 129964 78844
rect 130028 78780 130029 78844
rect 129963 78779 130029 78780
rect 129966 9077 130026 78779
rect 130150 68373 130210 79595
rect 130518 78845 130578 79595
rect 130515 78844 130581 78845
rect 130515 78780 130516 78844
rect 130580 78780 130581 78844
rect 130515 78779 130581 78780
rect 130331 78708 130397 78709
rect 130331 78644 130332 78708
rect 130396 78644 130397 78708
rect 130331 78643 130397 78644
rect 130334 69597 130394 78643
rect 130702 76533 130762 79867
rect 130699 76532 130765 76533
rect 130699 76468 130700 76532
rect 130764 76468 130765 76532
rect 130699 76467 130765 76468
rect 130331 69596 130397 69597
rect 130331 69532 130332 69596
rect 130396 69532 130397 69596
rect 130331 69531 130397 69532
rect 130147 68372 130213 68373
rect 130147 68308 130148 68372
rect 130212 68308 130213 68372
rect 130147 68307 130213 68308
rect 131254 65517 131314 79867
rect 131435 76668 131501 76669
rect 131435 76604 131436 76668
rect 131500 76604 131501 76668
rect 131435 76603 131501 76604
rect 131251 65516 131317 65517
rect 131251 65452 131252 65516
rect 131316 65452 131317 65516
rect 131251 65451 131317 65452
rect 131438 44845 131498 76603
rect 131622 75173 131682 79867
rect 131806 76669 131866 79867
rect 131803 76668 131869 76669
rect 131803 76604 131804 76668
rect 131868 76604 131869 76668
rect 131803 76603 131869 76604
rect 131619 75172 131685 75173
rect 131619 75108 131620 75172
rect 131684 75108 131685 75172
rect 131619 75107 131685 75108
rect 132294 61954 132914 78000
rect 132294 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 132914 61954
rect 132294 61634 132914 61718
rect 132294 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 132914 61634
rect 131435 44844 131501 44845
rect 131435 44780 131436 44844
rect 131500 44780 131501 44844
rect 131435 44779 131501 44780
rect 132294 25954 132914 61398
rect 132294 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 132914 25954
rect 132294 25634 132914 25718
rect 132294 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 132914 25634
rect 129963 9076 130029 9077
rect 129963 9012 129964 9076
rect 130028 9012 130029 9076
rect 129963 9011 130029 9012
rect 129779 8940 129845 8941
rect 129779 8876 129780 8940
rect 129844 8876 129845 8940
rect 129779 8875 129845 8876
rect 128675 7580 128741 7581
rect 128675 7516 128676 7580
rect 128740 7516 128741 7580
rect 128675 7515 128741 7516
rect 127794 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 128414 -4186
rect 127794 -4506 128414 -4422
rect 127794 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 128414 -4506
rect 127794 -7654 128414 -4742
rect 132294 -5146 132914 25398
rect 133094 9213 133154 79867
rect 133275 79796 133341 79797
rect 133275 79732 133276 79796
rect 133340 79732 133341 79796
rect 133275 79731 133341 79732
rect 133278 69733 133338 79731
rect 133643 77892 133709 77893
rect 133643 77828 133644 77892
rect 133708 77828 133709 77892
rect 133643 77827 133709 77828
rect 133275 69732 133341 69733
rect 133275 69668 133276 69732
rect 133340 69668 133341 69732
rect 133275 69667 133341 69668
rect 133646 9485 133706 77827
rect 133643 9484 133709 9485
rect 133643 9420 133644 9484
rect 133708 9420 133709 9484
rect 133643 9419 133709 9420
rect 133091 9212 133157 9213
rect 133091 9148 133092 9212
rect 133156 9148 133157 9212
rect 133091 9147 133157 9148
rect 133830 7717 133890 79867
rect 135486 77310 135546 79867
rect 135854 78709 135914 79867
rect 135851 78708 135917 78709
rect 135851 78644 135852 78708
rect 135916 78644 135917 78708
rect 135851 78643 135917 78644
rect 135302 77250 135546 77310
rect 134011 76668 134077 76669
rect 134011 76604 134012 76668
rect 134076 76604 134077 76668
rect 134011 76603 134077 76604
rect 135115 76668 135181 76669
rect 135115 76604 135116 76668
rect 135180 76604 135181 76668
rect 135115 76603 135181 76604
rect 134014 10301 134074 76603
rect 134011 10300 134077 10301
rect 134011 10236 134012 10300
rect 134076 10236 134077 10300
rect 134011 10235 134077 10236
rect 133827 7716 133893 7717
rect 133827 7652 133828 7716
rect 133892 7652 133893 7716
rect 133827 7651 133893 7652
rect 135118 3365 135178 76603
rect 135302 68237 135362 77250
rect 136219 76940 136285 76941
rect 136219 76876 136220 76940
rect 136284 76876 136285 76940
rect 136219 76875 136285 76876
rect 136035 76804 136101 76805
rect 136035 76740 136036 76804
rect 136100 76740 136101 76804
rect 136035 76739 136101 76740
rect 135299 68236 135365 68237
rect 135299 68172 135300 68236
rect 135364 68172 135365 68236
rect 135299 68171 135365 68172
rect 136038 3909 136098 76739
rect 136035 3908 136101 3909
rect 136035 3844 136036 3908
rect 136100 3844 136101 3908
rect 136035 3843 136101 3844
rect 136222 3637 136282 76875
rect 136403 76532 136469 76533
rect 136403 76468 136404 76532
rect 136468 76468 136469 76532
rect 136403 76467 136469 76468
rect 136219 3636 136285 3637
rect 136219 3572 136220 3636
rect 136284 3572 136285 3636
rect 136219 3571 136285 3572
rect 136406 3501 136466 76467
rect 136794 66454 137414 78000
rect 136794 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 137414 66454
rect 136794 66134 137414 66218
rect 136794 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 137414 66134
rect 136794 30454 137414 65898
rect 137694 43485 137754 79867
rect 137875 79796 137941 79797
rect 137875 79732 137876 79796
rect 137940 79732 137941 79796
rect 137875 79731 137941 79732
rect 137691 43484 137757 43485
rect 137691 43420 137692 43484
rect 137756 43420 137757 43484
rect 137691 43419 137757 43420
rect 136794 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 137414 30454
rect 136794 30134 137414 30218
rect 136794 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 137414 30134
rect 136403 3500 136469 3501
rect 136403 3436 136404 3500
rect 136468 3436 136469 3500
rect 136403 3435 136469 3436
rect 135115 3364 135181 3365
rect 135115 3300 135116 3364
rect 135180 3300 135181 3364
rect 135115 3299 135181 3300
rect 132294 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 132914 -5146
rect 132294 -5466 132914 -5382
rect 132294 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 132914 -5466
rect 132294 -7654 132914 -5702
rect 136794 -6106 137414 29898
rect 137878 6221 137938 79731
rect 138430 76533 138490 79867
rect 138611 79796 138677 79797
rect 138611 79732 138612 79796
rect 138676 79732 138677 79796
rect 138611 79731 138677 79732
rect 138427 76532 138493 76533
rect 138427 76468 138428 76532
rect 138492 76468 138493 76532
rect 138427 76467 138493 76468
rect 138614 67013 138674 79731
rect 138979 76668 139045 76669
rect 138979 76604 138980 76668
rect 139044 76604 139045 76668
rect 138979 76603 139045 76604
rect 140083 76668 140149 76669
rect 140083 76604 140084 76668
rect 140148 76604 140149 76668
rect 140083 76603 140149 76604
rect 138982 69597 139042 76603
rect 138979 69596 139045 69597
rect 138979 69532 138980 69596
rect 139044 69532 139045 69596
rect 138979 69531 139045 69532
rect 138611 67012 138677 67013
rect 138611 66948 138612 67012
rect 138676 66948 138677 67012
rect 138611 66947 138677 66948
rect 140086 27029 140146 76603
rect 140270 66877 140330 79867
rect 140451 79796 140517 79797
rect 140451 79732 140452 79796
rect 140516 79732 140517 79796
rect 140451 79731 140517 79732
rect 140267 66876 140333 66877
rect 140267 66812 140268 66876
rect 140332 66812 140333 66876
rect 140267 66811 140333 66812
rect 140454 47837 140514 79731
rect 140451 47836 140517 47837
rect 140451 47772 140452 47836
rect 140516 47772 140517 47836
rect 140451 47771 140517 47772
rect 140083 27028 140149 27029
rect 140083 26964 140084 27028
rect 140148 26964 140149 27028
rect 140083 26963 140149 26964
rect 141006 17373 141066 79867
rect 141294 70954 141914 78000
rect 142662 76397 142722 79867
rect 143211 76668 143277 76669
rect 143211 76604 143212 76668
rect 143276 76604 143277 76668
rect 143211 76603 143277 76604
rect 143395 76668 143461 76669
rect 143395 76604 143396 76668
rect 143460 76604 143461 76668
rect 143395 76603 143461 76604
rect 143027 76532 143093 76533
rect 143027 76468 143028 76532
rect 143092 76468 143093 76532
rect 143027 76467 143093 76468
rect 142659 76396 142725 76397
rect 142659 76332 142660 76396
rect 142724 76332 142725 76396
rect 142659 76331 142725 76332
rect 141294 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 141914 70954
rect 141294 70634 141914 70718
rect 141294 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 141914 70634
rect 141294 34954 141914 70398
rect 143030 61437 143090 76467
rect 143027 61436 143093 61437
rect 143027 61372 143028 61436
rect 143092 61372 143093 61436
rect 143027 61371 143093 61372
rect 141294 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 141914 34954
rect 141294 34634 141914 34718
rect 141294 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 141914 34634
rect 141003 17372 141069 17373
rect 141003 17308 141004 17372
rect 141068 17308 141069 17372
rect 141003 17307 141069 17308
rect 137875 6220 137941 6221
rect 137875 6156 137876 6220
rect 137940 6156 137941 6220
rect 137875 6155 137941 6156
rect 136794 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 137414 -6106
rect 136794 -6426 137414 -6342
rect 136794 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 137414 -6426
rect 136794 -7654 137414 -6662
rect 141294 -7066 141914 34398
rect 143214 32741 143274 76603
rect 143211 32740 143277 32741
rect 143211 32676 143212 32740
rect 143276 32676 143277 32740
rect 143211 32675 143277 32676
rect 143398 13293 143458 76603
rect 143766 74221 143826 79867
rect 144318 76669 144378 79867
rect 145235 79796 145301 79797
rect 145235 79732 145236 79796
rect 145300 79732 145301 79796
rect 145235 79731 145301 79732
rect 144499 76804 144565 76805
rect 144499 76740 144500 76804
rect 144564 76740 144565 76804
rect 144499 76739 144565 76740
rect 144315 76668 144381 76669
rect 144315 76604 144316 76668
rect 144380 76604 144381 76668
rect 144315 76603 144381 76604
rect 144131 76532 144197 76533
rect 144131 76468 144132 76532
rect 144196 76468 144197 76532
rect 144131 76467 144197 76468
rect 143763 74220 143829 74221
rect 143763 74156 143764 74220
rect 143828 74156 143829 74220
rect 143763 74155 143829 74156
rect 144134 20093 144194 76467
rect 144502 64293 144562 76739
rect 144499 64292 144565 64293
rect 144499 64228 144500 64292
rect 144564 64228 144565 64292
rect 144499 64227 144565 64228
rect 145238 62933 145298 79731
rect 145419 76668 145485 76669
rect 145419 76604 145420 76668
rect 145484 76604 145485 76668
rect 145419 76603 145485 76604
rect 145235 62932 145301 62933
rect 145235 62868 145236 62932
rect 145300 62868 145301 62932
rect 145235 62867 145301 62868
rect 145422 52053 145482 76603
rect 145419 52052 145485 52053
rect 145419 51988 145420 52052
rect 145484 51988 145485 52052
rect 145419 51987 145485 51988
rect 145606 39269 145666 79867
rect 146523 79796 146589 79797
rect 146523 79732 146524 79796
rect 146588 79732 146589 79796
rect 146523 79731 146589 79732
rect 146707 79796 146773 79797
rect 146707 79732 146708 79796
rect 146772 79732 146773 79796
rect 146707 79731 146773 79732
rect 145794 75454 146414 78000
rect 146526 76533 146586 79731
rect 146710 76805 146770 79731
rect 146707 76804 146773 76805
rect 146707 76740 146708 76804
rect 146772 76740 146773 76804
rect 146707 76739 146773 76740
rect 146894 76669 146954 79867
rect 146891 76668 146957 76669
rect 146891 76604 146892 76668
rect 146956 76604 146957 76668
rect 146891 76603 146957 76604
rect 146523 76532 146589 76533
rect 146523 76468 146524 76532
rect 146588 76468 146589 76532
rect 146523 76467 146589 76468
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 147075 75036 147141 75037
rect 147075 74972 147076 75036
rect 147140 74972 147141 75036
rect 147075 74971 147141 74972
rect 145794 39454 146414 74898
rect 145603 39268 145669 39269
rect 145603 39204 145604 39268
rect 145668 39204 145669 39268
rect 145603 39203 145669 39204
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 144131 20092 144197 20093
rect 144131 20028 144132 20092
rect 144196 20028 144197 20092
rect 144131 20027 144197 20028
rect 143395 13292 143461 13293
rect 143395 13228 143396 13292
rect 143460 13228 143461 13292
rect 143395 13227 143461 13228
rect 141294 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 141914 -7066
rect 141294 -7386 141914 -7302
rect 141294 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 141914 -7386
rect 141294 -7654 141914 -7622
rect 145794 3454 146414 38898
rect 147078 3773 147138 74971
rect 147262 9621 147322 79867
rect 148366 74493 148426 79867
rect 148547 79796 148613 79797
rect 148547 79732 148548 79796
rect 148612 79732 148613 79796
rect 148547 79731 148613 79732
rect 148363 74492 148429 74493
rect 148363 74428 148364 74492
rect 148428 74428 148429 74492
rect 148363 74427 148429 74428
rect 148550 17237 148610 79731
rect 148547 17236 148613 17237
rect 148547 17172 148548 17236
rect 148612 17172 148613 17236
rect 148547 17171 148613 17172
rect 147259 9620 147325 9621
rect 147259 9556 147260 9620
rect 147324 9556 147325 9620
rect 147259 9555 147325 9556
rect 148734 6493 148794 79867
rect 148915 76668 148981 76669
rect 148915 76604 148916 76668
rect 148980 76604 148981 76668
rect 148915 76603 148981 76604
rect 148918 6629 148978 76603
rect 149651 75172 149717 75173
rect 149651 75108 149652 75172
rect 149716 75108 149717 75172
rect 149651 75107 149717 75108
rect 149654 55997 149714 75107
rect 149651 55996 149717 55997
rect 149651 55932 149652 55996
rect 149716 55932 149717 55996
rect 149651 55931 149717 55932
rect 149838 42125 149898 79867
rect 150019 79796 150085 79797
rect 150019 79732 150020 79796
rect 150084 79732 150085 79796
rect 150019 79731 150085 79732
rect 149835 42124 149901 42125
rect 149835 42060 149836 42124
rect 149900 42060 149901 42124
rect 149835 42059 149901 42060
rect 150022 26893 150082 79731
rect 151491 78844 151557 78845
rect 151491 78780 151492 78844
rect 151556 78780 151557 78844
rect 151491 78779 151557 78780
rect 151307 78708 151373 78709
rect 151307 78644 151308 78708
rect 151372 78644 151373 78708
rect 151307 78643 151373 78644
rect 150294 43954 150914 78000
rect 151310 51917 151370 78643
rect 151307 51916 151373 51917
rect 151307 51852 151308 51916
rect 151372 51852 151373 51916
rect 151307 51851 151373 51852
rect 150294 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 150914 43954
rect 150294 43634 150914 43718
rect 150294 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 150914 43634
rect 150019 26892 150085 26893
rect 150019 26828 150020 26892
rect 150084 26828 150085 26892
rect 150019 26827 150085 26828
rect 150294 7954 150914 43398
rect 151494 35325 151554 78779
rect 151491 35324 151557 35325
rect 151491 35260 151492 35324
rect 151556 35260 151557 35324
rect 151491 35259 151557 35260
rect 151678 11797 151738 79867
rect 152411 79796 152477 79797
rect 152411 79732 152412 79796
rect 152476 79732 152477 79796
rect 152411 79731 152477 79732
rect 151859 79660 151925 79661
rect 151859 79596 151860 79660
rect 151924 79596 151925 79660
rect 151859 79595 151925 79596
rect 151862 77485 151922 79595
rect 151859 77484 151925 77485
rect 151859 77420 151860 77484
rect 151924 77420 151925 77484
rect 151859 77419 151925 77420
rect 152414 35189 152474 79731
rect 152598 68373 152658 79870
rect 152963 79868 152964 79870
rect 153028 79868 153029 79932
rect 152963 79867 153029 79868
rect 153699 79932 153765 79933
rect 153699 79868 153700 79932
rect 153764 79868 153765 79932
rect 153699 79867 153765 79868
rect 153883 79932 153949 79933
rect 153883 79868 153884 79932
rect 153948 79868 153949 79932
rect 153883 79867 153949 79868
rect 156827 79932 156893 79933
rect 156827 79868 156828 79932
rect 156892 79868 156893 79932
rect 156827 79867 156893 79868
rect 158115 79932 158181 79933
rect 158115 79868 158116 79932
rect 158180 79868 158181 79932
rect 158115 79867 158181 79868
rect 153702 78029 153762 79867
rect 153699 78028 153765 78029
rect 153699 77964 153700 78028
rect 153764 77964 153765 78028
rect 153699 77963 153765 77964
rect 152779 77348 152845 77349
rect 152779 77284 152780 77348
rect 152844 77284 152845 77348
rect 152779 77283 152845 77284
rect 152595 68372 152661 68373
rect 152595 68308 152596 68372
rect 152660 68308 152661 68372
rect 152595 68307 152661 68308
rect 152782 47701 152842 77283
rect 153886 51781 153946 79867
rect 154067 79796 154133 79797
rect 154067 79732 154068 79796
rect 154132 79732 154133 79796
rect 154067 79731 154133 79732
rect 154987 79796 155053 79797
rect 154987 79732 154988 79796
rect 155052 79732 155053 79796
rect 154987 79731 155053 79732
rect 155907 79796 155973 79797
rect 155907 79732 155908 79796
rect 155972 79732 155973 79796
rect 155907 79731 155973 79732
rect 156643 79796 156709 79797
rect 156643 79732 156644 79796
rect 156708 79732 156709 79796
rect 156643 79731 156709 79732
rect 153883 51780 153949 51781
rect 153883 51716 153884 51780
rect 153948 51716 153949 51780
rect 153883 51715 153949 51716
rect 152779 47700 152845 47701
rect 152779 47636 152780 47700
rect 152844 47636 152845 47700
rect 152779 47635 152845 47636
rect 152411 35188 152477 35189
rect 152411 35124 152412 35188
rect 152476 35124 152477 35188
rect 152411 35123 152477 35124
rect 154070 21589 154130 79731
rect 154990 78709 155050 79731
rect 154987 78708 155053 78709
rect 154987 78644 154988 78708
rect 155052 78644 155053 78708
rect 154987 78643 155053 78644
rect 154251 78164 154317 78165
rect 154251 78100 154252 78164
rect 154316 78100 154317 78164
rect 154251 78099 154317 78100
rect 154067 21588 154133 21589
rect 154067 21524 154068 21588
rect 154132 21524 154133 21588
rect 154067 21523 154133 21524
rect 154254 15877 154314 78099
rect 154435 77892 154501 77893
rect 154435 77828 154436 77892
rect 154500 77828 154501 77892
rect 154435 77827 154501 77828
rect 154251 15876 154317 15877
rect 154251 15812 154252 15876
rect 154316 15812 154317 15876
rect 154251 15811 154317 15812
rect 154438 13157 154498 77827
rect 154794 48454 155414 78000
rect 155723 77348 155789 77349
rect 155723 77284 155724 77348
rect 155788 77284 155789 77348
rect 155723 77283 155789 77284
rect 155726 55861 155786 77283
rect 155910 76669 155970 79731
rect 155907 76668 155973 76669
rect 155907 76604 155908 76668
rect 155972 76604 155973 76668
rect 155907 76603 155973 76604
rect 155723 55860 155789 55861
rect 155723 55796 155724 55860
rect 155788 55796 155789 55860
rect 155723 55795 155789 55796
rect 154794 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 155414 48454
rect 154794 48134 155414 48218
rect 154794 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 155414 48134
rect 154435 13156 154501 13157
rect 154435 13092 154436 13156
rect 154500 13092 154501 13156
rect 154435 13091 154501 13092
rect 154794 12454 155414 47898
rect 154794 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 155414 12454
rect 154794 12134 155414 12218
rect 154794 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 155414 12134
rect 151675 11796 151741 11797
rect 151675 11732 151676 11796
rect 151740 11732 151741 11796
rect 151675 11731 151741 11732
rect 150294 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 150914 7954
rect 150294 7634 150914 7718
rect 150294 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 150914 7634
rect 148915 6628 148981 6629
rect 148915 6564 148916 6628
rect 148980 6564 148981 6628
rect 148915 6563 148981 6564
rect 148731 6492 148797 6493
rect 148731 6428 148732 6492
rect 148796 6428 148797 6492
rect 148731 6427 148797 6428
rect 147075 3772 147141 3773
rect 147075 3708 147076 3772
rect 147140 3708 147141 3772
rect 147075 3707 147141 3708
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 150294 -1306 150914 7398
rect 150294 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 150914 -1306
rect 150294 -1626 150914 -1542
rect 150294 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 150914 -1626
rect 150294 -7654 150914 -1862
rect 154794 -2266 155414 11898
rect 156646 9349 156706 79731
rect 156830 47565 156890 79867
rect 157011 78844 157077 78845
rect 157011 78780 157012 78844
rect 157076 78780 157077 78844
rect 157011 78779 157077 78780
rect 157014 75581 157074 78779
rect 157195 78028 157261 78029
rect 157195 77964 157196 78028
rect 157260 77964 157261 78028
rect 157195 77963 157261 77964
rect 157931 78028 157997 78029
rect 157931 77964 157932 78028
rect 157996 77964 157997 78028
rect 157931 77963 157997 77964
rect 157011 75580 157077 75581
rect 157011 75516 157012 75580
rect 157076 75516 157077 75580
rect 157011 75515 157077 75516
rect 157198 70410 157258 77963
rect 157014 70350 157258 70410
rect 156827 47564 156893 47565
rect 156827 47500 156828 47564
rect 156892 47500 156893 47564
rect 156827 47499 156893 47500
rect 157014 18597 157074 70350
rect 157934 48925 157994 77963
rect 157931 48924 157997 48925
rect 157931 48860 157932 48924
rect 157996 48860 157997 48924
rect 157931 48859 157997 48860
rect 158118 19957 158178 79867
rect 158483 79796 158549 79797
rect 158483 79732 158484 79796
rect 158548 79732 158549 79796
rect 158483 79731 158549 79732
rect 158299 77892 158365 77893
rect 158299 77828 158300 77892
rect 158364 77828 158365 77892
rect 158299 77827 158365 77828
rect 158115 19956 158181 19957
rect 158115 19892 158116 19956
rect 158180 19892 158181 19956
rect 158115 19891 158181 19892
rect 157011 18596 157077 18597
rect 157011 18532 157012 18596
rect 157076 18532 157077 18596
rect 157011 18531 157077 18532
rect 158302 11661 158362 77827
rect 158299 11660 158365 11661
rect 158299 11596 158300 11660
rect 158364 11596 158365 11660
rect 158299 11595 158365 11596
rect 158486 10301 158546 79731
rect 159406 79253 159466 80139
rect 171317 79966 171383 79967
rect 160139 79932 160205 79933
rect 160139 79868 160140 79932
rect 160204 79868 160205 79932
rect 160139 79867 160205 79868
rect 160691 79932 160757 79933
rect 160691 79868 160692 79932
rect 160756 79868 160757 79932
rect 160691 79867 160757 79868
rect 161979 79932 162045 79933
rect 161979 79868 161980 79932
rect 162044 79868 162045 79932
rect 161979 79867 162045 79868
rect 162163 79932 162229 79933
rect 162163 79868 162164 79932
rect 162228 79868 162229 79932
rect 162163 79867 162229 79868
rect 163267 79932 163333 79933
rect 163267 79868 163268 79932
rect 163332 79868 163333 79932
rect 163267 79867 163333 79868
rect 163451 79932 163517 79933
rect 163451 79868 163452 79932
rect 163516 79868 163517 79932
rect 163451 79867 163517 79868
rect 164739 79932 164805 79933
rect 164739 79868 164740 79932
rect 164804 79868 164805 79932
rect 164739 79867 164805 79868
rect 165475 79932 165541 79933
rect 165475 79868 165476 79932
rect 165540 79868 165541 79932
rect 165475 79867 165541 79868
rect 166211 79932 166277 79933
rect 166211 79868 166212 79932
rect 166276 79868 166277 79932
rect 166211 79867 166277 79868
rect 168051 79932 168117 79933
rect 168051 79868 168052 79932
rect 168116 79868 168117 79932
rect 168051 79867 168117 79868
rect 168787 79932 168853 79933
rect 168787 79868 168788 79932
rect 168852 79868 168853 79932
rect 168787 79867 168853 79868
rect 169523 79932 169589 79933
rect 169523 79868 169524 79932
rect 169588 79868 169589 79932
rect 169523 79867 169589 79868
rect 170259 79932 170325 79933
rect 170259 79868 170260 79932
rect 170324 79868 170325 79932
rect 171317 79902 171318 79966
rect 171382 79930 171383 79966
rect 171550 79933 171610 80275
rect 171915 80204 171981 80205
rect 171915 80140 171916 80204
rect 171980 80202 171981 80204
rect 171980 80142 172162 80202
rect 171980 80140 171981 80142
rect 171915 80139 171981 80140
rect 171547 79932 171613 79933
rect 171382 79902 171426 79930
rect 171317 79901 171426 79902
rect 171320 79870 171426 79901
rect 170259 79867 170325 79868
rect 159771 79796 159837 79797
rect 159771 79732 159772 79796
rect 159836 79732 159837 79796
rect 159771 79731 159837 79732
rect 159403 79252 159469 79253
rect 159403 79188 159404 79252
rect 159468 79188 159469 79252
rect 159403 79187 159469 79188
rect 159035 78708 159101 78709
rect 159035 78644 159036 78708
rect 159100 78644 159101 78708
rect 159035 78643 159101 78644
rect 158851 78300 158917 78301
rect 158851 78236 158852 78300
rect 158916 78236 158917 78300
rect 158851 78235 158917 78236
rect 158854 31109 158914 78235
rect 158851 31108 158917 31109
rect 158851 31044 158852 31108
rect 158916 31044 158917 31108
rect 158851 31043 158917 31044
rect 159038 21453 159098 78643
rect 159774 78573 159834 79731
rect 159771 78572 159837 78573
rect 159771 78508 159772 78572
rect 159836 78508 159837 78572
rect 159771 78507 159837 78508
rect 159294 52954 159914 78000
rect 160142 77349 160202 79867
rect 160139 77348 160205 77349
rect 160139 77284 160140 77348
rect 160204 77284 160205 77348
rect 160139 77283 160205 77284
rect 159294 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 159914 52954
rect 159294 52634 159914 52718
rect 159294 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 159914 52634
rect 159035 21452 159101 21453
rect 159035 21388 159036 21452
rect 159100 21388 159101 21452
rect 159035 21387 159101 21388
rect 159294 16954 159914 52398
rect 159294 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 159914 16954
rect 159294 16634 159914 16718
rect 159294 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 159914 16634
rect 158483 10300 158549 10301
rect 158483 10236 158484 10300
rect 158548 10236 158549 10300
rect 158483 10235 158549 10236
rect 156643 9348 156709 9349
rect 156643 9284 156644 9348
rect 156708 9284 156709 9348
rect 156643 9283 156709 9284
rect 154794 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 155414 -2266
rect 154794 -2586 155414 -2502
rect 154794 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 155414 -2586
rect 154794 -7654 155414 -2822
rect 159294 -3226 159914 16398
rect 160694 9213 160754 79867
rect 160875 79796 160941 79797
rect 160875 79732 160876 79796
rect 160940 79732 160941 79796
rect 160875 79731 160941 79732
rect 160878 76533 160938 79731
rect 161982 76533 162042 79867
rect 160875 76532 160941 76533
rect 160875 76468 160876 76532
rect 160940 76468 160941 76532
rect 160875 76467 160941 76468
rect 161059 76532 161125 76533
rect 161059 76468 161060 76532
rect 161124 76468 161125 76532
rect 161059 76467 161125 76468
rect 161979 76532 162045 76533
rect 161979 76468 161980 76532
rect 162044 76468 162045 76532
rect 161979 76467 162045 76468
rect 161062 30973 161122 76467
rect 161059 30972 161125 30973
rect 161059 30908 161060 30972
rect 161124 30908 161125 30972
rect 161059 30907 161125 30908
rect 160691 9212 160757 9213
rect 160691 9148 160692 9212
rect 160756 9148 160757 9212
rect 160691 9147 160757 9148
rect 162166 6357 162226 79867
rect 162899 79796 162965 79797
rect 162899 79732 162900 79796
rect 162964 79732 162965 79796
rect 162899 79731 162965 79732
rect 162902 78709 162962 79731
rect 162899 78708 162965 78709
rect 162899 78644 162900 78708
rect 162964 78644 162965 78708
rect 162899 78643 162965 78644
rect 163270 76533 163330 79867
rect 162531 76532 162597 76533
rect 162531 76468 162532 76532
rect 162596 76468 162597 76532
rect 162531 76467 162597 76468
rect 163267 76532 163333 76533
rect 163267 76468 163268 76532
rect 163332 76468 163333 76532
rect 163267 76467 163333 76468
rect 162347 76396 162413 76397
rect 162347 76332 162348 76396
rect 162412 76332 162413 76396
rect 162347 76331 162413 76332
rect 162350 8941 162410 76331
rect 162534 9077 162594 76467
rect 163454 53141 163514 79867
rect 163635 79796 163701 79797
rect 163635 79732 163636 79796
rect 163700 79732 163701 79796
rect 163635 79731 163701 79732
rect 163451 53140 163517 53141
rect 163451 53076 163452 53140
rect 163516 53076 163517 53140
rect 163451 53075 163517 53076
rect 163638 43485 163698 79731
rect 163794 57454 164414 78000
rect 164742 75309 164802 79867
rect 165291 79796 165357 79797
rect 165291 79732 165292 79796
rect 165356 79732 165357 79796
rect 165291 79731 165357 79732
rect 164923 76532 164989 76533
rect 164923 76468 164924 76532
rect 164988 76468 164989 76532
rect 164923 76467 164989 76468
rect 164739 75308 164805 75309
rect 164739 75244 164740 75308
rect 164804 75244 164805 75308
rect 164739 75243 164805 75244
rect 164926 64157 164986 76467
rect 165107 76396 165173 76397
rect 165107 76332 165108 76396
rect 165172 76332 165173 76396
rect 165107 76331 165173 76332
rect 164923 64156 164989 64157
rect 164923 64092 164924 64156
rect 164988 64092 164989 64156
rect 164923 64091 164989 64092
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163635 43484 163701 43485
rect 163635 43420 163636 43484
rect 163700 43420 163701 43484
rect 163635 43419 163701 43420
rect 163794 21454 164414 56898
rect 165110 50285 165170 76331
rect 165107 50284 165173 50285
rect 165107 50220 165108 50284
rect 165172 50220 165173 50284
rect 165107 50219 165173 50220
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 165294 21317 165354 79731
rect 165291 21316 165357 21317
rect 165291 21252 165292 21316
rect 165356 21252 165357 21316
rect 165291 21251 165357 21252
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 162531 9076 162597 9077
rect 162531 9012 162532 9076
rect 162596 9012 162597 9076
rect 162531 9011 162597 9012
rect 162347 8940 162413 8941
rect 162347 8876 162348 8940
rect 162412 8876 162413 8940
rect 162347 8875 162413 8876
rect 162163 6356 162229 6357
rect 162163 6292 162164 6356
rect 162228 6292 162229 6356
rect 162163 6291 162229 6292
rect 159294 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 159914 -3226
rect 159294 -3546 159914 -3462
rect 159294 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 159914 -3546
rect 159294 -7654 159914 -3782
rect 163794 -4186 164414 20898
rect 165478 14517 165538 79867
rect 166214 68237 166274 79867
rect 166579 79796 166645 79797
rect 166579 79732 166580 79796
rect 166644 79732 166645 79796
rect 166579 79731 166645 79732
rect 167867 79796 167933 79797
rect 167867 79732 167868 79796
rect 167932 79732 167933 79796
rect 167867 79731 167933 79732
rect 166395 76396 166461 76397
rect 166395 76332 166396 76396
rect 166460 76332 166461 76396
rect 166395 76331 166461 76332
rect 166211 68236 166277 68237
rect 166211 68172 166212 68236
rect 166276 68172 166277 68236
rect 166211 68171 166277 68172
rect 166398 28253 166458 76331
rect 166395 28252 166461 28253
rect 166395 28188 166396 28252
rect 166460 28188 166461 28252
rect 166395 28187 166461 28188
rect 166582 24173 166642 79731
rect 166763 76532 166829 76533
rect 166763 76468 166764 76532
rect 166828 76468 166829 76532
rect 166763 76467 166829 76468
rect 167683 76532 167749 76533
rect 167683 76468 167684 76532
rect 167748 76468 167749 76532
rect 167683 76467 167749 76468
rect 166579 24172 166645 24173
rect 166579 24108 166580 24172
rect 166644 24108 166645 24172
rect 166579 24107 166645 24108
rect 165475 14516 165541 14517
rect 165475 14452 165476 14516
rect 165540 14452 165541 14516
rect 165475 14451 165541 14452
rect 166766 13021 166826 76467
rect 167686 46205 167746 76467
rect 167683 46204 167749 46205
rect 167683 46140 167684 46204
rect 167748 46140 167749 46204
rect 167683 46139 167749 46140
rect 167870 32605 167930 79731
rect 167867 32604 167933 32605
rect 167867 32540 167868 32604
rect 167932 32540 167933 32604
rect 167867 32539 167933 32540
rect 166763 13020 166829 13021
rect 166763 12956 166764 13020
rect 166828 12956 166829 13020
rect 166763 12955 166829 12956
rect 168054 6221 168114 79867
rect 168790 78437 168850 79867
rect 169339 79796 169405 79797
rect 169339 79732 169340 79796
rect 169404 79732 169405 79796
rect 169339 79731 169405 79732
rect 168787 78436 168853 78437
rect 168787 78372 168788 78436
rect 168852 78372 168853 78436
rect 168787 78371 168853 78372
rect 168294 61954 168914 78000
rect 168294 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 168914 61954
rect 168294 61634 168914 61718
rect 168294 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 168914 61634
rect 168294 25954 168914 61398
rect 169342 32469 169402 79731
rect 169526 77213 169586 79867
rect 169523 77212 169589 77213
rect 169523 77148 169524 77212
rect 169588 77148 169589 77212
rect 169523 77147 169589 77148
rect 170262 75989 170322 79867
rect 170811 79796 170877 79797
rect 170811 79732 170812 79796
rect 170876 79732 170877 79796
rect 170811 79731 170877 79732
rect 170995 79796 171061 79797
rect 170995 79732 170996 79796
rect 171060 79732 171061 79796
rect 170995 79731 171061 79732
rect 171179 79796 171245 79797
rect 171179 79732 171180 79796
rect 171244 79732 171245 79796
rect 171179 79731 171245 79732
rect 170627 76124 170693 76125
rect 170627 76060 170628 76124
rect 170692 76060 170693 76124
rect 170627 76059 170693 76060
rect 170259 75988 170325 75989
rect 170259 75924 170260 75988
rect 170324 75924 170325 75988
rect 170259 75923 170325 75924
rect 170443 75988 170509 75989
rect 170443 75924 170444 75988
rect 170508 75924 170509 75988
rect 170443 75923 170509 75924
rect 170446 62797 170506 75923
rect 170443 62796 170509 62797
rect 170443 62732 170444 62796
rect 170508 62732 170509 62796
rect 170443 62731 170509 62732
rect 170630 58581 170690 76059
rect 170627 58580 170693 58581
rect 170627 58516 170628 58580
rect 170692 58516 170693 58580
rect 170627 58515 170693 58516
rect 169339 32468 169405 32469
rect 169339 32404 169340 32468
rect 169404 32404 169405 32468
rect 169339 32403 169405 32404
rect 168294 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 168914 25954
rect 168294 25634 168914 25718
rect 168294 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 168914 25634
rect 168051 6220 168117 6221
rect 168051 6156 168052 6220
rect 168116 6156 168117 6220
rect 168051 6155 168117 6156
rect 163794 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 164414 -4186
rect 163794 -4506 164414 -4422
rect 163794 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 164414 -4506
rect 163794 -7654 164414 -4742
rect 168294 -5146 168914 25398
rect 170814 22677 170874 79731
rect 170998 77893 171058 79731
rect 171182 78981 171242 79731
rect 171179 78980 171245 78981
rect 171179 78916 171180 78980
rect 171244 78916 171245 78980
rect 171179 78915 171245 78916
rect 171366 78437 171426 79870
rect 171547 79868 171548 79932
rect 171612 79868 171613 79932
rect 171547 79867 171613 79868
rect 171731 79932 171797 79933
rect 171731 79868 171732 79932
rect 171796 79868 171797 79932
rect 171731 79867 171797 79868
rect 171363 78436 171429 78437
rect 171363 78372 171364 78436
rect 171428 78372 171429 78436
rect 171363 78371 171429 78372
rect 171734 78165 171794 79867
rect 172102 79661 172162 80142
rect 171915 79660 171981 79661
rect 171915 79596 171916 79660
rect 171980 79596 171981 79660
rect 171915 79595 171981 79596
rect 172099 79660 172165 79661
rect 172099 79596 172100 79660
rect 172164 79596 172165 79660
rect 172099 79595 172165 79596
rect 171731 78164 171797 78165
rect 171731 78100 171732 78164
rect 171796 78100 171797 78164
rect 171731 78099 171797 78100
rect 170995 77892 171061 77893
rect 170995 77828 170996 77892
rect 171060 77828 171061 77892
rect 170995 77827 171061 77828
rect 170995 77484 171061 77485
rect 170995 77420 170996 77484
rect 171060 77420 171061 77484
rect 170995 77419 171061 77420
rect 170811 22676 170877 22677
rect 170811 22612 170812 22676
rect 170876 22612 170877 22676
rect 170811 22611 170877 22612
rect 170998 4861 171058 77419
rect 170995 4860 171061 4861
rect 170995 4796 170996 4860
rect 171060 4796 171061 4860
rect 170995 4795 171061 4796
rect 171918 3501 171978 79595
rect 172286 78981 172346 80411
rect 186294 79954 186914 115398
rect 173019 79932 173085 79933
rect 173019 79868 173020 79932
rect 173084 79868 173085 79932
rect 173019 79867 173085 79868
rect 173203 79932 173269 79933
rect 173203 79868 173204 79932
rect 173268 79868 173269 79932
rect 173203 79867 173269 79868
rect 172283 78980 172349 78981
rect 172283 78916 172284 78980
rect 172348 78916 172349 78980
rect 172283 78915 172349 78916
rect 173022 78709 173082 79867
rect 173206 79117 173266 79867
rect 186294 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 186914 79954
rect 186294 79634 186914 79718
rect 186294 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 186914 79634
rect 173203 79116 173269 79117
rect 173203 79052 173204 79116
rect 173268 79052 173269 79116
rect 173203 79051 173269 79052
rect 173019 78708 173085 78709
rect 173019 78644 173020 78708
rect 173084 78644 173085 78708
rect 173019 78643 173085 78644
rect 172099 78572 172165 78573
rect 172099 78508 172100 78572
rect 172164 78508 172165 78572
rect 172099 78507 172165 78508
rect 172102 3637 172162 78507
rect 172283 77348 172349 77349
rect 172283 77284 172284 77348
rect 172348 77284 172349 77348
rect 172283 77283 172349 77284
rect 172099 3636 172165 3637
rect 172099 3572 172100 3636
rect 172164 3572 172165 3636
rect 172099 3571 172165 3572
rect 171915 3500 171981 3501
rect 171915 3436 171916 3500
rect 171980 3436 171981 3500
rect 171915 3435 171981 3436
rect 172286 3365 172346 77283
rect 172794 66454 173414 78000
rect 172794 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 173414 66454
rect 172794 66134 173414 66218
rect 172794 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 173414 66134
rect 172794 30454 173414 65898
rect 172794 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 173414 30454
rect 172794 30134 173414 30218
rect 172794 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 173414 30134
rect 172283 3364 172349 3365
rect 172283 3300 172284 3364
rect 172348 3300 172349 3364
rect 172283 3299 172349 3300
rect 168294 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 168914 -5146
rect 168294 -5466 168914 -5382
rect 168294 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 168914 -5466
rect 168294 -7654 168914 -5702
rect 172794 -6106 173414 29898
rect 172794 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 173414 -6106
rect 172794 -6426 173414 -6342
rect 172794 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 173414 -6426
rect 172794 -7654 173414 -6662
rect 177294 70954 177914 78000
rect 177294 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 177914 70954
rect 177294 70634 177914 70718
rect 177294 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 177914 70634
rect 177294 34954 177914 70398
rect 177294 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 177914 34954
rect 177294 34634 177914 34718
rect 177294 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 177914 34634
rect 177294 -7066 177914 34398
rect 177294 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 177914 -7066
rect 177294 -7386 177914 -7302
rect 177294 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 177914 -7386
rect 177294 -7654 177914 -7622
rect 181794 75454 182414 78000
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 186294 43954 186914 79398
rect 186294 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 186914 43954
rect 186294 43634 186914 43718
rect 186294 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 186914 43634
rect 186294 7954 186914 43398
rect 186294 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 186914 7954
rect 186294 7634 186914 7718
rect 186294 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 186914 7634
rect 186294 -1306 186914 7398
rect 186294 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 186914 -1306
rect 186294 -1626 186914 -1542
rect 186294 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 186914 -1626
rect 186294 -7654 186914 -1862
rect 190794 228453 191414 228484
rect 190794 228217 190826 228453
rect 191062 228217 191146 228453
rect 191382 228217 191414 228453
rect 190794 228133 191414 228217
rect 190794 227897 190826 228133
rect 191062 227897 191146 228133
rect 191382 227897 191414 228133
rect 190794 192454 191414 227897
rect 190794 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 191414 192454
rect 190794 192134 191414 192218
rect 190794 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 191414 192134
rect 190794 156454 191414 191898
rect 190794 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 191414 156454
rect 190794 156134 191414 156218
rect 190794 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 191414 156134
rect 190794 120454 191414 155898
rect 190794 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 191414 120454
rect 190794 120134 191414 120218
rect 190794 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 191414 120134
rect 190794 84454 191414 119898
rect 190794 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 191414 84454
rect 190794 84134 191414 84218
rect 190794 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 191414 84134
rect 190794 48454 191414 83898
rect 190794 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 191414 48454
rect 190794 48134 191414 48218
rect 190794 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 191414 48134
rect 190794 12454 191414 47898
rect 190794 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 191414 12454
rect 190794 12134 191414 12218
rect 190794 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 191414 12134
rect 190794 -2266 191414 11898
rect 190794 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 191414 -2266
rect 190794 -2586 191414 -2502
rect 190794 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 191414 -2586
rect 190794 -7654 191414 -2822
rect 195294 196954 195914 228484
rect 195294 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 195914 196954
rect 195294 196634 195914 196718
rect 195294 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 195914 196634
rect 195294 160954 195914 196398
rect 195294 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 195914 160954
rect 195294 160634 195914 160718
rect 195294 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 195914 160634
rect 195294 124954 195914 160398
rect 195294 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 195914 124954
rect 195294 124634 195914 124718
rect 195294 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 195914 124634
rect 195294 88954 195914 124398
rect 195294 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 195914 88954
rect 195294 88634 195914 88718
rect 195294 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 195914 88634
rect 195294 52954 195914 88398
rect 195294 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 195914 52954
rect 195294 52634 195914 52718
rect 195294 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 195914 52634
rect 195294 16954 195914 52398
rect 195294 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 195914 16954
rect 195294 16634 195914 16718
rect 195294 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 195914 16634
rect 195294 -3226 195914 16398
rect 195294 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 195914 -3226
rect 195294 -3546 195914 -3462
rect 195294 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 195914 -3546
rect 195294 -7654 195914 -3782
rect 199794 201454 200414 228484
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -4186 200414 20898
rect 199794 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 200414 -4186
rect 199794 -4506 200414 -4422
rect 199794 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 200414 -4506
rect 199794 -7654 200414 -4742
rect 204294 205954 204914 228484
rect 204294 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 204914 205954
rect 204294 205634 204914 205718
rect 204294 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 204914 205634
rect 204294 169954 204914 205398
rect 204294 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 204914 169954
rect 204294 169634 204914 169718
rect 204294 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 204914 169634
rect 204294 133954 204914 169398
rect 204294 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 204914 133954
rect 204294 133634 204914 133718
rect 204294 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 204914 133634
rect 204294 97954 204914 133398
rect 204294 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 204914 97954
rect 204294 97634 204914 97718
rect 204294 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 204914 97634
rect 204294 61954 204914 97398
rect 204294 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 204914 61954
rect 204294 61634 204914 61718
rect 204294 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 204914 61634
rect 204294 25954 204914 61398
rect 204294 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 204914 25954
rect 204294 25634 204914 25718
rect 204294 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 204914 25634
rect 204294 -5146 204914 25398
rect 204294 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 204914 -5146
rect 204294 -5466 204914 -5382
rect 204294 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 204914 -5466
rect 204294 -7654 204914 -5702
rect 208794 210454 209414 228484
rect 208794 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 209414 210454
rect 208794 210134 209414 210218
rect 208794 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 209414 210134
rect 208794 174454 209414 209898
rect 208794 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 209414 174454
rect 208794 174134 209414 174218
rect 208794 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 209414 174134
rect 208794 138454 209414 173898
rect 208794 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 209414 138454
rect 208794 138134 209414 138218
rect 208794 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 209414 138134
rect 208794 102454 209414 137898
rect 208794 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 209414 102454
rect 208794 102134 209414 102218
rect 208794 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 209414 102134
rect 208794 66454 209414 101898
rect 208794 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 209414 66454
rect 208794 66134 209414 66218
rect 208794 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 209414 66134
rect 208794 30454 209414 65898
rect 208794 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 209414 30454
rect 208794 30134 209414 30218
rect 208794 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 209414 30134
rect 208794 -6106 209414 29898
rect 208794 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 209414 -6106
rect 208794 -6426 209414 -6342
rect 208794 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 209414 -6426
rect 208794 -7654 209414 -6662
rect 213294 214954 213914 228484
rect 213294 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 213914 214954
rect 213294 214634 213914 214718
rect 213294 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 213914 214634
rect 213294 178954 213914 214398
rect 213294 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 213914 178954
rect 213294 178634 213914 178718
rect 213294 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 213914 178634
rect 213294 142954 213914 178398
rect 213294 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 213914 142954
rect 213294 142634 213914 142718
rect 213294 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 213914 142634
rect 213294 106954 213914 142398
rect 213294 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 213914 106954
rect 213294 106634 213914 106718
rect 213294 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 213914 106634
rect 213294 70954 213914 106398
rect 213294 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 213914 70954
rect 213294 70634 213914 70718
rect 213294 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 213914 70634
rect 213294 34954 213914 70398
rect 213294 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 213914 34954
rect 213294 34634 213914 34718
rect 213294 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 213914 34634
rect 213294 -7066 213914 34398
rect 213294 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 213914 -7066
rect 213294 -7386 213914 -7302
rect 213294 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 213914 -7386
rect 213294 -7654 213914 -7622
rect 217794 219454 218414 228484
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 147454 218414 182898
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 222294 223954 222914 228484
rect 222294 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 222914 223954
rect 222294 223634 222914 223718
rect 222294 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 222914 223634
rect 222294 187954 222914 223398
rect 222294 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 222914 187954
rect 222294 187634 222914 187718
rect 222294 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 222914 187634
rect 222294 151954 222914 187398
rect 222294 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 222914 151954
rect 222294 151634 222914 151718
rect 222294 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 222914 151634
rect 222294 115954 222914 151398
rect 222294 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 222914 115954
rect 222294 115634 222914 115718
rect 222294 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 222914 115634
rect 222294 79954 222914 115398
rect 222294 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 222914 79954
rect 222294 79634 222914 79718
rect 222294 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 222914 79634
rect 222294 43954 222914 79398
rect 222294 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 222914 43954
rect 222294 43634 222914 43718
rect 222294 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 222914 43634
rect 222294 7954 222914 43398
rect 222294 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 222914 7954
rect 222294 7634 222914 7718
rect 222294 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 222914 7634
rect 222294 -1306 222914 7398
rect 222294 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 222914 -1306
rect 222294 -1626 222914 -1542
rect 222294 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 222914 -1626
rect 222294 -7654 222914 -1862
rect 226794 228453 227414 228484
rect 226794 228217 226826 228453
rect 227062 228217 227146 228453
rect 227382 228217 227414 228453
rect 226794 228133 227414 228217
rect 226794 227897 226826 228133
rect 227062 227897 227146 228133
rect 227382 227897 227414 228133
rect 226794 192454 227414 227897
rect 226794 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 227414 192454
rect 226794 192134 227414 192218
rect 226794 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 227414 192134
rect 226794 156454 227414 191898
rect 226794 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 227414 156454
rect 226794 156134 227414 156218
rect 226794 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 227414 156134
rect 226794 120454 227414 155898
rect 226794 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 227414 120454
rect 226794 120134 227414 120218
rect 226794 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 227414 120134
rect 226794 84454 227414 119898
rect 226794 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 227414 84454
rect 226794 84134 227414 84218
rect 226794 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 227414 84134
rect 226794 48454 227414 83898
rect 226794 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 227414 48454
rect 226794 48134 227414 48218
rect 226794 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 227414 48134
rect 226794 12454 227414 47898
rect 226794 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 227414 12454
rect 226794 12134 227414 12218
rect 226794 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 227414 12134
rect 226794 -2266 227414 11898
rect 226794 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 227414 -2266
rect 226794 -2586 227414 -2502
rect 226794 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 227414 -2586
rect 226794 -7654 227414 -2822
rect 231294 196954 231914 228484
rect 231294 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 231914 196954
rect 231294 196634 231914 196718
rect 231294 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 231914 196634
rect 231294 160954 231914 196398
rect 231294 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 231914 160954
rect 231294 160634 231914 160718
rect 231294 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 231914 160634
rect 231294 124954 231914 160398
rect 231294 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 231914 124954
rect 231294 124634 231914 124718
rect 231294 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 231914 124634
rect 231294 88954 231914 124398
rect 231294 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 231914 88954
rect 231294 88634 231914 88718
rect 231294 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 231914 88634
rect 231294 52954 231914 88398
rect 231294 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 231914 52954
rect 231294 52634 231914 52718
rect 231294 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 231914 52634
rect 231294 16954 231914 52398
rect 231294 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 231914 16954
rect 231294 16634 231914 16718
rect 231294 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 231914 16634
rect 231294 -3226 231914 16398
rect 231294 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 231914 -3226
rect 231294 -3546 231914 -3462
rect 231294 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 231914 -3546
rect 231294 -7654 231914 -3782
rect 235794 201454 236414 228484
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 165454 236414 200898
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 235794 129454 236414 164898
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -4186 236414 20898
rect 235794 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 236414 -4186
rect 235794 -4506 236414 -4422
rect 235794 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 236414 -4506
rect 235794 -7654 236414 -4742
rect 240294 205954 240914 228484
rect 240294 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 240914 205954
rect 240294 205634 240914 205718
rect 240294 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 240914 205634
rect 240294 169954 240914 205398
rect 240294 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 240914 169954
rect 240294 169634 240914 169718
rect 240294 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 240914 169634
rect 240294 133954 240914 169398
rect 240294 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 240914 133954
rect 240294 133634 240914 133718
rect 240294 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 240914 133634
rect 240294 97954 240914 133398
rect 240294 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 240914 97954
rect 240294 97634 240914 97718
rect 240294 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 240914 97634
rect 240294 61954 240914 97398
rect 240294 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 240914 61954
rect 240294 61634 240914 61718
rect 240294 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 240914 61634
rect 240294 25954 240914 61398
rect 240294 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 240914 25954
rect 240294 25634 240914 25718
rect 240294 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 240914 25634
rect 240294 -5146 240914 25398
rect 240294 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 240914 -5146
rect 240294 -5466 240914 -5382
rect 240294 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 240914 -5466
rect 240294 -7654 240914 -5702
rect 244794 210454 245414 228484
rect 244794 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 245414 210454
rect 244794 210134 245414 210218
rect 244794 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 245414 210134
rect 244794 174454 245414 209898
rect 244794 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 245414 174454
rect 244794 174134 245414 174218
rect 244794 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 245414 174134
rect 244794 138454 245414 173898
rect 244794 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 245414 138454
rect 244794 138134 245414 138218
rect 244794 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 245414 138134
rect 244794 102454 245414 137898
rect 244794 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 245414 102454
rect 244794 102134 245414 102218
rect 244794 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 245414 102134
rect 244794 66454 245414 101898
rect 244794 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 245414 66454
rect 244794 66134 245414 66218
rect 244794 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 245414 66134
rect 244794 30454 245414 65898
rect 244794 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 245414 30454
rect 244794 30134 245414 30218
rect 244794 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 245414 30134
rect 244794 -6106 245414 29898
rect 244794 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 245414 -6106
rect 244794 -6426 245414 -6342
rect 244794 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 245414 -6426
rect 244794 -7654 245414 -6662
rect 249294 214954 249914 228484
rect 249294 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 249914 214954
rect 249294 214634 249914 214718
rect 249294 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 249914 214634
rect 249294 178954 249914 214398
rect 249294 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 249914 178954
rect 249294 178634 249914 178718
rect 249294 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 249914 178634
rect 249294 142954 249914 178398
rect 249294 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 249914 142954
rect 249294 142634 249914 142718
rect 249294 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 249914 142634
rect 249294 106954 249914 142398
rect 249294 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 249914 106954
rect 249294 106634 249914 106718
rect 249294 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 249914 106634
rect 249294 70954 249914 106398
rect 249294 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 249914 70954
rect 249294 70634 249914 70718
rect 249294 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 249914 70634
rect 249294 34954 249914 70398
rect 249294 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 249914 34954
rect 249294 34634 249914 34718
rect 249294 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 249914 34634
rect 249294 -7066 249914 34398
rect 249294 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 249914 -7066
rect 249294 -7386 249914 -7302
rect 249294 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 249914 -7386
rect 249294 -7654 249914 -7622
rect 253794 219454 254414 228484
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 258294 223954 258914 228484
rect 258294 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 258914 223954
rect 258294 223634 258914 223718
rect 258294 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 258914 223634
rect 258294 187954 258914 223398
rect 258294 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 258914 187954
rect 258294 187634 258914 187718
rect 258294 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 258914 187634
rect 258294 151954 258914 187398
rect 258294 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 258914 151954
rect 258294 151634 258914 151718
rect 258294 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 258914 151634
rect 258294 115954 258914 151398
rect 258294 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 258914 115954
rect 258294 115634 258914 115718
rect 258294 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 258914 115634
rect 258294 79954 258914 115398
rect 258294 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 258914 79954
rect 258294 79634 258914 79718
rect 258294 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 258914 79634
rect 258294 43954 258914 79398
rect 258294 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 258914 43954
rect 258294 43634 258914 43718
rect 258294 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 258914 43634
rect 258294 7954 258914 43398
rect 258294 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 258914 7954
rect 258294 7634 258914 7718
rect 258294 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 258914 7634
rect 258294 -1306 258914 7398
rect 258294 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 258914 -1306
rect 258294 -1626 258914 -1542
rect 258294 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 258914 -1626
rect 258294 -7654 258914 -1862
rect 262794 228453 263414 228484
rect 262794 228217 262826 228453
rect 263062 228217 263146 228453
rect 263382 228217 263414 228453
rect 262794 228133 263414 228217
rect 262794 227897 262826 228133
rect 263062 227897 263146 228133
rect 263382 227897 263414 228133
rect 262794 192454 263414 227897
rect 262794 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 263414 192454
rect 262794 192134 263414 192218
rect 262794 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 263414 192134
rect 262794 156454 263414 191898
rect 262794 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 263414 156454
rect 262794 156134 263414 156218
rect 262794 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 263414 156134
rect 262794 120454 263414 155898
rect 262794 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 263414 120454
rect 262794 120134 263414 120218
rect 262794 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 263414 120134
rect 262794 84454 263414 119898
rect 262794 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 263414 84454
rect 262794 84134 263414 84218
rect 262794 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 263414 84134
rect 262794 48454 263414 83898
rect 262794 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 263414 48454
rect 262794 48134 263414 48218
rect 262794 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 263414 48134
rect 262794 12454 263414 47898
rect 262794 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 263414 12454
rect 262794 12134 263414 12218
rect 262794 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 263414 12134
rect 262794 -2266 263414 11898
rect 262794 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 263414 -2266
rect 262794 -2586 263414 -2502
rect 262794 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 263414 -2586
rect 262794 -7654 263414 -2822
rect 267294 196954 267914 228484
rect 267294 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 267914 196954
rect 267294 196634 267914 196718
rect 267294 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 267914 196634
rect 267294 160954 267914 196398
rect 267294 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 267914 160954
rect 267294 160634 267914 160718
rect 267294 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 267914 160634
rect 267294 124954 267914 160398
rect 267294 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 267914 124954
rect 267294 124634 267914 124718
rect 267294 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 267914 124634
rect 267294 88954 267914 124398
rect 267294 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 267914 88954
rect 267294 88634 267914 88718
rect 267294 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 267914 88634
rect 267294 52954 267914 88398
rect 267294 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 267914 52954
rect 267294 52634 267914 52718
rect 267294 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 267914 52634
rect 267294 16954 267914 52398
rect 267294 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 267914 16954
rect 267294 16634 267914 16718
rect 267294 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 267914 16634
rect 267294 -3226 267914 16398
rect 267294 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 267914 -3226
rect 267294 -3546 267914 -3462
rect 267294 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 267914 -3546
rect 267294 -7654 267914 -3782
rect 271794 201454 272414 228484
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -4186 272414 20898
rect 271794 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 272414 -4186
rect 271794 -4506 272414 -4422
rect 271794 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 272414 -4506
rect 271794 -7654 272414 -4742
rect 276294 205954 276914 228484
rect 276294 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 276914 205954
rect 276294 205634 276914 205718
rect 276294 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 276914 205634
rect 276294 169954 276914 205398
rect 276294 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 276914 169954
rect 276294 169634 276914 169718
rect 276294 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 276914 169634
rect 276294 133954 276914 169398
rect 276294 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 276914 133954
rect 276294 133634 276914 133718
rect 276294 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 276914 133634
rect 276294 97954 276914 133398
rect 276294 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 276914 97954
rect 276294 97634 276914 97718
rect 276294 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 276914 97634
rect 276294 61954 276914 97398
rect 276294 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 276914 61954
rect 276294 61634 276914 61718
rect 276294 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 276914 61634
rect 276294 25954 276914 61398
rect 276294 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 276914 25954
rect 276294 25634 276914 25718
rect 276294 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 276914 25634
rect 276294 -5146 276914 25398
rect 276294 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 276914 -5146
rect 276294 -5466 276914 -5382
rect 276294 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 276914 -5466
rect 276294 -7654 276914 -5702
rect 280794 210454 281414 228484
rect 280794 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 281414 210454
rect 280794 210134 281414 210218
rect 280794 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 281414 210134
rect 280794 174454 281414 209898
rect 280794 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 281414 174454
rect 280794 174134 281414 174218
rect 280794 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 281414 174134
rect 280794 138454 281414 173898
rect 280794 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 281414 138454
rect 280794 138134 281414 138218
rect 280794 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 281414 138134
rect 280794 102454 281414 137898
rect 280794 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 281414 102454
rect 280794 102134 281414 102218
rect 280794 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 281414 102134
rect 280794 66454 281414 101898
rect 280794 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 281414 66454
rect 280794 66134 281414 66218
rect 280794 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 281414 66134
rect 280794 30454 281414 65898
rect 280794 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 281414 30454
rect 280794 30134 281414 30218
rect 280794 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 281414 30134
rect 280794 -6106 281414 29898
rect 280794 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 281414 -6106
rect 280794 -6426 281414 -6342
rect 280794 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 281414 -6426
rect 280794 -7654 281414 -6662
rect 285294 214954 285914 228484
rect 285294 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 285914 214954
rect 285294 214634 285914 214718
rect 285294 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 285914 214634
rect 285294 178954 285914 214398
rect 285294 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 285914 178954
rect 285294 178634 285914 178718
rect 285294 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 285914 178634
rect 285294 142954 285914 178398
rect 285294 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 285914 142954
rect 285294 142634 285914 142718
rect 285294 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 285914 142634
rect 285294 106954 285914 142398
rect 285294 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 285914 106954
rect 285294 106634 285914 106718
rect 285294 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 285914 106634
rect 285294 70954 285914 106398
rect 285294 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 285914 70954
rect 285294 70634 285914 70718
rect 285294 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 285914 70634
rect 285294 34954 285914 70398
rect 285294 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 285914 34954
rect 285294 34634 285914 34718
rect 285294 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 285914 34634
rect 285294 -7066 285914 34398
rect 285294 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 285914 -7066
rect 285294 -7386 285914 -7302
rect 285294 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 285914 -7386
rect 285294 -7654 285914 -7622
rect 289794 219454 290414 228484
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 294294 223954 294914 228484
rect 294294 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 294914 223954
rect 294294 223634 294914 223718
rect 294294 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 294914 223634
rect 294294 187954 294914 223398
rect 294294 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 294914 187954
rect 294294 187634 294914 187718
rect 294294 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 294914 187634
rect 294294 151954 294914 187398
rect 294294 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 294914 151954
rect 294294 151634 294914 151718
rect 294294 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 294914 151634
rect 294294 115954 294914 151398
rect 294294 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 294914 115954
rect 294294 115634 294914 115718
rect 294294 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 294914 115634
rect 294294 79954 294914 115398
rect 294294 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 294914 79954
rect 294294 79634 294914 79718
rect 294294 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 294914 79634
rect 294294 43954 294914 79398
rect 294294 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 294914 43954
rect 294294 43634 294914 43718
rect 294294 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 294914 43634
rect 294294 7954 294914 43398
rect 294294 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 294914 7954
rect 294294 7634 294914 7718
rect 294294 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 294914 7634
rect 294294 -1306 294914 7398
rect 294294 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 294914 -1306
rect 294294 -1626 294914 -1542
rect 294294 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 294914 -1626
rect 294294 -7654 294914 -1862
rect 298794 228453 299414 228484
rect 298794 228217 298826 228453
rect 299062 228217 299146 228453
rect 299382 228217 299414 228453
rect 298794 228133 299414 228217
rect 298794 227897 298826 228133
rect 299062 227897 299146 228133
rect 299382 227897 299414 228133
rect 298794 192454 299414 227897
rect 298794 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 299414 192454
rect 298794 192134 299414 192218
rect 298794 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 299414 192134
rect 298794 156454 299414 191898
rect 298794 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 299414 156454
rect 298794 156134 299414 156218
rect 298794 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 299414 156134
rect 298794 120454 299414 155898
rect 298794 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 299414 120454
rect 298794 120134 299414 120218
rect 298794 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 299414 120134
rect 298794 84454 299414 119898
rect 298794 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 299414 84454
rect 298794 84134 299414 84218
rect 298794 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 299414 84134
rect 298794 48454 299414 83898
rect 298794 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 299414 48454
rect 298794 48134 299414 48218
rect 298794 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 299414 48134
rect 298794 12454 299414 47898
rect 298794 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 299414 12454
rect 298794 12134 299414 12218
rect 298794 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 299414 12134
rect 298794 -2266 299414 11898
rect 298794 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 299414 -2266
rect 298794 -2586 299414 -2502
rect 298794 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 299414 -2586
rect 298794 -7654 299414 -2822
rect 303294 196954 303914 228484
rect 303294 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 303914 196954
rect 303294 196634 303914 196718
rect 303294 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 303914 196634
rect 303294 160954 303914 196398
rect 303294 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 303914 160954
rect 303294 160634 303914 160718
rect 303294 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 303914 160634
rect 303294 124954 303914 160398
rect 303294 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 303914 124954
rect 303294 124634 303914 124718
rect 303294 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 303914 124634
rect 303294 88954 303914 124398
rect 303294 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 303914 88954
rect 303294 88634 303914 88718
rect 303294 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 303914 88634
rect 303294 52954 303914 88398
rect 303294 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 303914 52954
rect 303294 52634 303914 52718
rect 303294 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 303914 52634
rect 303294 16954 303914 52398
rect 303294 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 303914 16954
rect 303294 16634 303914 16718
rect 303294 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 303914 16634
rect 303294 -3226 303914 16398
rect 303294 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 303914 -3226
rect 303294 -3546 303914 -3462
rect 303294 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 303914 -3546
rect 303294 -7654 303914 -3782
rect 307794 201454 308414 228484
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -4186 308414 20898
rect 307794 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 308414 -4186
rect 307794 -4506 308414 -4422
rect 307794 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 308414 -4506
rect 307794 -7654 308414 -4742
rect 312294 205954 312914 228484
rect 312294 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 312914 205954
rect 312294 205634 312914 205718
rect 312294 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 312914 205634
rect 312294 169954 312914 205398
rect 312294 169718 312326 169954
rect 312562 169718 312646 169954
rect 312882 169718 312914 169954
rect 312294 169634 312914 169718
rect 312294 169398 312326 169634
rect 312562 169398 312646 169634
rect 312882 169398 312914 169634
rect 312294 133954 312914 169398
rect 312294 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 312914 133954
rect 312294 133634 312914 133718
rect 312294 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 312914 133634
rect 312294 97954 312914 133398
rect 312294 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 312914 97954
rect 312294 97634 312914 97718
rect 312294 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 312914 97634
rect 312294 61954 312914 97398
rect 312294 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 312914 61954
rect 312294 61634 312914 61718
rect 312294 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 312914 61634
rect 312294 25954 312914 61398
rect 312294 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 312914 25954
rect 312294 25634 312914 25718
rect 312294 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 312914 25634
rect 312294 -5146 312914 25398
rect 312294 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 312914 -5146
rect 312294 -5466 312914 -5382
rect 312294 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 312914 -5466
rect 312294 -7654 312914 -5702
rect 316794 210454 317414 228484
rect 316794 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 317414 210454
rect 316794 210134 317414 210218
rect 316794 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 317414 210134
rect 316794 174454 317414 209898
rect 316794 174218 316826 174454
rect 317062 174218 317146 174454
rect 317382 174218 317414 174454
rect 316794 174134 317414 174218
rect 316794 173898 316826 174134
rect 317062 173898 317146 174134
rect 317382 173898 317414 174134
rect 316794 138454 317414 173898
rect 316794 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 317414 138454
rect 316794 138134 317414 138218
rect 316794 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 317414 138134
rect 316794 102454 317414 137898
rect 316794 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 317414 102454
rect 316794 102134 317414 102218
rect 316794 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 317414 102134
rect 316794 66454 317414 101898
rect 316794 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 317414 66454
rect 316794 66134 317414 66218
rect 316794 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 317414 66134
rect 316794 30454 317414 65898
rect 316794 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 317414 30454
rect 316794 30134 317414 30218
rect 316794 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 317414 30134
rect 316794 -6106 317414 29898
rect 316794 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 317414 -6106
rect 316794 -6426 317414 -6342
rect 316794 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 317414 -6426
rect 316794 -7654 317414 -6662
rect 321294 214954 321914 228484
rect 321294 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 321914 214954
rect 321294 214634 321914 214718
rect 321294 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 321914 214634
rect 321294 178954 321914 214398
rect 321294 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 321914 178954
rect 321294 178634 321914 178718
rect 321294 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 321914 178634
rect 321294 142954 321914 178398
rect 321294 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 321914 142954
rect 321294 142634 321914 142718
rect 321294 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 321914 142634
rect 321294 106954 321914 142398
rect 321294 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 321914 106954
rect 321294 106634 321914 106718
rect 321294 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 321914 106634
rect 321294 70954 321914 106398
rect 321294 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 321914 70954
rect 321294 70634 321914 70718
rect 321294 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 321914 70634
rect 321294 34954 321914 70398
rect 321294 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 321914 34954
rect 321294 34634 321914 34718
rect 321294 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 321914 34634
rect 321294 -7066 321914 34398
rect 321294 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 321914 -7066
rect 321294 -7386 321914 -7302
rect 321294 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 321914 -7386
rect 321294 -7654 321914 -7622
rect 325794 219454 326414 228484
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 330294 223954 330914 228484
rect 330294 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 330914 223954
rect 330294 223634 330914 223718
rect 330294 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 330914 223634
rect 330294 187954 330914 223398
rect 330294 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 330914 187954
rect 330294 187634 330914 187718
rect 330294 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 330914 187634
rect 330294 151954 330914 187398
rect 330294 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 330914 151954
rect 330294 151634 330914 151718
rect 330294 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 330914 151634
rect 330294 115954 330914 151398
rect 330294 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 330914 115954
rect 330294 115634 330914 115718
rect 330294 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 330914 115634
rect 330294 79954 330914 115398
rect 330294 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 330914 79954
rect 330294 79634 330914 79718
rect 330294 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 330914 79634
rect 330294 43954 330914 79398
rect 330294 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 330914 43954
rect 330294 43634 330914 43718
rect 330294 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 330914 43634
rect 330294 7954 330914 43398
rect 330294 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 330914 7954
rect 330294 7634 330914 7718
rect 330294 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 330914 7634
rect 330294 -1306 330914 7398
rect 330294 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 330914 -1306
rect 330294 -1626 330914 -1542
rect 330294 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 330914 -1626
rect 330294 -7654 330914 -1862
rect 334794 228453 335414 228484
rect 334794 228217 334826 228453
rect 335062 228217 335146 228453
rect 335382 228217 335414 228453
rect 334794 228133 335414 228217
rect 334794 227897 334826 228133
rect 335062 227897 335146 228133
rect 335382 227897 335414 228133
rect 334794 192454 335414 227897
rect 334794 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 335414 192454
rect 334794 192134 335414 192218
rect 334794 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 335414 192134
rect 334794 156454 335414 191898
rect 334794 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 335414 156454
rect 334794 156134 335414 156218
rect 334794 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 335414 156134
rect 334794 120454 335414 155898
rect 334794 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 335414 120454
rect 334794 120134 335414 120218
rect 334794 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 335414 120134
rect 334794 84454 335414 119898
rect 334794 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 335414 84454
rect 334794 84134 335414 84218
rect 334794 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 335414 84134
rect 334794 48454 335414 83898
rect 334794 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 335414 48454
rect 334794 48134 335414 48218
rect 334794 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 335414 48134
rect 334794 12454 335414 47898
rect 334794 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 335414 12454
rect 334794 12134 335414 12218
rect 334794 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 335414 12134
rect 334794 -2266 335414 11898
rect 334794 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 335414 -2266
rect 334794 -2586 335414 -2502
rect 334794 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 335414 -2586
rect 334794 -7654 335414 -2822
rect 339294 196954 339914 228484
rect 339294 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 339914 196954
rect 339294 196634 339914 196718
rect 339294 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 339914 196634
rect 339294 160954 339914 196398
rect 339294 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 339914 160954
rect 339294 160634 339914 160718
rect 339294 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 339914 160634
rect 339294 124954 339914 160398
rect 339294 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 339914 124954
rect 339294 124634 339914 124718
rect 339294 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 339914 124634
rect 339294 88954 339914 124398
rect 339294 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 339914 88954
rect 339294 88634 339914 88718
rect 339294 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 339914 88634
rect 339294 52954 339914 88398
rect 339294 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 339914 52954
rect 339294 52634 339914 52718
rect 339294 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 339914 52634
rect 339294 16954 339914 52398
rect 339294 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 339914 16954
rect 339294 16634 339914 16718
rect 339294 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 339914 16634
rect 339294 -3226 339914 16398
rect 339294 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 339914 -3226
rect 339294 -3546 339914 -3462
rect 339294 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 339914 -3546
rect 339294 -7654 339914 -3782
rect 343794 201454 344414 228484
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -4186 344414 20898
rect 343794 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 344414 -4186
rect 343794 -4506 344414 -4422
rect 343794 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 344414 -4506
rect 343794 -7654 344414 -4742
rect 348294 205954 348914 228484
rect 348294 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 348914 205954
rect 348294 205634 348914 205718
rect 348294 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 348914 205634
rect 348294 169954 348914 205398
rect 348294 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 348914 169954
rect 348294 169634 348914 169718
rect 348294 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 348914 169634
rect 348294 133954 348914 169398
rect 348294 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 348914 133954
rect 348294 133634 348914 133718
rect 348294 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 348914 133634
rect 348294 97954 348914 133398
rect 348294 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 348914 97954
rect 348294 97634 348914 97718
rect 348294 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 348914 97634
rect 348294 61954 348914 97398
rect 348294 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 348914 61954
rect 348294 61634 348914 61718
rect 348294 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 348914 61634
rect 348294 25954 348914 61398
rect 348294 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 348914 25954
rect 348294 25634 348914 25718
rect 348294 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 348914 25634
rect 348294 -5146 348914 25398
rect 348294 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 348914 -5146
rect 348294 -5466 348914 -5382
rect 348294 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 348914 -5466
rect 348294 -7654 348914 -5702
rect 352794 210454 353414 228484
rect 352794 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 353414 210454
rect 352794 210134 353414 210218
rect 352794 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 353414 210134
rect 352794 174454 353414 209898
rect 352794 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 353414 174454
rect 352794 174134 353414 174218
rect 352794 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 353414 174134
rect 352794 138454 353414 173898
rect 352794 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 353414 138454
rect 352794 138134 353414 138218
rect 352794 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 353414 138134
rect 352794 102454 353414 137898
rect 352794 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 353414 102454
rect 352794 102134 353414 102218
rect 352794 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 353414 102134
rect 352794 66454 353414 101898
rect 352794 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 353414 66454
rect 352794 66134 353414 66218
rect 352794 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 353414 66134
rect 352794 30454 353414 65898
rect 352794 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 353414 30454
rect 352794 30134 353414 30218
rect 352794 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 353414 30134
rect 352794 -6106 353414 29898
rect 352794 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 353414 -6106
rect 352794 -6426 353414 -6342
rect 352794 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 353414 -6426
rect 352794 -7654 353414 -6662
rect 357294 214954 357914 228484
rect 357294 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 357914 214954
rect 357294 214634 357914 214718
rect 357294 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 357914 214634
rect 357294 178954 357914 214398
rect 357294 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 357914 178954
rect 357294 178634 357914 178718
rect 357294 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 357914 178634
rect 357294 142954 357914 178398
rect 357294 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 357914 142954
rect 357294 142634 357914 142718
rect 357294 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 357914 142634
rect 357294 106954 357914 142398
rect 357294 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 357914 106954
rect 357294 106634 357914 106718
rect 357294 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 357914 106634
rect 357294 70954 357914 106398
rect 357294 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 357914 70954
rect 357294 70634 357914 70718
rect 357294 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 357914 70634
rect 357294 34954 357914 70398
rect 357294 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 357914 34954
rect 357294 34634 357914 34718
rect 357294 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 357914 34634
rect 357294 -7066 357914 34398
rect 357294 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 357914 -7066
rect 357294 -7386 357914 -7302
rect 357294 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 357914 -7386
rect 357294 -7654 357914 -7622
rect 361794 219454 362414 228484
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 366294 223954 366914 228484
rect 366294 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 366914 223954
rect 366294 223634 366914 223718
rect 366294 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 366914 223634
rect 366294 187954 366914 223398
rect 366294 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 366914 187954
rect 366294 187634 366914 187718
rect 366294 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 366914 187634
rect 366294 151954 366914 187398
rect 366294 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 366914 151954
rect 366294 151634 366914 151718
rect 366294 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 366914 151634
rect 366294 115954 366914 151398
rect 366294 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 366914 115954
rect 366294 115634 366914 115718
rect 366294 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 366914 115634
rect 366294 79954 366914 115398
rect 366294 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 366914 79954
rect 366294 79634 366914 79718
rect 366294 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 366914 79634
rect 366294 43954 366914 79398
rect 366294 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 366914 43954
rect 366294 43634 366914 43718
rect 366294 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 366914 43634
rect 366294 7954 366914 43398
rect 366294 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 366914 7954
rect 366294 7634 366914 7718
rect 366294 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 366914 7634
rect 366294 -1306 366914 7398
rect 366294 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 366914 -1306
rect 366294 -1626 366914 -1542
rect 366294 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 366914 -1626
rect 366294 -7654 366914 -1862
rect 370794 228453 371414 228484
rect 370794 228217 370826 228453
rect 371062 228217 371146 228453
rect 371382 228217 371414 228453
rect 370794 228133 371414 228217
rect 370794 227897 370826 228133
rect 371062 227897 371146 228133
rect 371382 227897 371414 228133
rect 370794 192454 371414 227897
rect 370794 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 371414 192454
rect 370794 192134 371414 192218
rect 370794 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 371414 192134
rect 370794 156454 371414 191898
rect 370794 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 371414 156454
rect 370794 156134 371414 156218
rect 370794 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 371414 156134
rect 370794 120454 371414 155898
rect 370794 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 371414 120454
rect 370794 120134 371414 120218
rect 370794 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 371414 120134
rect 370794 84454 371414 119898
rect 370794 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 371414 84454
rect 370794 84134 371414 84218
rect 370794 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 371414 84134
rect 370794 48454 371414 83898
rect 370794 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 371414 48454
rect 370794 48134 371414 48218
rect 370794 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 371414 48134
rect 370794 12454 371414 47898
rect 370794 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 371414 12454
rect 370794 12134 371414 12218
rect 370794 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 371414 12134
rect 370794 -2266 371414 11898
rect 370794 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 371414 -2266
rect 370794 -2586 371414 -2502
rect 370794 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 371414 -2586
rect 370794 -7654 371414 -2822
rect 375294 196954 375914 228484
rect 375294 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 375914 196954
rect 375294 196634 375914 196718
rect 375294 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 375914 196634
rect 375294 160954 375914 196398
rect 375294 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 375914 160954
rect 375294 160634 375914 160718
rect 375294 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 375914 160634
rect 375294 124954 375914 160398
rect 375294 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 375914 124954
rect 375294 124634 375914 124718
rect 375294 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 375914 124634
rect 375294 88954 375914 124398
rect 375294 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 375914 88954
rect 375294 88634 375914 88718
rect 375294 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 375914 88634
rect 375294 52954 375914 88398
rect 375294 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 375914 52954
rect 375294 52634 375914 52718
rect 375294 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 375914 52634
rect 375294 16954 375914 52398
rect 375294 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 375914 16954
rect 375294 16634 375914 16718
rect 375294 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 375914 16634
rect 375294 -3226 375914 16398
rect 375294 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 375914 -3226
rect 375294 -3546 375914 -3462
rect 375294 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 375914 -3546
rect 375294 -7654 375914 -3782
rect 379794 201454 380414 228484
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -4186 380414 20898
rect 379794 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 380414 -4186
rect 379794 -4506 380414 -4422
rect 379794 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 380414 -4506
rect 379794 -7654 380414 -4742
rect 384294 205954 384914 228484
rect 384294 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 384914 205954
rect 384294 205634 384914 205718
rect 384294 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 384914 205634
rect 384294 169954 384914 205398
rect 384294 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 384914 169954
rect 384294 169634 384914 169718
rect 384294 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 384914 169634
rect 384294 133954 384914 169398
rect 384294 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 384914 133954
rect 384294 133634 384914 133718
rect 384294 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 384914 133634
rect 384294 97954 384914 133398
rect 384294 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 384914 97954
rect 384294 97634 384914 97718
rect 384294 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 384914 97634
rect 384294 61954 384914 97398
rect 384294 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 384914 61954
rect 384294 61634 384914 61718
rect 384294 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 384914 61634
rect 384294 25954 384914 61398
rect 384294 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 384914 25954
rect 384294 25634 384914 25718
rect 384294 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 384914 25634
rect 384294 -5146 384914 25398
rect 384294 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 384914 -5146
rect 384294 -5466 384914 -5382
rect 384294 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 384914 -5466
rect 384294 -7654 384914 -5702
rect 388794 210454 389414 228484
rect 388794 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 389414 210454
rect 388794 210134 389414 210218
rect 388794 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 389414 210134
rect 388794 174454 389414 209898
rect 388794 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 389414 174454
rect 388794 174134 389414 174218
rect 388794 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 389414 174134
rect 388794 138454 389414 173898
rect 388794 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 389414 138454
rect 388794 138134 389414 138218
rect 388794 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 389414 138134
rect 388794 102454 389414 137898
rect 388794 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 389414 102454
rect 388794 102134 389414 102218
rect 388794 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 389414 102134
rect 388794 66454 389414 101898
rect 388794 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 389414 66454
rect 388794 66134 389414 66218
rect 388794 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 389414 66134
rect 388794 30454 389414 65898
rect 388794 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 389414 30454
rect 388794 30134 389414 30218
rect 388794 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 389414 30134
rect 388794 -6106 389414 29898
rect 388794 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 389414 -6106
rect 388794 -6426 389414 -6342
rect 388794 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 389414 -6426
rect 388794 -7654 389414 -6662
rect 393294 214954 393914 228484
rect 393294 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 393914 214954
rect 393294 214634 393914 214718
rect 393294 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 393914 214634
rect 393294 178954 393914 214398
rect 393294 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 393914 178954
rect 393294 178634 393914 178718
rect 393294 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 393914 178634
rect 393294 142954 393914 178398
rect 393294 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 393914 142954
rect 393294 142634 393914 142718
rect 393294 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 393914 142634
rect 393294 106954 393914 142398
rect 393294 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 393914 106954
rect 393294 106634 393914 106718
rect 393294 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 393914 106634
rect 393294 70954 393914 106398
rect 393294 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 393914 70954
rect 393294 70634 393914 70718
rect 393294 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 393914 70634
rect 393294 34954 393914 70398
rect 393294 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 393914 34954
rect 393294 34634 393914 34718
rect 393294 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 393914 34634
rect 393294 -7066 393914 34398
rect 393294 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 393914 -7066
rect 393294 -7386 393914 -7302
rect 393294 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 393914 -7386
rect 393294 -7654 393914 -7622
rect 397794 219454 398414 228484
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 402294 223954 402914 228484
rect 402294 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 402914 223954
rect 402294 223634 402914 223718
rect 402294 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 402914 223634
rect 402294 187954 402914 223398
rect 402294 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 402914 187954
rect 402294 187634 402914 187718
rect 402294 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 402914 187634
rect 402294 151954 402914 187398
rect 402294 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 402914 151954
rect 402294 151634 402914 151718
rect 402294 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 402914 151634
rect 402294 115954 402914 151398
rect 402294 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 402914 115954
rect 402294 115634 402914 115718
rect 402294 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 402914 115634
rect 402294 79954 402914 115398
rect 402294 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 402914 79954
rect 402294 79634 402914 79718
rect 402294 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 402914 79634
rect 402294 43954 402914 79398
rect 402294 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 402914 43954
rect 402294 43634 402914 43718
rect 402294 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 402914 43634
rect 402294 7954 402914 43398
rect 402294 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 402914 7954
rect 402294 7634 402914 7718
rect 402294 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 402914 7634
rect 402294 -1306 402914 7398
rect 402294 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 402914 -1306
rect 402294 -1626 402914 -1542
rect 402294 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 402914 -1626
rect 402294 -7654 402914 -1862
rect 406794 228454 407414 263898
rect 406794 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 407414 228454
rect 406794 228134 407414 228218
rect 406794 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 407414 228134
rect 406794 192454 407414 227898
rect 406794 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 407414 192454
rect 406794 192134 407414 192218
rect 406794 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 407414 192134
rect 406794 156454 407414 191898
rect 406794 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 407414 156454
rect 406794 156134 407414 156218
rect 406794 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 407414 156134
rect 406794 120454 407414 155898
rect 406794 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 407414 120454
rect 406794 120134 407414 120218
rect 406794 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 407414 120134
rect 406794 84454 407414 119898
rect 406794 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 407414 84454
rect 406794 84134 407414 84218
rect 406794 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 407414 84134
rect 406794 48454 407414 83898
rect 406794 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 407414 48454
rect 406794 48134 407414 48218
rect 406794 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 407414 48134
rect 406794 12454 407414 47898
rect 406794 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 407414 12454
rect 406794 12134 407414 12218
rect 406794 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 407414 12134
rect 406794 -2266 407414 11898
rect 406794 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 407414 -2266
rect 406794 -2586 407414 -2502
rect 406794 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 407414 -2586
rect 406794 -7654 407414 -2822
rect 411294 707718 411914 711590
rect 411294 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 411914 707718
rect 411294 707398 411914 707482
rect 411294 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 411914 707398
rect 411294 700954 411914 707162
rect 411294 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 411914 700954
rect 411294 700634 411914 700718
rect 411294 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 411914 700634
rect 411294 664954 411914 700398
rect 411294 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 411914 664954
rect 411294 664634 411914 664718
rect 411294 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 411914 664634
rect 411294 628954 411914 664398
rect 411294 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 411914 628954
rect 411294 628634 411914 628718
rect 411294 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 411914 628634
rect 411294 592954 411914 628398
rect 411294 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 411914 592954
rect 411294 592634 411914 592718
rect 411294 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 411914 592634
rect 411294 556954 411914 592398
rect 411294 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 411914 556954
rect 411294 556634 411914 556718
rect 411294 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 411914 556634
rect 411294 520954 411914 556398
rect 411294 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 411914 520954
rect 411294 520634 411914 520718
rect 411294 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 411914 520634
rect 411294 484954 411914 520398
rect 411294 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 411914 484954
rect 411294 484634 411914 484718
rect 411294 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 411914 484634
rect 411294 448954 411914 484398
rect 411294 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 411914 448954
rect 411294 448634 411914 448718
rect 411294 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 411914 448634
rect 411294 412954 411914 448398
rect 411294 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 411914 412954
rect 411294 412634 411914 412718
rect 411294 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 411914 412634
rect 411294 376954 411914 412398
rect 411294 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 411914 376954
rect 411294 376634 411914 376718
rect 411294 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 411914 376634
rect 411294 340954 411914 376398
rect 411294 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 411914 340954
rect 411294 340634 411914 340718
rect 411294 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 411914 340634
rect 411294 304954 411914 340398
rect 411294 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 411914 304954
rect 411294 304634 411914 304718
rect 411294 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 411914 304634
rect 411294 268954 411914 304398
rect 411294 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 411914 268954
rect 411294 268634 411914 268718
rect 411294 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 411914 268634
rect 411294 232954 411914 268398
rect 411294 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 411914 232954
rect 411294 232634 411914 232718
rect 411294 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 411914 232634
rect 411294 196954 411914 232398
rect 411294 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 411914 196954
rect 411294 196634 411914 196718
rect 411294 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 411914 196634
rect 411294 160954 411914 196398
rect 411294 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 411914 160954
rect 411294 160634 411914 160718
rect 411294 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 411914 160634
rect 411294 124954 411914 160398
rect 411294 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 411914 124954
rect 411294 124634 411914 124718
rect 411294 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 411914 124634
rect 411294 88954 411914 124398
rect 411294 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 411914 88954
rect 411294 88634 411914 88718
rect 411294 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 411914 88634
rect 411294 52954 411914 88398
rect 411294 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 411914 52954
rect 411294 52634 411914 52718
rect 411294 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 411914 52634
rect 411294 16954 411914 52398
rect 411294 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 411914 16954
rect 411294 16634 411914 16718
rect 411294 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 411914 16634
rect 411294 -3226 411914 16398
rect 411294 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 411914 -3226
rect 411294 -3546 411914 -3462
rect 411294 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 411914 -3546
rect 411294 -7654 411914 -3782
rect 415794 708678 416414 711590
rect 415794 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 416414 708678
rect 415794 708358 416414 708442
rect 415794 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 416414 708358
rect 415794 669454 416414 708122
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -4186 416414 20898
rect 415794 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 416414 -4186
rect 415794 -4506 416414 -4422
rect 415794 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 416414 -4506
rect 415794 -7654 416414 -4742
rect 420294 709638 420914 711590
rect 420294 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 420914 709638
rect 420294 709318 420914 709402
rect 420294 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 420914 709318
rect 420294 673954 420914 709082
rect 420294 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 420914 673954
rect 420294 673634 420914 673718
rect 420294 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 420914 673634
rect 420294 637954 420914 673398
rect 420294 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 420914 637954
rect 420294 637634 420914 637718
rect 420294 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 420914 637634
rect 420294 601954 420914 637398
rect 420294 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 420914 601954
rect 420294 601634 420914 601718
rect 420294 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 420914 601634
rect 420294 565954 420914 601398
rect 420294 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 420914 565954
rect 420294 565634 420914 565718
rect 420294 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 420914 565634
rect 420294 529954 420914 565398
rect 420294 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 420914 529954
rect 420294 529634 420914 529718
rect 420294 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 420914 529634
rect 420294 493954 420914 529398
rect 420294 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 420914 493954
rect 420294 493634 420914 493718
rect 420294 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 420914 493634
rect 420294 457954 420914 493398
rect 420294 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 420914 457954
rect 420294 457634 420914 457718
rect 420294 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 420914 457634
rect 420294 421954 420914 457398
rect 420294 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 420914 421954
rect 420294 421634 420914 421718
rect 420294 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 420914 421634
rect 420294 385954 420914 421398
rect 420294 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 420914 385954
rect 420294 385634 420914 385718
rect 420294 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 420914 385634
rect 420294 349954 420914 385398
rect 420294 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 420914 349954
rect 420294 349634 420914 349718
rect 420294 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 420914 349634
rect 420294 313954 420914 349398
rect 420294 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 420914 313954
rect 420294 313634 420914 313718
rect 420294 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 420914 313634
rect 420294 277954 420914 313398
rect 420294 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 420914 277954
rect 420294 277634 420914 277718
rect 420294 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 420914 277634
rect 420294 241954 420914 277398
rect 420294 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 420914 241954
rect 420294 241634 420914 241718
rect 420294 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 420914 241634
rect 420294 205954 420914 241398
rect 420294 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 420914 205954
rect 420294 205634 420914 205718
rect 420294 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 420914 205634
rect 420294 169954 420914 205398
rect 420294 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 420914 169954
rect 420294 169634 420914 169718
rect 420294 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 420914 169634
rect 420294 133954 420914 169398
rect 420294 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 420914 133954
rect 420294 133634 420914 133718
rect 420294 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 420914 133634
rect 420294 97954 420914 133398
rect 420294 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 420914 97954
rect 420294 97634 420914 97718
rect 420294 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 420914 97634
rect 420294 61954 420914 97398
rect 420294 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 420914 61954
rect 420294 61634 420914 61718
rect 420294 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 420914 61634
rect 420294 25954 420914 61398
rect 420294 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 420914 25954
rect 420294 25634 420914 25718
rect 420294 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 420914 25634
rect 420294 -5146 420914 25398
rect 420294 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 420914 -5146
rect 420294 -5466 420914 -5382
rect 420294 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 420914 -5466
rect 420294 -7654 420914 -5702
rect 424794 710598 425414 711590
rect 424794 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 425414 710598
rect 424794 710278 425414 710362
rect 424794 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 425414 710278
rect 424794 678454 425414 710042
rect 424794 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 425414 678454
rect 424794 678134 425414 678218
rect 424794 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 425414 678134
rect 424794 642454 425414 677898
rect 424794 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 425414 642454
rect 424794 642134 425414 642218
rect 424794 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 425414 642134
rect 424794 606454 425414 641898
rect 424794 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 425414 606454
rect 424794 606134 425414 606218
rect 424794 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 425414 606134
rect 424794 570454 425414 605898
rect 424794 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 425414 570454
rect 424794 570134 425414 570218
rect 424794 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 425414 570134
rect 424794 534454 425414 569898
rect 424794 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 425414 534454
rect 424794 534134 425414 534218
rect 424794 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 425414 534134
rect 424794 498454 425414 533898
rect 424794 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 425414 498454
rect 424794 498134 425414 498218
rect 424794 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 425414 498134
rect 424794 462454 425414 497898
rect 424794 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 425414 462454
rect 424794 462134 425414 462218
rect 424794 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 425414 462134
rect 424794 426454 425414 461898
rect 424794 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 425414 426454
rect 424794 426134 425414 426218
rect 424794 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 425414 426134
rect 424794 390454 425414 425898
rect 424794 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 425414 390454
rect 424794 390134 425414 390218
rect 424794 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 425414 390134
rect 424794 354454 425414 389898
rect 424794 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 425414 354454
rect 424794 354134 425414 354218
rect 424794 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 425414 354134
rect 424794 318454 425414 353898
rect 424794 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 425414 318454
rect 424794 318134 425414 318218
rect 424794 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 425414 318134
rect 424794 282454 425414 317898
rect 424794 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 425414 282454
rect 424794 282134 425414 282218
rect 424794 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 425414 282134
rect 424794 246454 425414 281898
rect 424794 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 425414 246454
rect 424794 246134 425414 246218
rect 424794 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 425414 246134
rect 424794 210454 425414 245898
rect 424794 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 425414 210454
rect 424794 210134 425414 210218
rect 424794 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 425414 210134
rect 424794 174454 425414 209898
rect 424794 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 425414 174454
rect 424794 174134 425414 174218
rect 424794 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 425414 174134
rect 424794 138454 425414 173898
rect 424794 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 425414 138454
rect 424794 138134 425414 138218
rect 424794 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 425414 138134
rect 424794 102454 425414 137898
rect 424794 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 425414 102454
rect 424794 102134 425414 102218
rect 424794 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 425414 102134
rect 424794 66454 425414 101898
rect 424794 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 425414 66454
rect 424794 66134 425414 66218
rect 424794 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 425414 66134
rect 424794 30454 425414 65898
rect 424794 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 425414 30454
rect 424794 30134 425414 30218
rect 424794 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 425414 30134
rect 424794 -6106 425414 29898
rect 424794 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 425414 -6106
rect 424794 -6426 425414 -6342
rect 424794 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 425414 -6426
rect 424794 -7654 425414 -6662
rect 429294 711558 429914 711590
rect 429294 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 429914 711558
rect 429294 711238 429914 711322
rect 429294 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 429914 711238
rect 429294 682954 429914 711002
rect 429294 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 429914 682954
rect 429294 682634 429914 682718
rect 429294 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 429914 682634
rect 429294 646954 429914 682398
rect 429294 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 429914 646954
rect 429294 646634 429914 646718
rect 429294 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 429914 646634
rect 429294 610954 429914 646398
rect 429294 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 429914 610954
rect 429294 610634 429914 610718
rect 429294 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 429914 610634
rect 429294 574954 429914 610398
rect 429294 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 429914 574954
rect 429294 574634 429914 574718
rect 429294 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 429914 574634
rect 429294 538954 429914 574398
rect 429294 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 429914 538954
rect 429294 538634 429914 538718
rect 429294 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 429914 538634
rect 429294 502954 429914 538398
rect 429294 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 429914 502954
rect 429294 502634 429914 502718
rect 429294 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 429914 502634
rect 429294 466954 429914 502398
rect 429294 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 429914 466954
rect 429294 466634 429914 466718
rect 429294 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 429914 466634
rect 429294 430954 429914 466398
rect 429294 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 429914 430954
rect 429294 430634 429914 430718
rect 429294 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 429914 430634
rect 429294 394954 429914 430398
rect 429294 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 429914 394954
rect 429294 394634 429914 394718
rect 429294 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 429914 394634
rect 429294 358954 429914 394398
rect 429294 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 429914 358954
rect 429294 358634 429914 358718
rect 429294 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 429914 358634
rect 429294 322954 429914 358398
rect 429294 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 429914 322954
rect 429294 322634 429914 322718
rect 429294 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 429914 322634
rect 429294 286954 429914 322398
rect 429294 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 429914 286954
rect 429294 286634 429914 286718
rect 429294 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 429914 286634
rect 429294 250954 429914 286398
rect 429294 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 429914 250954
rect 429294 250634 429914 250718
rect 429294 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 429914 250634
rect 429294 214954 429914 250398
rect 429294 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 429914 214954
rect 429294 214634 429914 214718
rect 429294 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 429914 214634
rect 429294 178954 429914 214398
rect 429294 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 429914 178954
rect 429294 178634 429914 178718
rect 429294 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 429914 178634
rect 429294 142954 429914 178398
rect 429294 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 429914 142954
rect 429294 142634 429914 142718
rect 429294 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 429914 142634
rect 429294 106954 429914 142398
rect 429294 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 429914 106954
rect 429294 106634 429914 106718
rect 429294 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 429914 106634
rect 429294 70954 429914 106398
rect 429294 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 429914 70954
rect 429294 70634 429914 70718
rect 429294 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 429914 70634
rect 429294 34954 429914 70398
rect 429294 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 429914 34954
rect 429294 34634 429914 34718
rect 429294 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 429914 34634
rect 429294 -7066 429914 34398
rect 429294 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 429914 -7066
rect 429294 -7386 429914 -7302
rect 429294 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 429914 -7386
rect 429294 -7654 429914 -7622
rect 433794 704838 434414 711590
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 438294 705798 438914 711590
rect 438294 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 438914 705798
rect 438294 705478 438914 705562
rect 438294 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 438914 705478
rect 438294 691954 438914 705242
rect 438294 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 438914 691954
rect 438294 691634 438914 691718
rect 438294 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 438914 691634
rect 438294 655954 438914 691398
rect 438294 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 438914 655954
rect 438294 655634 438914 655718
rect 438294 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 438914 655634
rect 438294 619954 438914 655398
rect 438294 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 438914 619954
rect 438294 619634 438914 619718
rect 438294 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 438914 619634
rect 438294 583954 438914 619398
rect 438294 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 438914 583954
rect 438294 583634 438914 583718
rect 438294 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 438914 583634
rect 438294 547954 438914 583398
rect 438294 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 438914 547954
rect 438294 547634 438914 547718
rect 438294 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 438914 547634
rect 438294 511954 438914 547398
rect 438294 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 438914 511954
rect 438294 511634 438914 511718
rect 438294 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 438914 511634
rect 438294 475954 438914 511398
rect 438294 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 438914 475954
rect 438294 475634 438914 475718
rect 438294 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 438914 475634
rect 438294 439954 438914 475398
rect 438294 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 438914 439954
rect 438294 439634 438914 439718
rect 438294 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 438914 439634
rect 438294 403954 438914 439398
rect 438294 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 438914 403954
rect 438294 403634 438914 403718
rect 438294 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 438914 403634
rect 438294 367954 438914 403398
rect 438294 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 438914 367954
rect 438294 367634 438914 367718
rect 438294 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 438914 367634
rect 438294 331954 438914 367398
rect 438294 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 438914 331954
rect 438294 331634 438914 331718
rect 438294 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 438914 331634
rect 438294 295954 438914 331398
rect 438294 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 438914 295954
rect 438294 295634 438914 295718
rect 438294 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 438914 295634
rect 438294 259954 438914 295398
rect 438294 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 438914 259954
rect 438294 259634 438914 259718
rect 438294 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 438914 259634
rect 438294 223954 438914 259398
rect 438294 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 438914 223954
rect 438294 223634 438914 223718
rect 438294 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 438914 223634
rect 438294 187954 438914 223398
rect 438294 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 438914 187954
rect 438294 187634 438914 187718
rect 438294 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 438914 187634
rect 438294 151954 438914 187398
rect 438294 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 438914 151954
rect 438294 151634 438914 151718
rect 438294 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 438914 151634
rect 438294 115954 438914 151398
rect 438294 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 438914 115954
rect 438294 115634 438914 115718
rect 438294 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 438914 115634
rect 438294 79954 438914 115398
rect 438294 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 438914 79954
rect 438294 79634 438914 79718
rect 438294 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 438914 79634
rect 438294 43954 438914 79398
rect 438294 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 438914 43954
rect 438294 43634 438914 43718
rect 438294 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 438914 43634
rect 438294 7954 438914 43398
rect 438294 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 438914 7954
rect 438294 7634 438914 7718
rect 438294 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 438914 7634
rect 438294 -1306 438914 7398
rect 438294 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 438914 -1306
rect 438294 -1626 438914 -1542
rect 438294 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 438914 -1626
rect 438294 -7654 438914 -1862
rect 442794 706758 443414 711590
rect 442794 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 443414 706758
rect 442794 706438 443414 706522
rect 442794 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 443414 706438
rect 442794 696454 443414 706202
rect 442794 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 443414 696454
rect 442794 696134 443414 696218
rect 442794 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 443414 696134
rect 442794 660454 443414 695898
rect 442794 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 443414 660454
rect 442794 660134 443414 660218
rect 442794 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 443414 660134
rect 442794 624454 443414 659898
rect 442794 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 443414 624454
rect 442794 624134 443414 624218
rect 442794 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 443414 624134
rect 442794 588454 443414 623898
rect 442794 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 443414 588454
rect 442794 588134 443414 588218
rect 442794 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 443414 588134
rect 442794 552454 443414 587898
rect 442794 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 443414 552454
rect 442794 552134 443414 552218
rect 442794 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 443414 552134
rect 442794 516454 443414 551898
rect 442794 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 443414 516454
rect 442794 516134 443414 516218
rect 442794 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 443414 516134
rect 442794 480454 443414 515898
rect 442794 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 443414 480454
rect 442794 480134 443414 480218
rect 442794 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 443414 480134
rect 442794 444454 443414 479898
rect 442794 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 443414 444454
rect 442794 444134 443414 444218
rect 442794 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 443414 444134
rect 442794 408454 443414 443898
rect 442794 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 443414 408454
rect 442794 408134 443414 408218
rect 442794 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 443414 408134
rect 442794 372454 443414 407898
rect 442794 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 443414 372454
rect 442794 372134 443414 372218
rect 442794 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 443414 372134
rect 442794 336454 443414 371898
rect 442794 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 443414 336454
rect 442794 336134 443414 336218
rect 442794 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 443414 336134
rect 442794 300454 443414 335898
rect 442794 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 443414 300454
rect 442794 300134 443414 300218
rect 442794 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 443414 300134
rect 442794 264454 443414 299898
rect 442794 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 443414 264454
rect 442794 264134 443414 264218
rect 442794 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 443414 264134
rect 442794 228454 443414 263898
rect 442794 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 443414 228454
rect 442794 228134 443414 228218
rect 442794 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 443414 228134
rect 442794 192454 443414 227898
rect 442794 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 443414 192454
rect 442794 192134 443414 192218
rect 442794 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 443414 192134
rect 442794 156454 443414 191898
rect 442794 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 443414 156454
rect 442794 156134 443414 156218
rect 442794 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 443414 156134
rect 442794 120454 443414 155898
rect 442794 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 443414 120454
rect 442794 120134 443414 120218
rect 442794 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 443414 120134
rect 442794 84454 443414 119898
rect 442794 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 443414 84454
rect 442794 84134 443414 84218
rect 442794 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 443414 84134
rect 442794 48454 443414 83898
rect 442794 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 443414 48454
rect 442794 48134 443414 48218
rect 442794 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 443414 48134
rect 442794 12454 443414 47898
rect 442794 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 443414 12454
rect 442794 12134 443414 12218
rect 442794 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 443414 12134
rect 442794 -2266 443414 11898
rect 442794 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 443414 -2266
rect 442794 -2586 443414 -2502
rect 442794 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 443414 -2586
rect 442794 -7654 443414 -2822
rect 447294 707718 447914 711590
rect 447294 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 447914 707718
rect 447294 707398 447914 707482
rect 447294 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 447914 707398
rect 447294 700954 447914 707162
rect 447294 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 447914 700954
rect 447294 700634 447914 700718
rect 447294 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 447914 700634
rect 447294 664954 447914 700398
rect 447294 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 447914 664954
rect 447294 664634 447914 664718
rect 447294 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 447914 664634
rect 447294 628954 447914 664398
rect 447294 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 447914 628954
rect 447294 628634 447914 628718
rect 447294 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 447914 628634
rect 447294 592954 447914 628398
rect 447294 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 447914 592954
rect 447294 592634 447914 592718
rect 447294 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 447914 592634
rect 447294 556954 447914 592398
rect 447294 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 447914 556954
rect 447294 556634 447914 556718
rect 447294 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 447914 556634
rect 447294 520954 447914 556398
rect 447294 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 447914 520954
rect 447294 520634 447914 520718
rect 447294 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 447914 520634
rect 447294 484954 447914 520398
rect 447294 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 447914 484954
rect 447294 484634 447914 484718
rect 447294 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 447914 484634
rect 447294 448954 447914 484398
rect 447294 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 447914 448954
rect 447294 448634 447914 448718
rect 447294 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 447914 448634
rect 447294 412954 447914 448398
rect 447294 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 447914 412954
rect 447294 412634 447914 412718
rect 447294 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 447914 412634
rect 447294 376954 447914 412398
rect 447294 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 447914 376954
rect 447294 376634 447914 376718
rect 447294 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 447914 376634
rect 447294 340954 447914 376398
rect 447294 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 447914 340954
rect 447294 340634 447914 340718
rect 447294 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 447914 340634
rect 447294 304954 447914 340398
rect 447294 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 447914 304954
rect 447294 304634 447914 304718
rect 447294 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 447914 304634
rect 447294 268954 447914 304398
rect 447294 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 447914 268954
rect 447294 268634 447914 268718
rect 447294 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 447914 268634
rect 447294 232954 447914 268398
rect 447294 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 447914 232954
rect 447294 232634 447914 232718
rect 447294 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 447914 232634
rect 447294 196954 447914 232398
rect 447294 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 447914 196954
rect 447294 196634 447914 196718
rect 447294 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 447914 196634
rect 447294 160954 447914 196398
rect 447294 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 447914 160954
rect 447294 160634 447914 160718
rect 447294 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 447914 160634
rect 447294 124954 447914 160398
rect 447294 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 447914 124954
rect 447294 124634 447914 124718
rect 447294 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 447914 124634
rect 447294 88954 447914 124398
rect 447294 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 447914 88954
rect 447294 88634 447914 88718
rect 447294 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 447914 88634
rect 447294 52954 447914 88398
rect 447294 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 447914 52954
rect 447294 52634 447914 52718
rect 447294 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 447914 52634
rect 447294 16954 447914 52398
rect 447294 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 447914 16954
rect 447294 16634 447914 16718
rect 447294 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 447914 16634
rect 447294 -3226 447914 16398
rect 447294 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 447914 -3226
rect 447294 -3546 447914 -3462
rect 447294 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 447914 -3546
rect 447294 -7654 447914 -3782
rect 451794 708678 452414 711590
rect 451794 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 452414 708678
rect 451794 708358 452414 708442
rect 451794 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 452414 708358
rect 451794 669454 452414 708122
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -4186 452414 20898
rect 451794 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 452414 -4186
rect 451794 -4506 452414 -4422
rect 451794 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 452414 -4506
rect 451794 -7654 452414 -4742
rect 456294 709638 456914 711590
rect 456294 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 456914 709638
rect 456294 709318 456914 709402
rect 456294 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 456914 709318
rect 456294 673954 456914 709082
rect 456294 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 456914 673954
rect 456294 673634 456914 673718
rect 456294 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 456914 673634
rect 456294 637954 456914 673398
rect 456294 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 456914 637954
rect 456294 637634 456914 637718
rect 456294 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 456914 637634
rect 456294 601954 456914 637398
rect 456294 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 456914 601954
rect 456294 601634 456914 601718
rect 456294 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 456914 601634
rect 456294 565954 456914 601398
rect 456294 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 456914 565954
rect 456294 565634 456914 565718
rect 456294 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 456914 565634
rect 456294 529954 456914 565398
rect 456294 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 456914 529954
rect 456294 529634 456914 529718
rect 456294 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 456914 529634
rect 456294 493954 456914 529398
rect 456294 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 456914 493954
rect 456294 493634 456914 493718
rect 456294 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 456914 493634
rect 456294 457954 456914 493398
rect 456294 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 456914 457954
rect 456294 457634 456914 457718
rect 456294 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 456914 457634
rect 456294 421954 456914 457398
rect 456294 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 456914 421954
rect 456294 421634 456914 421718
rect 456294 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 456914 421634
rect 456294 385954 456914 421398
rect 456294 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 456914 385954
rect 456294 385634 456914 385718
rect 456294 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 456914 385634
rect 456294 349954 456914 385398
rect 456294 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 456914 349954
rect 456294 349634 456914 349718
rect 456294 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 456914 349634
rect 456294 313954 456914 349398
rect 456294 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 456914 313954
rect 456294 313634 456914 313718
rect 456294 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 456914 313634
rect 456294 277954 456914 313398
rect 456294 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 456914 277954
rect 456294 277634 456914 277718
rect 456294 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 456914 277634
rect 456294 241954 456914 277398
rect 456294 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 456914 241954
rect 456294 241634 456914 241718
rect 456294 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 456914 241634
rect 456294 205954 456914 241398
rect 456294 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 456914 205954
rect 456294 205634 456914 205718
rect 456294 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 456914 205634
rect 456294 169954 456914 205398
rect 456294 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 456914 169954
rect 456294 169634 456914 169718
rect 456294 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 456914 169634
rect 456294 133954 456914 169398
rect 456294 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 456914 133954
rect 456294 133634 456914 133718
rect 456294 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 456914 133634
rect 456294 97954 456914 133398
rect 456294 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 456914 97954
rect 456294 97634 456914 97718
rect 456294 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 456914 97634
rect 456294 61954 456914 97398
rect 456294 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 456914 61954
rect 456294 61634 456914 61718
rect 456294 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 456914 61634
rect 456294 25954 456914 61398
rect 456294 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 456914 25954
rect 456294 25634 456914 25718
rect 456294 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 456914 25634
rect 456294 -5146 456914 25398
rect 456294 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 456914 -5146
rect 456294 -5466 456914 -5382
rect 456294 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 456914 -5466
rect 456294 -7654 456914 -5702
rect 460794 710598 461414 711590
rect 460794 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 461414 710598
rect 460794 710278 461414 710362
rect 460794 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 461414 710278
rect 460794 678454 461414 710042
rect 460794 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 461414 678454
rect 460794 678134 461414 678218
rect 460794 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 461414 678134
rect 460794 642454 461414 677898
rect 460794 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 461414 642454
rect 460794 642134 461414 642218
rect 460794 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 461414 642134
rect 460794 606454 461414 641898
rect 460794 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 461414 606454
rect 460794 606134 461414 606218
rect 460794 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 461414 606134
rect 460794 570454 461414 605898
rect 460794 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 461414 570454
rect 460794 570134 461414 570218
rect 460794 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 461414 570134
rect 460794 534454 461414 569898
rect 460794 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 461414 534454
rect 460794 534134 461414 534218
rect 460794 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 461414 534134
rect 460794 498454 461414 533898
rect 460794 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 461414 498454
rect 460794 498134 461414 498218
rect 460794 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 461414 498134
rect 460794 462454 461414 497898
rect 460794 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 461414 462454
rect 460794 462134 461414 462218
rect 460794 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 461414 462134
rect 460794 426454 461414 461898
rect 460794 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 461414 426454
rect 460794 426134 461414 426218
rect 460794 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 461414 426134
rect 460794 390454 461414 425898
rect 460794 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 461414 390454
rect 460794 390134 461414 390218
rect 460794 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 461414 390134
rect 460794 354454 461414 389898
rect 460794 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 461414 354454
rect 460794 354134 461414 354218
rect 460794 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 461414 354134
rect 460794 318454 461414 353898
rect 460794 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 461414 318454
rect 460794 318134 461414 318218
rect 460794 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 461414 318134
rect 460794 282454 461414 317898
rect 460794 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 461414 282454
rect 460794 282134 461414 282218
rect 460794 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 461414 282134
rect 460794 246454 461414 281898
rect 460794 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 461414 246454
rect 460794 246134 461414 246218
rect 460794 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 461414 246134
rect 460794 210454 461414 245898
rect 460794 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 461414 210454
rect 460794 210134 461414 210218
rect 460794 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 461414 210134
rect 460794 174454 461414 209898
rect 460794 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 461414 174454
rect 460794 174134 461414 174218
rect 460794 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 461414 174134
rect 460794 138454 461414 173898
rect 460794 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 461414 138454
rect 460794 138134 461414 138218
rect 460794 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 461414 138134
rect 460794 102454 461414 137898
rect 460794 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 461414 102454
rect 460794 102134 461414 102218
rect 460794 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 461414 102134
rect 460794 66454 461414 101898
rect 460794 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 461414 66454
rect 460794 66134 461414 66218
rect 460794 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 461414 66134
rect 460794 30454 461414 65898
rect 460794 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 461414 30454
rect 460794 30134 461414 30218
rect 460794 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 461414 30134
rect 460794 -6106 461414 29898
rect 460794 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 461414 -6106
rect 460794 -6426 461414 -6342
rect 460794 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 461414 -6426
rect 460794 -7654 461414 -6662
rect 465294 711558 465914 711590
rect 465294 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 465914 711558
rect 465294 711238 465914 711322
rect 465294 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 465914 711238
rect 465294 682954 465914 711002
rect 465294 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 465914 682954
rect 465294 682634 465914 682718
rect 465294 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 465914 682634
rect 465294 646954 465914 682398
rect 465294 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 465914 646954
rect 465294 646634 465914 646718
rect 465294 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 465914 646634
rect 465294 610954 465914 646398
rect 465294 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 465914 610954
rect 465294 610634 465914 610718
rect 465294 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 465914 610634
rect 465294 574954 465914 610398
rect 465294 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 465914 574954
rect 465294 574634 465914 574718
rect 465294 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 465914 574634
rect 465294 538954 465914 574398
rect 465294 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 465914 538954
rect 465294 538634 465914 538718
rect 465294 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 465914 538634
rect 465294 502954 465914 538398
rect 465294 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 465914 502954
rect 465294 502634 465914 502718
rect 465294 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 465914 502634
rect 465294 466954 465914 502398
rect 465294 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 465914 466954
rect 465294 466634 465914 466718
rect 465294 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 465914 466634
rect 465294 430954 465914 466398
rect 465294 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 465914 430954
rect 465294 430634 465914 430718
rect 465294 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 465914 430634
rect 465294 394954 465914 430398
rect 465294 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 465914 394954
rect 465294 394634 465914 394718
rect 465294 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 465914 394634
rect 465294 358954 465914 394398
rect 465294 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 465914 358954
rect 465294 358634 465914 358718
rect 465294 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 465914 358634
rect 465294 322954 465914 358398
rect 465294 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 465914 322954
rect 465294 322634 465914 322718
rect 465294 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 465914 322634
rect 465294 286954 465914 322398
rect 465294 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 465914 286954
rect 465294 286634 465914 286718
rect 465294 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 465914 286634
rect 465294 250954 465914 286398
rect 465294 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 465914 250954
rect 465294 250634 465914 250718
rect 465294 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 465914 250634
rect 465294 214954 465914 250398
rect 465294 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 465914 214954
rect 465294 214634 465914 214718
rect 465294 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 465914 214634
rect 465294 178954 465914 214398
rect 465294 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 465914 178954
rect 465294 178634 465914 178718
rect 465294 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 465914 178634
rect 465294 142954 465914 178398
rect 465294 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 465914 142954
rect 465294 142634 465914 142718
rect 465294 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 465914 142634
rect 465294 106954 465914 142398
rect 465294 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 465914 106954
rect 465294 106634 465914 106718
rect 465294 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 465914 106634
rect 465294 70954 465914 106398
rect 465294 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 465914 70954
rect 465294 70634 465914 70718
rect 465294 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 465914 70634
rect 465294 34954 465914 70398
rect 465294 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 465914 34954
rect 465294 34634 465914 34718
rect 465294 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 465914 34634
rect 465294 -7066 465914 34398
rect 465294 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 465914 -7066
rect 465294 -7386 465914 -7302
rect 465294 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 465914 -7386
rect 465294 -7654 465914 -7622
rect 469794 704838 470414 711590
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 474294 705798 474914 711590
rect 474294 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 474914 705798
rect 474294 705478 474914 705562
rect 474294 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 474914 705478
rect 474294 691954 474914 705242
rect 474294 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 474914 691954
rect 474294 691634 474914 691718
rect 474294 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 474914 691634
rect 474294 655954 474914 691398
rect 474294 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 474914 655954
rect 474294 655634 474914 655718
rect 474294 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 474914 655634
rect 474294 619954 474914 655398
rect 474294 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 474914 619954
rect 474294 619634 474914 619718
rect 474294 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 474914 619634
rect 474294 583954 474914 619398
rect 474294 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 474914 583954
rect 474294 583634 474914 583718
rect 474294 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 474914 583634
rect 474294 547954 474914 583398
rect 474294 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 474914 547954
rect 474294 547634 474914 547718
rect 474294 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 474914 547634
rect 474294 511954 474914 547398
rect 474294 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 474914 511954
rect 474294 511634 474914 511718
rect 474294 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 474914 511634
rect 474294 475954 474914 511398
rect 474294 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 474914 475954
rect 474294 475634 474914 475718
rect 474294 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 474914 475634
rect 474294 439954 474914 475398
rect 474294 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 474914 439954
rect 474294 439634 474914 439718
rect 474294 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 474914 439634
rect 474294 403954 474914 439398
rect 474294 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 474914 403954
rect 474294 403634 474914 403718
rect 474294 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 474914 403634
rect 474294 367954 474914 403398
rect 474294 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 474914 367954
rect 474294 367634 474914 367718
rect 474294 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 474914 367634
rect 474294 331954 474914 367398
rect 474294 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 474914 331954
rect 474294 331634 474914 331718
rect 474294 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 474914 331634
rect 474294 295954 474914 331398
rect 474294 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 474914 295954
rect 474294 295634 474914 295718
rect 474294 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 474914 295634
rect 474294 259954 474914 295398
rect 474294 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 474914 259954
rect 474294 259634 474914 259718
rect 474294 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 474914 259634
rect 474294 223954 474914 259398
rect 474294 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 474914 223954
rect 474294 223634 474914 223718
rect 474294 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 474914 223634
rect 474294 187954 474914 223398
rect 474294 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 474914 187954
rect 474294 187634 474914 187718
rect 474294 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 474914 187634
rect 474294 151954 474914 187398
rect 474294 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 474914 151954
rect 474294 151634 474914 151718
rect 474294 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 474914 151634
rect 474294 115954 474914 151398
rect 474294 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 474914 115954
rect 474294 115634 474914 115718
rect 474294 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 474914 115634
rect 474294 79954 474914 115398
rect 474294 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 474914 79954
rect 474294 79634 474914 79718
rect 474294 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 474914 79634
rect 474294 43954 474914 79398
rect 474294 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 474914 43954
rect 474294 43634 474914 43718
rect 474294 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 474914 43634
rect 474294 7954 474914 43398
rect 474294 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 474914 7954
rect 474294 7634 474914 7718
rect 474294 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 474914 7634
rect 474294 -1306 474914 7398
rect 474294 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 474914 -1306
rect 474294 -1626 474914 -1542
rect 474294 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 474914 -1626
rect 474294 -7654 474914 -1862
rect 478794 706758 479414 711590
rect 478794 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 479414 706758
rect 478794 706438 479414 706522
rect 478794 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 479414 706438
rect 478794 696454 479414 706202
rect 478794 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 479414 696454
rect 478794 696134 479414 696218
rect 478794 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 479414 696134
rect 478794 660454 479414 695898
rect 478794 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 479414 660454
rect 478794 660134 479414 660218
rect 478794 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 479414 660134
rect 478794 624454 479414 659898
rect 478794 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 479414 624454
rect 478794 624134 479414 624218
rect 478794 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 479414 624134
rect 478794 588454 479414 623898
rect 478794 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 479414 588454
rect 478794 588134 479414 588218
rect 478794 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 479414 588134
rect 478794 552454 479414 587898
rect 478794 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 479414 552454
rect 478794 552134 479414 552218
rect 478794 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 479414 552134
rect 478794 516454 479414 551898
rect 478794 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 479414 516454
rect 478794 516134 479414 516218
rect 478794 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 479414 516134
rect 478794 480454 479414 515898
rect 478794 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 479414 480454
rect 478794 480134 479414 480218
rect 478794 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 479414 480134
rect 478794 444454 479414 479898
rect 478794 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 479414 444454
rect 478794 444134 479414 444218
rect 478794 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 479414 444134
rect 478794 408454 479414 443898
rect 478794 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 479414 408454
rect 478794 408134 479414 408218
rect 478794 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 479414 408134
rect 478794 372454 479414 407898
rect 478794 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 479414 372454
rect 478794 372134 479414 372218
rect 478794 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 479414 372134
rect 478794 336454 479414 371898
rect 478794 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 479414 336454
rect 478794 336134 479414 336218
rect 478794 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 479414 336134
rect 478794 300454 479414 335898
rect 478794 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 479414 300454
rect 478794 300134 479414 300218
rect 478794 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 479414 300134
rect 478794 264454 479414 299898
rect 478794 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 479414 264454
rect 478794 264134 479414 264218
rect 478794 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 479414 264134
rect 478794 228454 479414 263898
rect 478794 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 479414 228454
rect 478794 228134 479414 228218
rect 478794 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 479414 228134
rect 478794 192454 479414 227898
rect 478794 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 479414 192454
rect 478794 192134 479414 192218
rect 478794 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 479414 192134
rect 478794 156454 479414 191898
rect 478794 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 479414 156454
rect 478794 156134 479414 156218
rect 478794 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 479414 156134
rect 478794 120454 479414 155898
rect 478794 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 479414 120454
rect 478794 120134 479414 120218
rect 478794 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 479414 120134
rect 478794 84454 479414 119898
rect 478794 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 479414 84454
rect 478794 84134 479414 84218
rect 478794 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 479414 84134
rect 478794 48454 479414 83898
rect 478794 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 479414 48454
rect 478794 48134 479414 48218
rect 478794 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 479414 48134
rect 478794 12454 479414 47898
rect 478794 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 479414 12454
rect 478794 12134 479414 12218
rect 478794 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 479414 12134
rect 478794 -2266 479414 11898
rect 478794 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 479414 -2266
rect 478794 -2586 479414 -2502
rect 478794 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 479414 -2586
rect 478794 -7654 479414 -2822
rect 483294 707718 483914 711590
rect 483294 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 483914 707718
rect 483294 707398 483914 707482
rect 483294 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 483914 707398
rect 483294 700954 483914 707162
rect 483294 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 483914 700954
rect 483294 700634 483914 700718
rect 483294 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 483914 700634
rect 483294 664954 483914 700398
rect 483294 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 483914 664954
rect 483294 664634 483914 664718
rect 483294 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 483914 664634
rect 483294 628954 483914 664398
rect 483294 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 483914 628954
rect 483294 628634 483914 628718
rect 483294 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 483914 628634
rect 483294 592954 483914 628398
rect 483294 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 483914 592954
rect 483294 592634 483914 592718
rect 483294 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 483914 592634
rect 483294 556954 483914 592398
rect 483294 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 483914 556954
rect 483294 556634 483914 556718
rect 483294 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 483914 556634
rect 483294 520954 483914 556398
rect 483294 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 483914 520954
rect 483294 520634 483914 520718
rect 483294 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 483914 520634
rect 483294 484954 483914 520398
rect 483294 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 483914 484954
rect 483294 484634 483914 484718
rect 483294 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 483914 484634
rect 483294 448954 483914 484398
rect 483294 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 483914 448954
rect 483294 448634 483914 448718
rect 483294 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 483914 448634
rect 483294 412954 483914 448398
rect 483294 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 483914 412954
rect 483294 412634 483914 412718
rect 483294 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 483914 412634
rect 483294 376954 483914 412398
rect 483294 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 483914 376954
rect 483294 376634 483914 376718
rect 483294 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 483914 376634
rect 483294 340954 483914 376398
rect 483294 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 483914 340954
rect 483294 340634 483914 340718
rect 483294 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 483914 340634
rect 483294 304954 483914 340398
rect 483294 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 483914 304954
rect 483294 304634 483914 304718
rect 483294 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 483914 304634
rect 483294 268954 483914 304398
rect 483294 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 483914 268954
rect 483294 268634 483914 268718
rect 483294 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 483914 268634
rect 483294 232954 483914 268398
rect 483294 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 483914 232954
rect 483294 232634 483914 232718
rect 483294 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 483914 232634
rect 483294 196954 483914 232398
rect 483294 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 483914 196954
rect 483294 196634 483914 196718
rect 483294 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 483914 196634
rect 483294 160954 483914 196398
rect 483294 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 483914 160954
rect 483294 160634 483914 160718
rect 483294 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 483914 160634
rect 483294 124954 483914 160398
rect 483294 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 483914 124954
rect 483294 124634 483914 124718
rect 483294 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 483914 124634
rect 483294 88954 483914 124398
rect 483294 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 483914 88954
rect 483294 88634 483914 88718
rect 483294 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 483914 88634
rect 483294 52954 483914 88398
rect 483294 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 483914 52954
rect 483294 52634 483914 52718
rect 483294 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 483914 52634
rect 483294 16954 483914 52398
rect 483294 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 483914 16954
rect 483294 16634 483914 16718
rect 483294 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 483914 16634
rect 483294 -3226 483914 16398
rect 483294 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 483914 -3226
rect 483294 -3546 483914 -3462
rect 483294 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 483914 -3546
rect 483294 -7654 483914 -3782
rect 487794 708678 488414 711590
rect 487794 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 488414 708678
rect 487794 708358 488414 708442
rect 487794 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 488414 708358
rect 487794 669454 488414 708122
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -4186 488414 20898
rect 487794 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 488414 -4186
rect 487794 -4506 488414 -4422
rect 487794 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 488414 -4506
rect 487794 -7654 488414 -4742
rect 492294 709638 492914 711590
rect 492294 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 492914 709638
rect 492294 709318 492914 709402
rect 492294 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 492914 709318
rect 492294 673954 492914 709082
rect 492294 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 492914 673954
rect 492294 673634 492914 673718
rect 492294 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 492914 673634
rect 492294 637954 492914 673398
rect 492294 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 492914 637954
rect 492294 637634 492914 637718
rect 492294 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 492914 637634
rect 492294 601954 492914 637398
rect 492294 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 492914 601954
rect 492294 601634 492914 601718
rect 492294 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 492914 601634
rect 492294 565954 492914 601398
rect 492294 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 492914 565954
rect 492294 565634 492914 565718
rect 492294 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 492914 565634
rect 492294 529954 492914 565398
rect 492294 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 492914 529954
rect 492294 529634 492914 529718
rect 492294 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 492914 529634
rect 492294 493954 492914 529398
rect 492294 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 492914 493954
rect 492294 493634 492914 493718
rect 492294 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 492914 493634
rect 492294 457954 492914 493398
rect 492294 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 492914 457954
rect 492294 457634 492914 457718
rect 492294 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 492914 457634
rect 492294 421954 492914 457398
rect 492294 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 492914 421954
rect 492294 421634 492914 421718
rect 492294 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 492914 421634
rect 492294 385954 492914 421398
rect 492294 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 492914 385954
rect 492294 385634 492914 385718
rect 492294 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 492914 385634
rect 492294 349954 492914 385398
rect 492294 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 492914 349954
rect 492294 349634 492914 349718
rect 492294 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 492914 349634
rect 492294 313954 492914 349398
rect 492294 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 492914 313954
rect 492294 313634 492914 313718
rect 492294 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 492914 313634
rect 492294 277954 492914 313398
rect 492294 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 492914 277954
rect 492294 277634 492914 277718
rect 492294 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 492914 277634
rect 492294 241954 492914 277398
rect 492294 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 492914 241954
rect 492294 241634 492914 241718
rect 492294 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 492914 241634
rect 492294 205954 492914 241398
rect 492294 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 492914 205954
rect 492294 205634 492914 205718
rect 492294 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 492914 205634
rect 492294 169954 492914 205398
rect 492294 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 492914 169954
rect 492294 169634 492914 169718
rect 492294 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 492914 169634
rect 492294 133954 492914 169398
rect 492294 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 492914 133954
rect 492294 133634 492914 133718
rect 492294 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 492914 133634
rect 492294 97954 492914 133398
rect 492294 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 492914 97954
rect 492294 97634 492914 97718
rect 492294 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 492914 97634
rect 492294 61954 492914 97398
rect 492294 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 492914 61954
rect 492294 61634 492914 61718
rect 492294 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 492914 61634
rect 492294 25954 492914 61398
rect 492294 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 492914 25954
rect 492294 25634 492914 25718
rect 492294 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 492914 25634
rect 492294 -5146 492914 25398
rect 492294 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 492914 -5146
rect 492294 -5466 492914 -5382
rect 492294 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 492914 -5466
rect 492294 -7654 492914 -5702
rect 496794 710598 497414 711590
rect 496794 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 497414 710598
rect 496794 710278 497414 710362
rect 496794 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 497414 710278
rect 496794 678454 497414 710042
rect 496794 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 497414 678454
rect 496794 678134 497414 678218
rect 496794 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 497414 678134
rect 496794 642454 497414 677898
rect 496794 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 497414 642454
rect 496794 642134 497414 642218
rect 496794 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 497414 642134
rect 496794 606454 497414 641898
rect 496794 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 497414 606454
rect 496794 606134 497414 606218
rect 496794 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 497414 606134
rect 496794 570454 497414 605898
rect 496794 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 497414 570454
rect 496794 570134 497414 570218
rect 496794 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 497414 570134
rect 496794 534454 497414 569898
rect 496794 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 497414 534454
rect 496794 534134 497414 534218
rect 496794 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 497414 534134
rect 496794 498454 497414 533898
rect 496794 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 497414 498454
rect 496794 498134 497414 498218
rect 496794 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 497414 498134
rect 496794 462454 497414 497898
rect 496794 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 497414 462454
rect 496794 462134 497414 462218
rect 496794 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 497414 462134
rect 496794 426454 497414 461898
rect 496794 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 497414 426454
rect 496794 426134 497414 426218
rect 496794 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 497414 426134
rect 496794 390454 497414 425898
rect 496794 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 497414 390454
rect 496794 390134 497414 390218
rect 496794 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 497414 390134
rect 496794 354454 497414 389898
rect 496794 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 497414 354454
rect 496794 354134 497414 354218
rect 496794 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 497414 354134
rect 496794 318454 497414 353898
rect 496794 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 497414 318454
rect 496794 318134 497414 318218
rect 496794 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 497414 318134
rect 496794 282454 497414 317898
rect 496794 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 497414 282454
rect 496794 282134 497414 282218
rect 496794 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 497414 282134
rect 496794 246454 497414 281898
rect 496794 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 497414 246454
rect 496794 246134 497414 246218
rect 496794 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 497414 246134
rect 496794 210454 497414 245898
rect 496794 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 497414 210454
rect 496794 210134 497414 210218
rect 496794 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 497414 210134
rect 496794 174454 497414 209898
rect 496794 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 497414 174454
rect 496794 174134 497414 174218
rect 496794 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 497414 174134
rect 496794 138454 497414 173898
rect 496794 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 497414 138454
rect 496794 138134 497414 138218
rect 496794 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 497414 138134
rect 496794 102454 497414 137898
rect 496794 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 497414 102454
rect 496794 102134 497414 102218
rect 496794 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 497414 102134
rect 496794 66454 497414 101898
rect 496794 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 497414 66454
rect 496794 66134 497414 66218
rect 496794 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 497414 66134
rect 496794 30454 497414 65898
rect 496794 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 497414 30454
rect 496794 30134 497414 30218
rect 496794 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 497414 30134
rect 496794 -6106 497414 29898
rect 496794 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 497414 -6106
rect 496794 -6426 497414 -6342
rect 496794 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 497414 -6426
rect 496794 -7654 497414 -6662
rect 501294 711558 501914 711590
rect 501294 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 501914 711558
rect 501294 711238 501914 711322
rect 501294 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 501914 711238
rect 501294 682954 501914 711002
rect 501294 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 501914 682954
rect 501294 682634 501914 682718
rect 501294 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 501914 682634
rect 501294 646954 501914 682398
rect 501294 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 501914 646954
rect 501294 646634 501914 646718
rect 501294 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 501914 646634
rect 501294 610954 501914 646398
rect 501294 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 501914 610954
rect 501294 610634 501914 610718
rect 501294 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 501914 610634
rect 501294 574954 501914 610398
rect 501294 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 501914 574954
rect 501294 574634 501914 574718
rect 501294 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 501914 574634
rect 501294 538954 501914 574398
rect 501294 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 501914 538954
rect 501294 538634 501914 538718
rect 501294 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 501914 538634
rect 501294 502954 501914 538398
rect 501294 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 501914 502954
rect 501294 502634 501914 502718
rect 501294 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 501914 502634
rect 501294 466954 501914 502398
rect 501294 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 501914 466954
rect 501294 466634 501914 466718
rect 501294 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 501914 466634
rect 501294 430954 501914 466398
rect 501294 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 501914 430954
rect 501294 430634 501914 430718
rect 501294 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 501914 430634
rect 501294 394954 501914 430398
rect 501294 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 501914 394954
rect 501294 394634 501914 394718
rect 501294 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 501914 394634
rect 501294 358954 501914 394398
rect 501294 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 501914 358954
rect 501294 358634 501914 358718
rect 501294 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 501914 358634
rect 501294 322954 501914 358398
rect 501294 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 501914 322954
rect 501294 322634 501914 322718
rect 501294 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 501914 322634
rect 501294 286954 501914 322398
rect 501294 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 501914 286954
rect 501294 286634 501914 286718
rect 501294 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 501914 286634
rect 501294 250954 501914 286398
rect 501294 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 501914 250954
rect 501294 250634 501914 250718
rect 501294 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 501914 250634
rect 501294 214954 501914 250398
rect 501294 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 501914 214954
rect 501294 214634 501914 214718
rect 501294 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 501914 214634
rect 501294 178954 501914 214398
rect 501294 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 501914 178954
rect 501294 178634 501914 178718
rect 501294 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 501914 178634
rect 501294 142954 501914 178398
rect 501294 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 501914 142954
rect 501294 142634 501914 142718
rect 501294 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 501914 142634
rect 501294 106954 501914 142398
rect 501294 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 501914 106954
rect 501294 106634 501914 106718
rect 501294 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 501914 106634
rect 501294 70954 501914 106398
rect 501294 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 501914 70954
rect 501294 70634 501914 70718
rect 501294 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 501914 70634
rect 501294 34954 501914 70398
rect 501294 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 501914 34954
rect 501294 34634 501914 34718
rect 501294 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 501914 34634
rect 501294 -7066 501914 34398
rect 501294 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 501914 -7066
rect 501294 -7386 501914 -7302
rect 501294 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 501914 -7386
rect 501294 -7654 501914 -7622
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 510294 705798 510914 711590
rect 510294 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 510914 705798
rect 510294 705478 510914 705562
rect 510294 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 510914 705478
rect 510294 691954 510914 705242
rect 510294 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 510914 691954
rect 510294 691634 510914 691718
rect 510294 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 510914 691634
rect 510294 655954 510914 691398
rect 510294 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 510914 655954
rect 510294 655634 510914 655718
rect 510294 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 510914 655634
rect 510294 619954 510914 655398
rect 510294 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 510914 619954
rect 510294 619634 510914 619718
rect 510294 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 510914 619634
rect 510294 583954 510914 619398
rect 510294 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 510914 583954
rect 510294 583634 510914 583718
rect 510294 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 510914 583634
rect 510294 547954 510914 583398
rect 510294 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 510914 547954
rect 510294 547634 510914 547718
rect 510294 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 510914 547634
rect 510294 511954 510914 547398
rect 510294 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 510914 511954
rect 510294 511634 510914 511718
rect 510294 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 510914 511634
rect 510294 475954 510914 511398
rect 510294 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 510914 475954
rect 510294 475634 510914 475718
rect 510294 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 510914 475634
rect 510294 439954 510914 475398
rect 510294 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 510914 439954
rect 510294 439634 510914 439718
rect 510294 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 510914 439634
rect 510294 403954 510914 439398
rect 510294 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 510914 403954
rect 510294 403634 510914 403718
rect 510294 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 510914 403634
rect 510294 367954 510914 403398
rect 510294 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 510914 367954
rect 510294 367634 510914 367718
rect 510294 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 510914 367634
rect 510294 331954 510914 367398
rect 510294 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 510914 331954
rect 510294 331634 510914 331718
rect 510294 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 510914 331634
rect 510294 295954 510914 331398
rect 510294 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 510914 295954
rect 510294 295634 510914 295718
rect 510294 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 510914 295634
rect 510294 259954 510914 295398
rect 510294 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 510914 259954
rect 510294 259634 510914 259718
rect 510294 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 510914 259634
rect 510294 223954 510914 259398
rect 510294 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 510914 223954
rect 510294 223634 510914 223718
rect 510294 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 510914 223634
rect 510294 187954 510914 223398
rect 510294 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 510914 187954
rect 510294 187634 510914 187718
rect 510294 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 510914 187634
rect 510294 151954 510914 187398
rect 510294 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 510914 151954
rect 510294 151634 510914 151718
rect 510294 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 510914 151634
rect 510294 115954 510914 151398
rect 510294 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 510914 115954
rect 510294 115634 510914 115718
rect 510294 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 510914 115634
rect 510294 79954 510914 115398
rect 510294 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 510914 79954
rect 510294 79634 510914 79718
rect 510294 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 510914 79634
rect 510294 43954 510914 79398
rect 510294 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 510914 43954
rect 510294 43634 510914 43718
rect 510294 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 510914 43634
rect 510294 7954 510914 43398
rect 510294 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 510914 7954
rect 510294 7634 510914 7718
rect 510294 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 510914 7634
rect 510294 -1306 510914 7398
rect 510294 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 510914 -1306
rect 510294 -1626 510914 -1542
rect 510294 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 510914 -1626
rect 510294 -7654 510914 -1862
rect 514794 706758 515414 711590
rect 514794 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 515414 706758
rect 514794 706438 515414 706522
rect 514794 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 515414 706438
rect 514794 696454 515414 706202
rect 514794 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 515414 696454
rect 514794 696134 515414 696218
rect 514794 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 515414 696134
rect 514794 660454 515414 695898
rect 514794 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 515414 660454
rect 514794 660134 515414 660218
rect 514794 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 515414 660134
rect 514794 624454 515414 659898
rect 514794 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 515414 624454
rect 514794 624134 515414 624218
rect 514794 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 515414 624134
rect 514794 588454 515414 623898
rect 514794 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 515414 588454
rect 514794 588134 515414 588218
rect 514794 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 515414 588134
rect 514794 552454 515414 587898
rect 514794 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 515414 552454
rect 514794 552134 515414 552218
rect 514794 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 515414 552134
rect 514794 516454 515414 551898
rect 514794 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 515414 516454
rect 514794 516134 515414 516218
rect 514794 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 515414 516134
rect 514794 480454 515414 515898
rect 514794 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 515414 480454
rect 514794 480134 515414 480218
rect 514794 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 515414 480134
rect 514794 444454 515414 479898
rect 514794 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 515414 444454
rect 514794 444134 515414 444218
rect 514794 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 515414 444134
rect 514794 408454 515414 443898
rect 514794 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 515414 408454
rect 514794 408134 515414 408218
rect 514794 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 515414 408134
rect 514794 372454 515414 407898
rect 514794 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 515414 372454
rect 514794 372134 515414 372218
rect 514794 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 515414 372134
rect 514794 336454 515414 371898
rect 514794 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 515414 336454
rect 514794 336134 515414 336218
rect 514794 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 515414 336134
rect 514794 300454 515414 335898
rect 514794 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 515414 300454
rect 514794 300134 515414 300218
rect 514794 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 515414 300134
rect 514794 264454 515414 299898
rect 514794 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 515414 264454
rect 514794 264134 515414 264218
rect 514794 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 515414 264134
rect 514794 228454 515414 263898
rect 514794 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 515414 228454
rect 514794 228134 515414 228218
rect 514794 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 515414 228134
rect 514794 192454 515414 227898
rect 514794 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 515414 192454
rect 514794 192134 515414 192218
rect 514794 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 515414 192134
rect 514794 156454 515414 191898
rect 514794 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 515414 156454
rect 514794 156134 515414 156218
rect 514794 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 515414 156134
rect 514794 120454 515414 155898
rect 514794 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 515414 120454
rect 514794 120134 515414 120218
rect 514794 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 515414 120134
rect 514794 84454 515414 119898
rect 514794 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 515414 84454
rect 514794 84134 515414 84218
rect 514794 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 515414 84134
rect 514794 48454 515414 83898
rect 514794 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 515414 48454
rect 514794 48134 515414 48218
rect 514794 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 515414 48134
rect 514794 12454 515414 47898
rect 514794 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 515414 12454
rect 514794 12134 515414 12218
rect 514794 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 515414 12134
rect 514794 -2266 515414 11898
rect 514794 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 515414 -2266
rect 514794 -2586 515414 -2502
rect 514794 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 515414 -2586
rect 514794 -7654 515414 -2822
rect 519294 707718 519914 711590
rect 519294 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 519914 707718
rect 519294 707398 519914 707482
rect 519294 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 519914 707398
rect 519294 700954 519914 707162
rect 519294 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 519914 700954
rect 519294 700634 519914 700718
rect 519294 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 519914 700634
rect 519294 664954 519914 700398
rect 519294 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 519914 664954
rect 519294 664634 519914 664718
rect 519294 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 519914 664634
rect 519294 628954 519914 664398
rect 519294 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 519914 628954
rect 519294 628634 519914 628718
rect 519294 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 519914 628634
rect 519294 592954 519914 628398
rect 519294 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 519914 592954
rect 519294 592634 519914 592718
rect 519294 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 519914 592634
rect 519294 556954 519914 592398
rect 519294 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 519914 556954
rect 519294 556634 519914 556718
rect 519294 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 519914 556634
rect 519294 520954 519914 556398
rect 519294 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 519914 520954
rect 519294 520634 519914 520718
rect 519294 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 519914 520634
rect 519294 484954 519914 520398
rect 519294 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 519914 484954
rect 519294 484634 519914 484718
rect 519294 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 519914 484634
rect 519294 448954 519914 484398
rect 519294 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 519914 448954
rect 519294 448634 519914 448718
rect 519294 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 519914 448634
rect 519294 412954 519914 448398
rect 519294 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 519914 412954
rect 519294 412634 519914 412718
rect 519294 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 519914 412634
rect 519294 376954 519914 412398
rect 519294 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 519914 376954
rect 519294 376634 519914 376718
rect 519294 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 519914 376634
rect 519294 340954 519914 376398
rect 519294 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 519914 340954
rect 519294 340634 519914 340718
rect 519294 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 519914 340634
rect 519294 304954 519914 340398
rect 519294 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 519914 304954
rect 519294 304634 519914 304718
rect 519294 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 519914 304634
rect 519294 268954 519914 304398
rect 519294 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 519914 268954
rect 519294 268634 519914 268718
rect 519294 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 519914 268634
rect 519294 232954 519914 268398
rect 519294 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 519914 232954
rect 519294 232634 519914 232718
rect 519294 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 519914 232634
rect 519294 196954 519914 232398
rect 519294 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 519914 196954
rect 519294 196634 519914 196718
rect 519294 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 519914 196634
rect 519294 160954 519914 196398
rect 519294 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 519914 160954
rect 519294 160634 519914 160718
rect 519294 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 519914 160634
rect 519294 124954 519914 160398
rect 519294 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 519914 124954
rect 519294 124634 519914 124718
rect 519294 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 519914 124634
rect 519294 88954 519914 124398
rect 519294 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 519914 88954
rect 519294 88634 519914 88718
rect 519294 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 519914 88634
rect 519294 52954 519914 88398
rect 519294 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 519914 52954
rect 519294 52634 519914 52718
rect 519294 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 519914 52634
rect 519294 16954 519914 52398
rect 519294 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 519914 16954
rect 519294 16634 519914 16718
rect 519294 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 519914 16634
rect 519294 -3226 519914 16398
rect 519294 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 519914 -3226
rect 519294 -3546 519914 -3462
rect 519294 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 519914 -3546
rect 519294 -7654 519914 -3782
rect 523794 708678 524414 711590
rect 523794 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 524414 708678
rect 523794 708358 524414 708442
rect 523794 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 524414 708358
rect 523794 669454 524414 708122
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -4186 524414 20898
rect 523794 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 524414 -4186
rect 523794 -4506 524414 -4422
rect 523794 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 524414 -4506
rect 523794 -7654 524414 -4742
rect 528294 709638 528914 711590
rect 528294 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 528914 709638
rect 528294 709318 528914 709402
rect 528294 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 528914 709318
rect 528294 673954 528914 709082
rect 528294 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 528914 673954
rect 528294 673634 528914 673718
rect 528294 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 528914 673634
rect 528294 637954 528914 673398
rect 528294 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 528914 637954
rect 528294 637634 528914 637718
rect 528294 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 528914 637634
rect 528294 601954 528914 637398
rect 528294 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 528914 601954
rect 528294 601634 528914 601718
rect 528294 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 528914 601634
rect 528294 565954 528914 601398
rect 528294 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 528914 565954
rect 528294 565634 528914 565718
rect 528294 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 528914 565634
rect 528294 529954 528914 565398
rect 528294 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 528914 529954
rect 528294 529634 528914 529718
rect 528294 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 528914 529634
rect 528294 493954 528914 529398
rect 528294 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 528914 493954
rect 528294 493634 528914 493718
rect 528294 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 528914 493634
rect 528294 457954 528914 493398
rect 528294 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 528914 457954
rect 528294 457634 528914 457718
rect 528294 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 528914 457634
rect 528294 421954 528914 457398
rect 528294 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 528914 421954
rect 528294 421634 528914 421718
rect 528294 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 528914 421634
rect 528294 385954 528914 421398
rect 528294 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 528914 385954
rect 528294 385634 528914 385718
rect 528294 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 528914 385634
rect 528294 349954 528914 385398
rect 528294 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 528914 349954
rect 528294 349634 528914 349718
rect 528294 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 528914 349634
rect 528294 313954 528914 349398
rect 528294 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 528914 313954
rect 528294 313634 528914 313718
rect 528294 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 528914 313634
rect 528294 277954 528914 313398
rect 528294 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 528914 277954
rect 528294 277634 528914 277718
rect 528294 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 528914 277634
rect 528294 241954 528914 277398
rect 528294 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 528914 241954
rect 528294 241634 528914 241718
rect 528294 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 528914 241634
rect 528294 205954 528914 241398
rect 528294 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 528914 205954
rect 528294 205634 528914 205718
rect 528294 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 528914 205634
rect 528294 169954 528914 205398
rect 528294 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 528914 169954
rect 528294 169634 528914 169718
rect 528294 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 528914 169634
rect 528294 133954 528914 169398
rect 528294 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 528914 133954
rect 528294 133634 528914 133718
rect 528294 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 528914 133634
rect 528294 97954 528914 133398
rect 528294 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 528914 97954
rect 528294 97634 528914 97718
rect 528294 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 528914 97634
rect 528294 61954 528914 97398
rect 528294 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 528914 61954
rect 528294 61634 528914 61718
rect 528294 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 528914 61634
rect 528294 25954 528914 61398
rect 528294 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 528914 25954
rect 528294 25634 528914 25718
rect 528294 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 528914 25634
rect 528294 -5146 528914 25398
rect 528294 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 528914 -5146
rect 528294 -5466 528914 -5382
rect 528294 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 528914 -5466
rect 528294 -7654 528914 -5702
rect 532794 710598 533414 711590
rect 532794 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 533414 710598
rect 532794 710278 533414 710362
rect 532794 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 533414 710278
rect 532794 678454 533414 710042
rect 532794 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 533414 678454
rect 532794 678134 533414 678218
rect 532794 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 533414 678134
rect 532794 642454 533414 677898
rect 532794 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 533414 642454
rect 532794 642134 533414 642218
rect 532794 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 533414 642134
rect 532794 606454 533414 641898
rect 532794 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 533414 606454
rect 532794 606134 533414 606218
rect 532794 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 533414 606134
rect 532794 570454 533414 605898
rect 532794 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 533414 570454
rect 532794 570134 533414 570218
rect 532794 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 533414 570134
rect 532794 534454 533414 569898
rect 532794 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 533414 534454
rect 532794 534134 533414 534218
rect 532794 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 533414 534134
rect 532794 498454 533414 533898
rect 532794 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 533414 498454
rect 532794 498134 533414 498218
rect 532794 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 533414 498134
rect 532794 462454 533414 497898
rect 532794 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 533414 462454
rect 532794 462134 533414 462218
rect 532794 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 533414 462134
rect 532794 426454 533414 461898
rect 532794 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 533414 426454
rect 532794 426134 533414 426218
rect 532794 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 533414 426134
rect 532794 390454 533414 425898
rect 532794 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 533414 390454
rect 532794 390134 533414 390218
rect 532794 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 533414 390134
rect 532794 354454 533414 389898
rect 532794 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 533414 354454
rect 532794 354134 533414 354218
rect 532794 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 533414 354134
rect 532794 318454 533414 353898
rect 532794 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 533414 318454
rect 532794 318134 533414 318218
rect 532794 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 533414 318134
rect 532794 282454 533414 317898
rect 532794 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 533414 282454
rect 532794 282134 533414 282218
rect 532794 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 533414 282134
rect 532794 246454 533414 281898
rect 532794 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 533414 246454
rect 532794 246134 533414 246218
rect 532794 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 533414 246134
rect 532794 210454 533414 245898
rect 532794 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 533414 210454
rect 532794 210134 533414 210218
rect 532794 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 533414 210134
rect 532794 174454 533414 209898
rect 532794 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 533414 174454
rect 532794 174134 533414 174218
rect 532794 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 533414 174134
rect 532794 138454 533414 173898
rect 532794 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 533414 138454
rect 532794 138134 533414 138218
rect 532794 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 533414 138134
rect 532794 102454 533414 137898
rect 532794 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 533414 102454
rect 532794 102134 533414 102218
rect 532794 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 533414 102134
rect 532794 66454 533414 101898
rect 532794 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 533414 66454
rect 532794 66134 533414 66218
rect 532794 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 533414 66134
rect 532794 30454 533414 65898
rect 532794 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 533414 30454
rect 532794 30134 533414 30218
rect 532794 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 533414 30134
rect 532794 -6106 533414 29898
rect 532794 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 533414 -6106
rect 532794 -6426 533414 -6342
rect 532794 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 533414 -6426
rect 532794 -7654 533414 -6662
rect 537294 711558 537914 711590
rect 537294 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 537914 711558
rect 537294 711238 537914 711322
rect 537294 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 537914 711238
rect 537294 682954 537914 711002
rect 537294 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 537914 682954
rect 537294 682634 537914 682718
rect 537294 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 537914 682634
rect 537294 646954 537914 682398
rect 537294 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 537914 646954
rect 537294 646634 537914 646718
rect 537294 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 537914 646634
rect 537294 610954 537914 646398
rect 537294 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 537914 610954
rect 537294 610634 537914 610718
rect 537294 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 537914 610634
rect 537294 574954 537914 610398
rect 537294 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 537914 574954
rect 537294 574634 537914 574718
rect 537294 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 537914 574634
rect 537294 538954 537914 574398
rect 537294 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 537914 538954
rect 537294 538634 537914 538718
rect 537294 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 537914 538634
rect 537294 502954 537914 538398
rect 537294 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 537914 502954
rect 537294 502634 537914 502718
rect 537294 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 537914 502634
rect 537294 466954 537914 502398
rect 537294 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 537914 466954
rect 537294 466634 537914 466718
rect 537294 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 537914 466634
rect 537294 430954 537914 466398
rect 537294 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 537914 430954
rect 537294 430634 537914 430718
rect 537294 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 537914 430634
rect 537294 394954 537914 430398
rect 537294 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 537914 394954
rect 537294 394634 537914 394718
rect 537294 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 537914 394634
rect 537294 358954 537914 394398
rect 537294 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 537914 358954
rect 537294 358634 537914 358718
rect 537294 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 537914 358634
rect 537294 322954 537914 358398
rect 537294 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 537914 322954
rect 537294 322634 537914 322718
rect 537294 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 537914 322634
rect 537294 286954 537914 322398
rect 537294 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 537914 286954
rect 537294 286634 537914 286718
rect 537294 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 537914 286634
rect 537294 250954 537914 286398
rect 537294 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 537914 250954
rect 537294 250634 537914 250718
rect 537294 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 537914 250634
rect 537294 214954 537914 250398
rect 537294 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 537914 214954
rect 537294 214634 537914 214718
rect 537294 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 537914 214634
rect 537294 178954 537914 214398
rect 537294 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 537914 178954
rect 537294 178634 537914 178718
rect 537294 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 537914 178634
rect 537294 142954 537914 178398
rect 537294 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 537914 142954
rect 537294 142634 537914 142718
rect 537294 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 537914 142634
rect 537294 106954 537914 142398
rect 537294 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 537914 106954
rect 537294 106634 537914 106718
rect 537294 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 537914 106634
rect 537294 70954 537914 106398
rect 537294 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 537914 70954
rect 537294 70634 537914 70718
rect 537294 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 537914 70634
rect 537294 34954 537914 70398
rect 537294 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 537914 34954
rect 537294 34634 537914 34718
rect 537294 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 537914 34634
rect 537294 -7066 537914 34398
rect 537294 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 537914 -7066
rect 537294 -7386 537914 -7302
rect 537294 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 537914 -7386
rect 537294 -7654 537914 -7622
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 546294 705798 546914 711590
rect 546294 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 546914 705798
rect 546294 705478 546914 705562
rect 546294 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 546914 705478
rect 546294 691954 546914 705242
rect 546294 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 546914 691954
rect 546294 691634 546914 691718
rect 546294 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 546914 691634
rect 546294 655954 546914 691398
rect 546294 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 546914 655954
rect 546294 655634 546914 655718
rect 546294 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 546914 655634
rect 546294 619954 546914 655398
rect 546294 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 546914 619954
rect 546294 619634 546914 619718
rect 546294 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 546914 619634
rect 546294 583954 546914 619398
rect 546294 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 546914 583954
rect 546294 583634 546914 583718
rect 546294 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 546914 583634
rect 546294 547954 546914 583398
rect 546294 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 546914 547954
rect 546294 547634 546914 547718
rect 546294 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 546914 547634
rect 546294 511954 546914 547398
rect 546294 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 546914 511954
rect 546294 511634 546914 511718
rect 546294 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 546914 511634
rect 546294 475954 546914 511398
rect 546294 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 546914 475954
rect 546294 475634 546914 475718
rect 546294 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 546914 475634
rect 546294 439954 546914 475398
rect 546294 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 546914 439954
rect 546294 439634 546914 439718
rect 546294 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 546914 439634
rect 546294 403954 546914 439398
rect 546294 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 546914 403954
rect 546294 403634 546914 403718
rect 546294 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 546914 403634
rect 546294 367954 546914 403398
rect 546294 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 546914 367954
rect 546294 367634 546914 367718
rect 546294 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 546914 367634
rect 546294 331954 546914 367398
rect 546294 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 546914 331954
rect 546294 331634 546914 331718
rect 546294 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 546914 331634
rect 546294 295954 546914 331398
rect 546294 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 546914 295954
rect 546294 295634 546914 295718
rect 546294 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 546914 295634
rect 546294 259954 546914 295398
rect 546294 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 546914 259954
rect 546294 259634 546914 259718
rect 546294 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 546914 259634
rect 546294 223954 546914 259398
rect 546294 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 546914 223954
rect 546294 223634 546914 223718
rect 546294 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 546914 223634
rect 546294 187954 546914 223398
rect 546294 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 546914 187954
rect 546294 187634 546914 187718
rect 546294 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 546914 187634
rect 546294 151954 546914 187398
rect 546294 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 546914 151954
rect 546294 151634 546914 151718
rect 546294 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 546914 151634
rect 546294 115954 546914 151398
rect 546294 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 546914 115954
rect 546294 115634 546914 115718
rect 546294 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 546914 115634
rect 546294 79954 546914 115398
rect 546294 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 546914 79954
rect 546294 79634 546914 79718
rect 546294 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 546914 79634
rect 546294 43954 546914 79398
rect 546294 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 546914 43954
rect 546294 43634 546914 43718
rect 546294 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 546914 43634
rect 546294 7954 546914 43398
rect 546294 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 546914 7954
rect 546294 7634 546914 7718
rect 546294 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 546914 7634
rect 546294 -1306 546914 7398
rect 546294 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 546914 -1306
rect 546294 -1626 546914 -1542
rect 546294 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 546914 -1626
rect 546294 -7654 546914 -1862
rect 550794 706758 551414 711590
rect 550794 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 551414 706758
rect 550794 706438 551414 706522
rect 550794 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 551414 706438
rect 550794 696454 551414 706202
rect 550794 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 551414 696454
rect 550794 696134 551414 696218
rect 550794 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 551414 696134
rect 550794 660454 551414 695898
rect 550794 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 551414 660454
rect 550794 660134 551414 660218
rect 550794 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 551414 660134
rect 550794 624454 551414 659898
rect 550794 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 551414 624454
rect 550794 624134 551414 624218
rect 550794 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 551414 624134
rect 550794 588454 551414 623898
rect 550794 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 551414 588454
rect 550794 588134 551414 588218
rect 550794 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 551414 588134
rect 550794 552454 551414 587898
rect 550794 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 551414 552454
rect 550794 552134 551414 552218
rect 550794 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 551414 552134
rect 550794 516454 551414 551898
rect 550794 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 551414 516454
rect 550794 516134 551414 516218
rect 550794 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 551414 516134
rect 550794 480454 551414 515898
rect 550794 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 551414 480454
rect 550794 480134 551414 480218
rect 550794 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 551414 480134
rect 550794 444454 551414 479898
rect 550794 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 551414 444454
rect 550794 444134 551414 444218
rect 550794 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 551414 444134
rect 550794 408454 551414 443898
rect 550794 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 551414 408454
rect 550794 408134 551414 408218
rect 550794 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 551414 408134
rect 550794 372454 551414 407898
rect 550794 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 551414 372454
rect 550794 372134 551414 372218
rect 550794 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 551414 372134
rect 550794 336454 551414 371898
rect 550794 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 551414 336454
rect 550794 336134 551414 336218
rect 550794 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 551414 336134
rect 550794 300454 551414 335898
rect 550794 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 551414 300454
rect 550794 300134 551414 300218
rect 550794 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 551414 300134
rect 550794 264454 551414 299898
rect 550794 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 551414 264454
rect 550794 264134 551414 264218
rect 550794 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 551414 264134
rect 550794 228454 551414 263898
rect 550794 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 551414 228454
rect 550794 228134 551414 228218
rect 550794 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 551414 228134
rect 550794 192454 551414 227898
rect 550794 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 551414 192454
rect 550794 192134 551414 192218
rect 550794 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 551414 192134
rect 550794 156454 551414 191898
rect 550794 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 551414 156454
rect 550794 156134 551414 156218
rect 550794 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 551414 156134
rect 550794 120454 551414 155898
rect 550794 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 551414 120454
rect 550794 120134 551414 120218
rect 550794 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 551414 120134
rect 550794 84454 551414 119898
rect 550794 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 551414 84454
rect 550794 84134 551414 84218
rect 550794 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 551414 84134
rect 550794 48454 551414 83898
rect 550794 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 551414 48454
rect 550794 48134 551414 48218
rect 550794 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 551414 48134
rect 550794 12454 551414 47898
rect 550794 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 551414 12454
rect 550794 12134 551414 12218
rect 550794 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 551414 12134
rect 550794 -2266 551414 11898
rect 550794 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 551414 -2266
rect 550794 -2586 551414 -2502
rect 550794 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 551414 -2586
rect 550794 -7654 551414 -2822
rect 555294 707718 555914 711590
rect 555294 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 555914 707718
rect 555294 707398 555914 707482
rect 555294 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 555914 707398
rect 555294 700954 555914 707162
rect 555294 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 555914 700954
rect 555294 700634 555914 700718
rect 555294 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 555914 700634
rect 555294 664954 555914 700398
rect 555294 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 555914 664954
rect 555294 664634 555914 664718
rect 555294 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 555914 664634
rect 555294 628954 555914 664398
rect 555294 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 555914 628954
rect 555294 628634 555914 628718
rect 555294 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 555914 628634
rect 555294 592954 555914 628398
rect 555294 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 555914 592954
rect 555294 592634 555914 592718
rect 555294 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 555914 592634
rect 555294 556954 555914 592398
rect 555294 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 555914 556954
rect 555294 556634 555914 556718
rect 555294 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 555914 556634
rect 555294 520954 555914 556398
rect 555294 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 555914 520954
rect 555294 520634 555914 520718
rect 555294 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 555914 520634
rect 555294 484954 555914 520398
rect 555294 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 555914 484954
rect 555294 484634 555914 484718
rect 555294 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 555914 484634
rect 555294 448954 555914 484398
rect 555294 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 555914 448954
rect 555294 448634 555914 448718
rect 555294 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 555914 448634
rect 555294 412954 555914 448398
rect 555294 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 555914 412954
rect 555294 412634 555914 412718
rect 555294 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 555914 412634
rect 555294 376954 555914 412398
rect 555294 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 555914 376954
rect 555294 376634 555914 376718
rect 555294 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 555914 376634
rect 555294 340954 555914 376398
rect 555294 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 555914 340954
rect 555294 340634 555914 340718
rect 555294 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 555914 340634
rect 555294 304954 555914 340398
rect 555294 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 555914 304954
rect 555294 304634 555914 304718
rect 555294 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 555914 304634
rect 555294 268954 555914 304398
rect 555294 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 555914 268954
rect 555294 268634 555914 268718
rect 555294 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 555914 268634
rect 555294 232954 555914 268398
rect 555294 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 555914 232954
rect 555294 232634 555914 232718
rect 555294 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 555914 232634
rect 555294 196954 555914 232398
rect 555294 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 555914 196954
rect 555294 196634 555914 196718
rect 555294 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 555914 196634
rect 555294 160954 555914 196398
rect 555294 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 555914 160954
rect 555294 160634 555914 160718
rect 555294 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 555914 160634
rect 555294 124954 555914 160398
rect 555294 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 555914 124954
rect 555294 124634 555914 124718
rect 555294 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 555914 124634
rect 555294 88954 555914 124398
rect 555294 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 555914 88954
rect 555294 88634 555914 88718
rect 555294 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 555914 88634
rect 555294 52954 555914 88398
rect 555294 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 555914 52954
rect 555294 52634 555914 52718
rect 555294 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 555914 52634
rect 555294 16954 555914 52398
rect 555294 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 555914 16954
rect 555294 16634 555914 16718
rect 555294 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 555914 16634
rect 555294 -3226 555914 16398
rect 555294 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 555914 -3226
rect 555294 -3546 555914 -3462
rect 555294 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 555914 -3546
rect 555294 -7654 555914 -3782
rect 559794 708678 560414 711590
rect 559794 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 560414 708678
rect 559794 708358 560414 708442
rect 559794 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 560414 708358
rect 559794 669454 560414 708122
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -4186 560414 20898
rect 559794 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 560414 -4186
rect 559794 -4506 560414 -4422
rect 559794 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 560414 -4506
rect 559794 -7654 560414 -4742
rect 564294 709638 564914 711590
rect 564294 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 564914 709638
rect 564294 709318 564914 709402
rect 564294 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 564914 709318
rect 564294 673954 564914 709082
rect 564294 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 564914 673954
rect 564294 673634 564914 673718
rect 564294 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 564914 673634
rect 564294 637954 564914 673398
rect 564294 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 564914 637954
rect 564294 637634 564914 637718
rect 564294 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 564914 637634
rect 564294 601954 564914 637398
rect 564294 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 564914 601954
rect 564294 601634 564914 601718
rect 564294 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 564914 601634
rect 564294 565954 564914 601398
rect 564294 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 564914 565954
rect 564294 565634 564914 565718
rect 564294 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 564914 565634
rect 564294 529954 564914 565398
rect 564294 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 564914 529954
rect 564294 529634 564914 529718
rect 564294 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 564914 529634
rect 564294 493954 564914 529398
rect 564294 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 564914 493954
rect 564294 493634 564914 493718
rect 564294 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 564914 493634
rect 564294 457954 564914 493398
rect 564294 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 564914 457954
rect 564294 457634 564914 457718
rect 564294 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 564914 457634
rect 564294 421954 564914 457398
rect 564294 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 564914 421954
rect 564294 421634 564914 421718
rect 564294 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 564914 421634
rect 564294 385954 564914 421398
rect 564294 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 564914 385954
rect 564294 385634 564914 385718
rect 564294 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 564914 385634
rect 564294 349954 564914 385398
rect 564294 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 564914 349954
rect 564294 349634 564914 349718
rect 564294 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 564914 349634
rect 564294 313954 564914 349398
rect 564294 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 564914 313954
rect 564294 313634 564914 313718
rect 564294 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 564914 313634
rect 564294 277954 564914 313398
rect 564294 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 564914 277954
rect 564294 277634 564914 277718
rect 564294 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 564914 277634
rect 564294 241954 564914 277398
rect 564294 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 564914 241954
rect 564294 241634 564914 241718
rect 564294 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 564914 241634
rect 564294 205954 564914 241398
rect 564294 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 564914 205954
rect 564294 205634 564914 205718
rect 564294 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 564914 205634
rect 564294 169954 564914 205398
rect 564294 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 564914 169954
rect 564294 169634 564914 169718
rect 564294 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 564914 169634
rect 564294 133954 564914 169398
rect 564294 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 564914 133954
rect 564294 133634 564914 133718
rect 564294 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 564914 133634
rect 564294 97954 564914 133398
rect 564294 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 564914 97954
rect 564294 97634 564914 97718
rect 564294 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 564914 97634
rect 564294 61954 564914 97398
rect 564294 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 564914 61954
rect 564294 61634 564914 61718
rect 564294 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 564914 61634
rect 564294 25954 564914 61398
rect 564294 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 564914 25954
rect 564294 25634 564914 25718
rect 564294 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 564914 25634
rect 564294 -5146 564914 25398
rect 564294 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 564914 -5146
rect 564294 -5466 564914 -5382
rect 564294 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 564914 -5466
rect 564294 -7654 564914 -5702
rect 568794 710598 569414 711590
rect 568794 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 569414 710598
rect 568794 710278 569414 710362
rect 568794 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 569414 710278
rect 568794 678454 569414 710042
rect 568794 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 569414 678454
rect 568794 678134 569414 678218
rect 568794 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 569414 678134
rect 568794 642454 569414 677898
rect 568794 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 569414 642454
rect 568794 642134 569414 642218
rect 568794 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 569414 642134
rect 568794 606454 569414 641898
rect 568794 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 569414 606454
rect 568794 606134 569414 606218
rect 568794 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 569414 606134
rect 568794 570454 569414 605898
rect 568794 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 569414 570454
rect 568794 570134 569414 570218
rect 568794 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 569414 570134
rect 568794 534454 569414 569898
rect 568794 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 569414 534454
rect 568794 534134 569414 534218
rect 568794 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 569414 534134
rect 568794 498454 569414 533898
rect 568794 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 569414 498454
rect 568794 498134 569414 498218
rect 568794 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 569414 498134
rect 568794 462454 569414 497898
rect 568794 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 569414 462454
rect 568794 462134 569414 462218
rect 568794 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 569414 462134
rect 568794 426454 569414 461898
rect 568794 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 569414 426454
rect 568794 426134 569414 426218
rect 568794 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 569414 426134
rect 568794 390454 569414 425898
rect 568794 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 569414 390454
rect 568794 390134 569414 390218
rect 568794 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 569414 390134
rect 568794 354454 569414 389898
rect 568794 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 569414 354454
rect 568794 354134 569414 354218
rect 568794 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 569414 354134
rect 568794 318454 569414 353898
rect 568794 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 569414 318454
rect 568794 318134 569414 318218
rect 568794 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 569414 318134
rect 568794 282454 569414 317898
rect 568794 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 569414 282454
rect 568794 282134 569414 282218
rect 568794 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 569414 282134
rect 568794 246454 569414 281898
rect 568794 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 569414 246454
rect 568794 246134 569414 246218
rect 568794 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 569414 246134
rect 568794 210454 569414 245898
rect 568794 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 569414 210454
rect 568794 210134 569414 210218
rect 568794 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 569414 210134
rect 568794 174454 569414 209898
rect 568794 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 569414 174454
rect 568794 174134 569414 174218
rect 568794 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 569414 174134
rect 568794 138454 569414 173898
rect 568794 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 569414 138454
rect 568794 138134 569414 138218
rect 568794 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 569414 138134
rect 568794 102454 569414 137898
rect 568794 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 569414 102454
rect 568794 102134 569414 102218
rect 568794 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 569414 102134
rect 568794 66454 569414 101898
rect 568794 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 569414 66454
rect 568794 66134 569414 66218
rect 568794 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 569414 66134
rect 568794 30454 569414 65898
rect 568794 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 569414 30454
rect 568794 30134 569414 30218
rect 568794 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 569414 30134
rect 568794 -6106 569414 29898
rect 568794 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 569414 -6106
rect 568794 -6426 569414 -6342
rect 568794 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 569414 -6426
rect 568794 -7654 569414 -6662
rect 573294 711558 573914 711590
rect 573294 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 573914 711558
rect 573294 711238 573914 711322
rect 573294 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 573914 711238
rect 573294 682954 573914 711002
rect 573294 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 573914 682954
rect 573294 682634 573914 682718
rect 573294 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 573914 682634
rect 573294 646954 573914 682398
rect 573294 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 573914 646954
rect 573294 646634 573914 646718
rect 573294 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 573914 646634
rect 573294 610954 573914 646398
rect 573294 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 573914 610954
rect 573294 610634 573914 610718
rect 573294 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 573914 610634
rect 573294 574954 573914 610398
rect 573294 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 573914 574954
rect 573294 574634 573914 574718
rect 573294 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 573914 574634
rect 573294 538954 573914 574398
rect 573294 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 573914 538954
rect 573294 538634 573914 538718
rect 573294 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 573914 538634
rect 573294 502954 573914 538398
rect 573294 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 573914 502954
rect 573294 502634 573914 502718
rect 573294 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 573914 502634
rect 573294 466954 573914 502398
rect 573294 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 573914 466954
rect 573294 466634 573914 466718
rect 573294 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 573914 466634
rect 573294 430954 573914 466398
rect 573294 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 573914 430954
rect 573294 430634 573914 430718
rect 573294 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 573914 430634
rect 573294 394954 573914 430398
rect 573294 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 573914 394954
rect 573294 394634 573914 394718
rect 573294 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 573914 394634
rect 573294 358954 573914 394398
rect 573294 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 573914 358954
rect 573294 358634 573914 358718
rect 573294 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 573914 358634
rect 573294 322954 573914 358398
rect 573294 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 573914 322954
rect 573294 322634 573914 322718
rect 573294 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 573914 322634
rect 573294 286954 573914 322398
rect 573294 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 573914 286954
rect 573294 286634 573914 286718
rect 573294 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 573914 286634
rect 573294 250954 573914 286398
rect 573294 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 573914 250954
rect 573294 250634 573914 250718
rect 573294 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 573914 250634
rect 573294 214954 573914 250398
rect 573294 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 573914 214954
rect 573294 214634 573914 214718
rect 573294 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 573914 214634
rect 573294 178954 573914 214398
rect 573294 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 573914 178954
rect 573294 178634 573914 178718
rect 573294 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 573914 178634
rect 573294 142954 573914 178398
rect 573294 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 573914 142954
rect 573294 142634 573914 142718
rect 573294 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 573914 142634
rect 573294 106954 573914 142398
rect 573294 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 573914 106954
rect 573294 106634 573914 106718
rect 573294 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 573914 106634
rect 573294 70954 573914 106398
rect 573294 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 573914 70954
rect 573294 70634 573914 70718
rect 573294 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 573914 70634
rect 573294 34954 573914 70398
rect 573294 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 573914 34954
rect 573294 34634 573914 34718
rect 573294 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 573914 34634
rect 573294 -7066 573914 34398
rect 573294 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 573914 -7066
rect 573294 -7386 573914 -7302
rect 573294 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 573914 -7386
rect 573294 -7654 573914 -7622
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 582294 705798 582914 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 582294 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 582914 705798
rect 582294 705478 582914 705562
rect 582294 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 582914 705478
rect 582294 691954 582914 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 582294 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 582914 691954
rect 582294 691634 582914 691718
rect 582294 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 582914 691634
rect 582294 655954 582914 691398
rect 582294 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 582914 655954
rect 582294 655634 582914 655718
rect 582294 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 582914 655634
rect 582294 619954 582914 655398
rect 582294 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 582914 619954
rect 582294 619634 582914 619718
rect 582294 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 582914 619634
rect 582294 583954 582914 619398
rect 582294 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 582914 583954
rect 582294 583634 582914 583718
rect 582294 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 582914 583634
rect 582294 547954 582914 583398
rect 582294 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 582914 547954
rect 582294 547634 582914 547718
rect 582294 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 582914 547634
rect 582294 511954 582914 547398
rect 582294 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 582914 511954
rect 582294 511634 582914 511718
rect 582294 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 582914 511634
rect 582294 475954 582914 511398
rect 582294 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 582914 475954
rect 582294 475634 582914 475718
rect 582294 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 582914 475634
rect 582294 439954 582914 475398
rect 582294 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 582914 439954
rect 582294 439634 582914 439718
rect 582294 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 582914 439634
rect 582294 403954 582914 439398
rect 582294 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 582914 403954
rect 582294 403634 582914 403718
rect 582294 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 582914 403634
rect 582294 367954 582914 403398
rect 582294 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 582914 367954
rect 582294 367634 582914 367718
rect 582294 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 582914 367634
rect 582294 331954 582914 367398
rect 582294 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 582914 331954
rect 582294 331634 582914 331718
rect 582294 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 582914 331634
rect 582294 295954 582914 331398
rect 582294 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 582914 295954
rect 582294 295634 582914 295718
rect 582294 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 582914 295634
rect 582294 259954 582914 295398
rect 582294 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 582914 259954
rect 582294 259634 582914 259718
rect 582294 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 582914 259634
rect 582294 223954 582914 259398
rect 582294 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 582914 223954
rect 582294 223634 582914 223718
rect 582294 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 582914 223634
rect 582294 187954 582914 223398
rect 582294 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 582914 187954
rect 582294 187634 582914 187718
rect 582294 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 582914 187634
rect 582294 151954 582914 187398
rect 582294 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 582914 151954
rect 582294 151634 582914 151718
rect 582294 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 582914 151634
rect 582294 115954 582914 151398
rect 582294 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 582914 115954
rect 582294 115634 582914 115718
rect 582294 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 582914 115634
rect 582294 79954 582914 115398
rect 582294 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 582914 79954
rect 582294 79634 582914 79718
rect 582294 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 582914 79634
rect 582294 43954 582914 79398
rect 582294 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 582914 43954
rect 582294 43634 582914 43718
rect 582294 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 582914 43634
rect 582294 7954 582914 43398
rect 582294 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 582914 7954
rect 582294 7634 582914 7718
rect 582294 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 582914 7634
rect 582294 -1306 582914 7398
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691954 586890 705242
rect 586270 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 586890 691954
rect 586270 691634 586890 691718
rect 586270 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 586890 691634
rect 586270 655954 586890 691398
rect 586270 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 586890 655954
rect 586270 655634 586890 655718
rect 586270 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 586890 655634
rect 586270 619954 586890 655398
rect 586270 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 586890 619954
rect 586270 619634 586890 619718
rect 586270 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 586890 619634
rect 586270 583954 586890 619398
rect 586270 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 586890 583954
rect 586270 583634 586890 583718
rect 586270 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 586890 583634
rect 586270 547954 586890 583398
rect 586270 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 586890 547954
rect 586270 547634 586890 547718
rect 586270 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 586890 547634
rect 586270 511954 586890 547398
rect 586270 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 586890 511954
rect 586270 511634 586890 511718
rect 586270 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 586890 511634
rect 586270 475954 586890 511398
rect 586270 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 586890 475954
rect 586270 475634 586890 475718
rect 586270 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 586890 475634
rect 586270 439954 586890 475398
rect 586270 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 586890 439954
rect 586270 439634 586890 439718
rect 586270 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 586890 439634
rect 586270 403954 586890 439398
rect 586270 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 586890 403954
rect 586270 403634 586890 403718
rect 586270 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 586890 403634
rect 586270 367954 586890 403398
rect 586270 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 586890 367954
rect 586270 367634 586890 367718
rect 586270 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 586890 367634
rect 586270 331954 586890 367398
rect 586270 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 586890 331954
rect 586270 331634 586890 331718
rect 586270 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 586890 331634
rect 586270 295954 586890 331398
rect 586270 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 586890 295954
rect 586270 295634 586890 295718
rect 586270 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 586890 295634
rect 586270 259954 586890 295398
rect 586270 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 586890 259954
rect 586270 259634 586890 259718
rect 586270 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 586890 259634
rect 586270 223954 586890 259398
rect 586270 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 586890 223954
rect 586270 223634 586890 223718
rect 586270 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 586890 223634
rect 586270 187954 586890 223398
rect 586270 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 586890 187954
rect 586270 187634 586890 187718
rect 586270 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 586890 187634
rect 586270 151954 586890 187398
rect 586270 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 586890 151954
rect 586270 151634 586890 151718
rect 586270 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 586890 151634
rect 586270 115954 586890 151398
rect 586270 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 586890 115954
rect 586270 115634 586890 115718
rect 586270 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 586890 115634
rect 586270 79954 586890 115398
rect 586270 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 586890 79954
rect 586270 79634 586890 79718
rect 586270 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 586890 79634
rect 586270 43954 586890 79398
rect 586270 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 586890 43954
rect 586270 43634 586890 43718
rect 586270 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 586890 43634
rect 586270 7954 586890 43398
rect 586270 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 586890 7954
rect 586270 7634 586890 7718
rect 586270 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 586890 7634
rect 582294 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 582914 -1306
rect 582294 -1626 582914 -1542
rect 582294 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 582914 -1626
rect 582294 -7654 582914 -1862
rect 586270 -1306 586890 7398
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 696454 587850 706202
rect 587230 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 587850 696454
rect 587230 696134 587850 696218
rect 587230 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 587850 696134
rect 587230 660454 587850 695898
rect 587230 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 587850 660454
rect 587230 660134 587850 660218
rect 587230 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 587850 660134
rect 587230 624454 587850 659898
rect 587230 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 587850 624454
rect 587230 624134 587850 624218
rect 587230 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 587850 624134
rect 587230 588454 587850 623898
rect 587230 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 587850 588454
rect 587230 588134 587850 588218
rect 587230 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 587850 588134
rect 587230 552454 587850 587898
rect 587230 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 587850 552454
rect 587230 552134 587850 552218
rect 587230 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 587850 552134
rect 587230 516454 587850 551898
rect 587230 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 587850 516454
rect 587230 516134 587850 516218
rect 587230 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 587850 516134
rect 587230 480454 587850 515898
rect 587230 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 587850 480454
rect 587230 480134 587850 480218
rect 587230 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 587850 480134
rect 587230 444454 587850 479898
rect 587230 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 587850 444454
rect 587230 444134 587850 444218
rect 587230 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 587850 444134
rect 587230 408454 587850 443898
rect 587230 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 587850 408454
rect 587230 408134 587850 408218
rect 587230 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 587850 408134
rect 587230 372454 587850 407898
rect 587230 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 587850 372454
rect 587230 372134 587850 372218
rect 587230 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 587850 372134
rect 587230 336454 587850 371898
rect 587230 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 587850 336454
rect 587230 336134 587850 336218
rect 587230 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 587850 336134
rect 587230 300454 587850 335898
rect 587230 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 587850 300454
rect 587230 300134 587850 300218
rect 587230 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 587850 300134
rect 587230 264454 587850 299898
rect 587230 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 587850 264454
rect 587230 264134 587850 264218
rect 587230 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 587850 264134
rect 587230 228454 587850 263898
rect 587230 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 587850 228454
rect 587230 228134 587850 228218
rect 587230 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 587850 228134
rect 587230 192454 587850 227898
rect 587230 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 587850 192454
rect 587230 192134 587850 192218
rect 587230 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 587850 192134
rect 587230 156454 587850 191898
rect 587230 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 587850 156454
rect 587230 156134 587850 156218
rect 587230 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 587850 156134
rect 587230 120454 587850 155898
rect 587230 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 587850 120454
rect 587230 120134 587850 120218
rect 587230 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 587850 120134
rect 587230 84454 587850 119898
rect 587230 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 587850 84454
rect 587230 84134 587850 84218
rect 587230 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 587850 84134
rect 587230 48454 587850 83898
rect 587230 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 587850 48454
rect 587230 48134 587850 48218
rect 587230 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 587850 48134
rect 587230 12454 587850 47898
rect 587230 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 587850 12454
rect 587230 12134 587850 12218
rect 587230 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 587850 12134
rect 587230 -2266 587850 11898
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 700954 588810 707162
rect 588190 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 588810 700954
rect 588190 700634 588810 700718
rect 588190 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 588810 700634
rect 588190 664954 588810 700398
rect 588190 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 588810 664954
rect 588190 664634 588810 664718
rect 588190 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 588810 664634
rect 588190 628954 588810 664398
rect 588190 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 588810 628954
rect 588190 628634 588810 628718
rect 588190 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 588810 628634
rect 588190 592954 588810 628398
rect 588190 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 588810 592954
rect 588190 592634 588810 592718
rect 588190 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 588810 592634
rect 588190 556954 588810 592398
rect 588190 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 588810 556954
rect 588190 556634 588810 556718
rect 588190 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 588810 556634
rect 588190 520954 588810 556398
rect 588190 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 588810 520954
rect 588190 520634 588810 520718
rect 588190 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 588810 520634
rect 588190 484954 588810 520398
rect 588190 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 588810 484954
rect 588190 484634 588810 484718
rect 588190 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 588810 484634
rect 588190 448954 588810 484398
rect 588190 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 588810 448954
rect 588190 448634 588810 448718
rect 588190 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 588810 448634
rect 588190 412954 588810 448398
rect 588190 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 588810 412954
rect 588190 412634 588810 412718
rect 588190 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 588810 412634
rect 588190 376954 588810 412398
rect 588190 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 588810 376954
rect 588190 376634 588810 376718
rect 588190 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 588810 376634
rect 588190 340954 588810 376398
rect 588190 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 588810 340954
rect 588190 340634 588810 340718
rect 588190 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 588810 340634
rect 588190 304954 588810 340398
rect 588190 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 588810 304954
rect 588190 304634 588810 304718
rect 588190 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 588810 304634
rect 588190 268954 588810 304398
rect 588190 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 588810 268954
rect 588190 268634 588810 268718
rect 588190 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 588810 268634
rect 588190 232954 588810 268398
rect 588190 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 588810 232954
rect 588190 232634 588810 232718
rect 588190 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 588810 232634
rect 588190 196954 588810 232398
rect 588190 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 588810 196954
rect 588190 196634 588810 196718
rect 588190 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 588810 196634
rect 588190 160954 588810 196398
rect 588190 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 588810 160954
rect 588190 160634 588810 160718
rect 588190 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 588810 160634
rect 588190 124954 588810 160398
rect 588190 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 588810 124954
rect 588190 124634 588810 124718
rect 588190 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 588810 124634
rect 588190 88954 588810 124398
rect 588190 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 588810 88954
rect 588190 88634 588810 88718
rect 588190 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 588810 88634
rect 588190 52954 588810 88398
rect 588190 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 588810 52954
rect 588190 52634 588810 52718
rect 588190 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 588810 52634
rect 588190 16954 588810 52398
rect 588190 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 588810 16954
rect 588190 16634 588810 16718
rect 588190 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 588810 16634
rect 588190 -3226 588810 16398
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 669454 589770 708122
rect 589150 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 589770 669454
rect 589150 669134 589770 669218
rect 589150 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 589770 669134
rect 589150 633454 589770 668898
rect 589150 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 589770 633454
rect 589150 633134 589770 633218
rect 589150 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 589770 633134
rect 589150 597454 589770 632898
rect 589150 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 589770 597454
rect 589150 597134 589770 597218
rect 589150 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 589770 597134
rect 589150 561454 589770 596898
rect 589150 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 589770 561454
rect 589150 561134 589770 561218
rect 589150 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 589770 561134
rect 589150 525454 589770 560898
rect 589150 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 589770 525454
rect 589150 525134 589770 525218
rect 589150 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 589770 525134
rect 589150 489454 589770 524898
rect 589150 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 589770 489454
rect 589150 489134 589770 489218
rect 589150 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 589770 489134
rect 589150 453454 589770 488898
rect 589150 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 589770 453454
rect 589150 453134 589770 453218
rect 589150 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 589770 453134
rect 589150 417454 589770 452898
rect 589150 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 589770 417454
rect 589150 417134 589770 417218
rect 589150 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 589770 417134
rect 589150 381454 589770 416898
rect 589150 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 589770 381454
rect 589150 381134 589770 381218
rect 589150 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 589770 381134
rect 589150 345454 589770 380898
rect 589150 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 589770 345454
rect 589150 345134 589770 345218
rect 589150 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 589770 345134
rect 589150 309454 589770 344898
rect 589150 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 589770 309454
rect 589150 309134 589770 309218
rect 589150 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 589770 309134
rect 589150 273454 589770 308898
rect 589150 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 589770 273454
rect 589150 273134 589770 273218
rect 589150 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 589770 273134
rect 589150 237454 589770 272898
rect 589150 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 589770 237454
rect 589150 237134 589770 237218
rect 589150 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 589770 237134
rect 589150 201454 589770 236898
rect 589150 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 589770 201454
rect 589150 201134 589770 201218
rect 589150 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 589770 201134
rect 589150 165454 589770 200898
rect 589150 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 589770 165454
rect 589150 165134 589770 165218
rect 589150 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 589770 165134
rect 589150 129454 589770 164898
rect 589150 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 589770 129454
rect 589150 129134 589770 129218
rect 589150 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 589770 129134
rect 589150 93454 589770 128898
rect 589150 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 589770 93454
rect 589150 93134 589770 93218
rect 589150 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 589770 93134
rect 589150 57454 589770 92898
rect 589150 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 589770 57454
rect 589150 57134 589770 57218
rect 589150 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 589770 57134
rect 589150 21454 589770 56898
rect 589150 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 589770 21454
rect 589150 21134 589770 21218
rect 589150 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 589770 21134
rect 589150 -4186 589770 20898
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 673954 590730 709082
rect 590110 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 590730 673954
rect 590110 673634 590730 673718
rect 590110 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 590730 673634
rect 590110 637954 590730 673398
rect 590110 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 590730 637954
rect 590110 637634 590730 637718
rect 590110 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 590730 637634
rect 590110 601954 590730 637398
rect 590110 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 590730 601954
rect 590110 601634 590730 601718
rect 590110 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 590730 601634
rect 590110 565954 590730 601398
rect 590110 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 590730 565954
rect 590110 565634 590730 565718
rect 590110 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 590730 565634
rect 590110 529954 590730 565398
rect 590110 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 590730 529954
rect 590110 529634 590730 529718
rect 590110 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 590730 529634
rect 590110 493954 590730 529398
rect 590110 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 590730 493954
rect 590110 493634 590730 493718
rect 590110 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 590730 493634
rect 590110 457954 590730 493398
rect 590110 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 590730 457954
rect 590110 457634 590730 457718
rect 590110 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 590730 457634
rect 590110 421954 590730 457398
rect 590110 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 590730 421954
rect 590110 421634 590730 421718
rect 590110 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 590730 421634
rect 590110 385954 590730 421398
rect 590110 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 590730 385954
rect 590110 385634 590730 385718
rect 590110 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 590730 385634
rect 590110 349954 590730 385398
rect 590110 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 590730 349954
rect 590110 349634 590730 349718
rect 590110 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 590730 349634
rect 590110 313954 590730 349398
rect 590110 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 590730 313954
rect 590110 313634 590730 313718
rect 590110 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 590730 313634
rect 590110 277954 590730 313398
rect 590110 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 590730 277954
rect 590110 277634 590730 277718
rect 590110 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 590730 277634
rect 590110 241954 590730 277398
rect 590110 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 590730 241954
rect 590110 241634 590730 241718
rect 590110 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 590730 241634
rect 590110 205954 590730 241398
rect 590110 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 590730 205954
rect 590110 205634 590730 205718
rect 590110 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 590730 205634
rect 590110 169954 590730 205398
rect 590110 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 590730 169954
rect 590110 169634 590730 169718
rect 590110 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 590730 169634
rect 590110 133954 590730 169398
rect 590110 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 590730 133954
rect 590110 133634 590730 133718
rect 590110 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 590730 133634
rect 590110 97954 590730 133398
rect 590110 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 590730 97954
rect 590110 97634 590730 97718
rect 590110 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 590730 97634
rect 590110 61954 590730 97398
rect 590110 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 590730 61954
rect 590110 61634 590730 61718
rect 590110 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 590730 61634
rect 590110 25954 590730 61398
rect 590110 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 590730 25954
rect 590110 25634 590730 25718
rect 590110 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 590730 25634
rect 590110 -5146 590730 25398
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 678454 591690 710042
rect 591070 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 591690 678454
rect 591070 678134 591690 678218
rect 591070 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 591690 678134
rect 591070 642454 591690 677898
rect 591070 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 591690 642454
rect 591070 642134 591690 642218
rect 591070 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 591690 642134
rect 591070 606454 591690 641898
rect 591070 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 591690 606454
rect 591070 606134 591690 606218
rect 591070 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 591690 606134
rect 591070 570454 591690 605898
rect 591070 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 591690 570454
rect 591070 570134 591690 570218
rect 591070 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 591690 570134
rect 591070 534454 591690 569898
rect 591070 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 591690 534454
rect 591070 534134 591690 534218
rect 591070 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 591690 534134
rect 591070 498454 591690 533898
rect 591070 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 591690 498454
rect 591070 498134 591690 498218
rect 591070 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 591690 498134
rect 591070 462454 591690 497898
rect 591070 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 591690 462454
rect 591070 462134 591690 462218
rect 591070 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 591690 462134
rect 591070 426454 591690 461898
rect 591070 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 591690 426454
rect 591070 426134 591690 426218
rect 591070 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 591690 426134
rect 591070 390454 591690 425898
rect 591070 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 591690 390454
rect 591070 390134 591690 390218
rect 591070 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 591690 390134
rect 591070 354454 591690 389898
rect 591070 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 591690 354454
rect 591070 354134 591690 354218
rect 591070 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 591690 354134
rect 591070 318454 591690 353898
rect 591070 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 591690 318454
rect 591070 318134 591690 318218
rect 591070 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 591690 318134
rect 591070 282454 591690 317898
rect 591070 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 591690 282454
rect 591070 282134 591690 282218
rect 591070 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 591690 282134
rect 591070 246454 591690 281898
rect 591070 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 591690 246454
rect 591070 246134 591690 246218
rect 591070 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 591690 246134
rect 591070 210454 591690 245898
rect 591070 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 591690 210454
rect 591070 210134 591690 210218
rect 591070 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 591690 210134
rect 591070 174454 591690 209898
rect 591070 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 591690 174454
rect 591070 174134 591690 174218
rect 591070 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 591690 174134
rect 591070 138454 591690 173898
rect 591070 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 591690 138454
rect 591070 138134 591690 138218
rect 591070 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 591690 138134
rect 591070 102454 591690 137898
rect 591070 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 591690 102454
rect 591070 102134 591690 102218
rect 591070 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 591690 102134
rect 591070 66454 591690 101898
rect 591070 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 591690 66454
rect 591070 66134 591690 66218
rect 591070 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 591690 66134
rect 591070 30454 591690 65898
rect 591070 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 591690 30454
rect 591070 30134 591690 30218
rect 591070 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 591690 30134
rect 591070 -6106 591690 29898
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 682954 592650 711002
rect 592030 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect 592030 682634 592650 682718
rect 592030 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect 592030 646954 592650 682398
rect 592030 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect 592030 646634 592650 646718
rect 592030 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect 592030 610954 592650 646398
rect 592030 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect 592030 610634 592650 610718
rect 592030 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect 592030 574954 592650 610398
rect 592030 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect 592030 574634 592650 574718
rect 592030 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect 592030 538954 592650 574398
rect 592030 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect 592030 538634 592650 538718
rect 592030 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect 592030 502954 592650 538398
rect 592030 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect 592030 502634 592650 502718
rect 592030 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect 592030 466954 592650 502398
rect 592030 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect 592030 466634 592650 466718
rect 592030 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect 592030 430954 592650 466398
rect 592030 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect 592030 430634 592650 430718
rect 592030 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect 592030 394954 592650 430398
rect 592030 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect 592030 394634 592650 394718
rect 592030 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect 592030 358954 592650 394398
rect 592030 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect 592030 358634 592650 358718
rect 592030 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect 592030 322954 592650 358398
rect 592030 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect 592030 322634 592650 322718
rect 592030 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect 592030 286954 592650 322398
rect 592030 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect 592030 286634 592650 286718
rect 592030 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect 592030 250954 592650 286398
rect 592030 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect 592030 250634 592650 250718
rect 592030 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect 592030 214954 592650 250398
rect 592030 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect 592030 214634 592650 214718
rect 592030 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect 592030 178954 592650 214398
rect 592030 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect 592030 178634 592650 178718
rect 592030 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect 592030 142954 592650 178398
rect 592030 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect 592030 142634 592650 142718
rect 592030 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect 592030 106954 592650 142398
rect 592030 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect 592030 106634 592650 106718
rect 592030 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect 592030 70954 592650 106398
rect 592030 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect 592030 70634 592650 70718
rect 592030 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect 592030 34954 592650 70398
rect 592030 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect 592030 34634 592650 34718
rect 592030 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect 592030 -7066 592650 34398
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 682718 -8458 682954
rect -8374 682718 -8138 682954
rect -8694 682398 -8458 682634
rect -8374 682398 -8138 682634
rect -8694 646718 -8458 646954
rect -8374 646718 -8138 646954
rect -8694 646398 -8458 646634
rect -8374 646398 -8138 646634
rect -8694 610718 -8458 610954
rect -8374 610718 -8138 610954
rect -8694 610398 -8458 610634
rect -8374 610398 -8138 610634
rect -8694 574718 -8458 574954
rect -8374 574718 -8138 574954
rect -8694 574398 -8458 574634
rect -8374 574398 -8138 574634
rect -8694 538718 -8458 538954
rect -8374 538718 -8138 538954
rect -8694 538398 -8458 538634
rect -8374 538398 -8138 538634
rect -8694 502718 -8458 502954
rect -8374 502718 -8138 502954
rect -8694 502398 -8458 502634
rect -8374 502398 -8138 502634
rect -8694 466718 -8458 466954
rect -8374 466718 -8138 466954
rect -8694 466398 -8458 466634
rect -8374 466398 -8138 466634
rect -8694 430718 -8458 430954
rect -8374 430718 -8138 430954
rect -8694 430398 -8458 430634
rect -8374 430398 -8138 430634
rect -8694 394718 -8458 394954
rect -8374 394718 -8138 394954
rect -8694 394398 -8458 394634
rect -8374 394398 -8138 394634
rect -8694 358718 -8458 358954
rect -8374 358718 -8138 358954
rect -8694 358398 -8458 358634
rect -8374 358398 -8138 358634
rect -8694 322718 -8458 322954
rect -8374 322718 -8138 322954
rect -8694 322398 -8458 322634
rect -8374 322398 -8138 322634
rect -8694 286718 -8458 286954
rect -8374 286718 -8138 286954
rect -8694 286398 -8458 286634
rect -8374 286398 -8138 286634
rect -8694 250718 -8458 250954
rect -8374 250718 -8138 250954
rect -8694 250398 -8458 250634
rect -8374 250398 -8138 250634
rect -8694 214718 -8458 214954
rect -8374 214718 -8138 214954
rect -8694 214398 -8458 214634
rect -8374 214398 -8138 214634
rect -8694 178718 -8458 178954
rect -8374 178718 -8138 178954
rect -8694 178398 -8458 178634
rect -8374 178398 -8138 178634
rect -8694 142718 -8458 142954
rect -8374 142718 -8138 142954
rect -8694 142398 -8458 142634
rect -8374 142398 -8138 142634
rect -8694 106718 -8458 106954
rect -8374 106718 -8138 106954
rect -8694 106398 -8458 106634
rect -8374 106398 -8138 106634
rect -8694 70718 -8458 70954
rect -8374 70718 -8138 70954
rect -8694 70398 -8458 70634
rect -8374 70398 -8138 70634
rect -8694 34718 -8458 34954
rect -8374 34718 -8138 34954
rect -8694 34398 -8458 34634
rect -8374 34398 -8138 34634
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 678218 -7498 678454
rect -7414 678218 -7178 678454
rect -7734 677898 -7498 678134
rect -7414 677898 -7178 678134
rect -7734 642218 -7498 642454
rect -7414 642218 -7178 642454
rect -7734 641898 -7498 642134
rect -7414 641898 -7178 642134
rect -7734 606218 -7498 606454
rect -7414 606218 -7178 606454
rect -7734 605898 -7498 606134
rect -7414 605898 -7178 606134
rect -7734 570218 -7498 570454
rect -7414 570218 -7178 570454
rect -7734 569898 -7498 570134
rect -7414 569898 -7178 570134
rect -7734 534218 -7498 534454
rect -7414 534218 -7178 534454
rect -7734 533898 -7498 534134
rect -7414 533898 -7178 534134
rect -7734 498218 -7498 498454
rect -7414 498218 -7178 498454
rect -7734 497898 -7498 498134
rect -7414 497898 -7178 498134
rect -7734 462218 -7498 462454
rect -7414 462218 -7178 462454
rect -7734 461898 -7498 462134
rect -7414 461898 -7178 462134
rect -7734 426218 -7498 426454
rect -7414 426218 -7178 426454
rect -7734 425898 -7498 426134
rect -7414 425898 -7178 426134
rect -7734 390218 -7498 390454
rect -7414 390218 -7178 390454
rect -7734 389898 -7498 390134
rect -7414 389898 -7178 390134
rect -7734 354218 -7498 354454
rect -7414 354218 -7178 354454
rect -7734 353898 -7498 354134
rect -7414 353898 -7178 354134
rect -7734 318218 -7498 318454
rect -7414 318218 -7178 318454
rect -7734 317898 -7498 318134
rect -7414 317898 -7178 318134
rect -7734 282218 -7498 282454
rect -7414 282218 -7178 282454
rect -7734 281898 -7498 282134
rect -7414 281898 -7178 282134
rect -7734 246218 -7498 246454
rect -7414 246218 -7178 246454
rect -7734 245898 -7498 246134
rect -7414 245898 -7178 246134
rect -7734 210218 -7498 210454
rect -7414 210218 -7178 210454
rect -7734 209898 -7498 210134
rect -7414 209898 -7178 210134
rect -7734 174218 -7498 174454
rect -7414 174218 -7178 174454
rect -7734 173898 -7498 174134
rect -7414 173898 -7178 174134
rect -7734 138218 -7498 138454
rect -7414 138218 -7178 138454
rect -7734 137898 -7498 138134
rect -7414 137898 -7178 138134
rect -7734 102218 -7498 102454
rect -7414 102218 -7178 102454
rect -7734 101898 -7498 102134
rect -7414 101898 -7178 102134
rect -7734 66218 -7498 66454
rect -7414 66218 -7178 66454
rect -7734 65898 -7498 66134
rect -7414 65898 -7178 66134
rect -7734 30218 -7498 30454
rect -7414 30218 -7178 30454
rect -7734 29898 -7498 30134
rect -7414 29898 -7178 30134
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 673718 -6538 673954
rect -6454 673718 -6218 673954
rect -6774 673398 -6538 673634
rect -6454 673398 -6218 673634
rect -6774 637718 -6538 637954
rect -6454 637718 -6218 637954
rect -6774 637398 -6538 637634
rect -6454 637398 -6218 637634
rect -6774 601718 -6538 601954
rect -6454 601718 -6218 601954
rect -6774 601398 -6538 601634
rect -6454 601398 -6218 601634
rect -6774 565718 -6538 565954
rect -6454 565718 -6218 565954
rect -6774 565398 -6538 565634
rect -6454 565398 -6218 565634
rect -6774 529718 -6538 529954
rect -6454 529718 -6218 529954
rect -6774 529398 -6538 529634
rect -6454 529398 -6218 529634
rect -6774 493718 -6538 493954
rect -6454 493718 -6218 493954
rect -6774 493398 -6538 493634
rect -6454 493398 -6218 493634
rect -6774 457718 -6538 457954
rect -6454 457718 -6218 457954
rect -6774 457398 -6538 457634
rect -6454 457398 -6218 457634
rect -6774 421718 -6538 421954
rect -6454 421718 -6218 421954
rect -6774 421398 -6538 421634
rect -6454 421398 -6218 421634
rect -6774 385718 -6538 385954
rect -6454 385718 -6218 385954
rect -6774 385398 -6538 385634
rect -6454 385398 -6218 385634
rect -6774 349718 -6538 349954
rect -6454 349718 -6218 349954
rect -6774 349398 -6538 349634
rect -6454 349398 -6218 349634
rect -6774 313718 -6538 313954
rect -6454 313718 -6218 313954
rect -6774 313398 -6538 313634
rect -6454 313398 -6218 313634
rect -6774 277718 -6538 277954
rect -6454 277718 -6218 277954
rect -6774 277398 -6538 277634
rect -6454 277398 -6218 277634
rect -6774 241718 -6538 241954
rect -6454 241718 -6218 241954
rect -6774 241398 -6538 241634
rect -6454 241398 -6218 241634
rect -6774 205718 -6538 205954
rect -6454 205718 -6218 205954
rect -6774 205398 -6538 205634
rect -6454 205398 -6218 205634
rect -6774 169718 -6538 169954
rect -6454 169718 -6218 169954
rect -6774 169398 -6538 169634
rect -6454 169398 -6218 169634
rect -6774 133718 -6538 133954
rect -6454 133718 -6218 133954
rect -6774 133398 -6538 133634
rect -6454 133398 -6218 133634
rect -6774 97718 -6538 97954
rect -6454 97718 -6218 97954
rect -6774 97398 -6538 97634
rect -6454 97398 -6218 97634
rect -6774 61718 -6538 61954
rect -6454 61718 -6218 61954
rect -6774 61398 -6538 61634
rect -6454 61398 -6218 61634
rect -6774 25718 -6538 25954
rect -6454 25718 -6218 25954
rect -6774 25398 -6538 25634
rect -6454 25398 -6218 25634
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 669218 -5578 669454
rect -5494 669218 -5258 669454
rect -5814 668898 -5578 669134
rect -5494 668898 -5258 669134
rect -5814 633218 -5578 633454
rect -5494 633218 -5258 633454
rect -5814 632898 -5578 633134
rect -5494 632898 -5258 633134
rect -5814 597218 -5578 597454
rect -5494 597218 -5258 597454
rect -5814 596898 -5578 597134
rect -5494 596898 -5258 597134
rect -5814 561218 -5578 561454
rect -5494 561218 -5258 561454
rect -5814 560898 -5578 561134
rect -5494 560898 -5258 561134
rect -5814 525218 -5578 525454
rect -5494 525218 -5258 525454
rect -5814 524898 -5578 525134
rect -5494 524898 -5258 525134
rect -5814 489218 -5578 489454
rect -5494 489218 -5258 489454
rect -5814 488898 -5578 489134
rect -5494 488898 -5258 489134
rect -5814 453218 -5578 453454
rect -5494 453218 -5258 453454
rect -5814 452898 -5578 453134
rect -5494 452898 -5258 453134
rect -5814 417218 -5578 417454
rect -5494 417218 -5258 417454
rect -5814 416898 -5578 417134
rect -5494 416898 -5258 417134
rect -5814 381218 -5578 381454
rect -5494 381218 -5258 381454
rect -5814 380898 -5578 381134
rect -5494 380898 -5258 381134
rect -5814 345218 -5578 345454
rect -5494 345218 -5258 345454
rect -5814 344898 -5578 345134
rect -5494 344898 -5258 345134
rect -5814 309218 -5578 309454
rect -5494 309218 -5258 309454
rect -5814 308898 -5578 309134
rect -5494 308898 -5258 309134
rect -5814 273218 -5578 273454
rect -5494 273218 -5258 273454
rect -5814 272898 -5578 273134
rect -5494 272898 -5258 273134
rect -5814 237218 -5578 237454
rect -5494 237218 -5258 237454
rect -5814 236898 -5578 237134
rect -5494 236898 -5258 237134
rect -5814 201218 -5578 201454
rect -5494 201218 -5258 201454
rect -5814 200898 -5578 201134
rect -5494 200898 -5258 201134
rect -5814 165218 -5578 165454
rect -5494 165218 -5258 165454
rect -5814 164898 -5578 165134
rect -5494 164898 -5258 165134
rect -5814 129218 -5578 129454
rect -5494 129218 -5258 129454
rect -5814 128898 -5578 129134
rect -5494 128898 -5258 129134
rect -5814 93218 -5578 93454
rect -5494 93218 -5258 93454
rect -5814 92898 -5578 93134
rect -5494 92898 -5258 93134
rect -5814 57218 -5578 57454
rect -5494 57218 -5258 57454
rect -5814 56898 -5578 57134
rect -5494 56898 -5258 57134
rect -5814 21218 -5578 21454
rect -5494 21218 -5258 21454
rect -5814 20898 -5578 21134
rect -5494 20898 -5258 21134
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 700718 -4618 700954
rect -4534 700718 -4298 700954
rect -4854 700398 -4618 700634
rect -4534 700398 -4298 700634
rect -4854 664718 -4618 664954
rect -4534 664718 -4298 664954
rect -4854 664398 -4618 664634
rect -4534 664398 -4298 664634
rect -4854 628718 -4618 628954
rect -4534 628718 -4298 628954
rect -4854 628398 -4618 628634
rect -4534 628398 -4298 628634
rect -4854 592718 -4618 592954
rect -4534 592718 -4298 592954
rect -4854 592398 -4618 592634
rect -4534 592398 -4298 592634
rect -4854 556718 -4618 556954
rect -4534 556718 -4298 556954
rect -4854 556398 -4618 556634
rect -4534 556398 -4298 556634
rect -4854 520718 -4618 520954
rect -4534 520718 -4298 520954
rect -4854 520398 -4618 520634
rect -4534 520398 -4298 520634
rect -4854 484718 -4618 484954
rect -4534 484718 -4298 484954
rect -4854 484398 -4618 484634
rect -4534 484398 -4298 484634
rect -4854 448718 -4618 448954
rect -4534 448718 -4298 448954
rect -4854 448398 -4618 448634
rect -4534 448398 -4298 448634
rect -4854 412718 -4618 412954
rect -4534 412718 -4298 412954
rect -4854 412398 -4618 412634
rect -4534 412398 -4298 412634
rect -4854 376718 -4618 376954
rect -4534 376718 -4298 376954
rect -4854 376398 -4618 376634
rect -4534 376398 -4298 376634
rect -4854 340718 -4618 340954
rect -4534 340718 -4298 340954
rect -4854 340398 -4618 340634
rect -4534 340398 -4298 340634
rect -4854 304718 -4618 304954
rect -4534 304718 -4298 304954
rect -4854 304398 -4618 304634
rect -4534 304398 -4298 304634
rect -4854 268718 -4618 268954
rect -4534 268718 -4298 268954
rect -4854 268398 -4618 268634
rect -4534 268398 -4298 268634
rect -4854 232718 -4618 232954
rect -4534 232718 -4298 232954
rect -4854 232398 -4618 232634
rect -4534 232398 -4298 232634
rect -4854 196718 -4618 196954
rect -4534 196718 -4298 196954
rect -4854 196398 -4618 196634
rect -4534 196398 -4298 196634
rect -4854 160718 -4618 160954
rect -4534 160718 -4298 160954
rect -4854 160398 -4618 160634
rect -4534 160398 -4298 160634
rect -4854 124718 -4618 124954
rect -4534 124718 -4298 124954
rect -4854 124398 -4618 124634
rect -4534 124398 -4298 124634
rect -4854 88718 -4618 88954
rect -4534 88718 -4298 88954
rect -4854 88398 -4618 88634
rect -4534 88398 -4298 88634
rect -4854 52718 -4618 52954
rect -4534 52718 -4298 52954
rect -4854 52398 -4618 52634
rect -4534 52398 -4298 52634
rect -4854 16718 -4618 16954
rect -4534 16718 -4298 16954
rect -4854 16398 -4618 16634
rect -4534 16398 -4298 16634
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 696218 -3658 696454
rect -3574 696218 -3338 696454
rect -3894 695898 -3658 696134
rect -3574 695898 -3338 696134
rect -3894 660218 -3658 660454
rect -3574 660218 -3338 660454
rect -3894 659898 -3658 660134
rect -3574 659898 -3338 660134
rect -3894 624218 -3658 624454
rect -3574 624218 -3338 624454
rect -3894 623898 -3658 624134
rect -3574 623898 -3338 624134
rect -3894 588218 -3658 588454
rect -3574 588218 -3338 588454
rect -3894 587898 -3658 588134
rect -3574 587898 -3338 588134
rect -3894 552218 -3658 552454
rect -3574 552218 -3338 552454
rect -3894 551898 -3658 552134
rect -3574 551898 -3338 552134
rect -3894 516218 -3658 516454
rect -3574 516218 -3338 516454
rect -3894 515898 -3658 516134
rect -3574 515898 -3338 516134
rect -3894 480218 -3658 480454
rect -3574 480218 -3338 480454
rect -3894 479898 -3658 480134
rect -3574 479898 -3338 480134
rect -3894 444218 -3658 444454
rect -3574 444218 -3338 444454
rect -3894 443898 -3658 444134
rect -3574 443898 -3338 444134
rect -3894 408218 -3658 408454
rect -3574 408218 -3338 408454
rect -3894 407898 -3658 408134
rect -3574 407898 -3338 408134
rect -3894 372218 -3658 372454
rect -3574 372218 -3338 372454
rect -3894 371898 -3658 372134
rect -3574 371898 -3338 372134
rect -3894 336218 -3658 336454
rect -3574 336218 -3338 336454
rect -3894 335898 -3658 336134
rect -3574 335898 -3338 336134
rect -3894 300218 -3658 300454
rect -3574 300218 -3338 300454
rect -3894 299898 -3658 300134
rect -3574 299898 -3338 300134
rect -3894 264218 -3658 264454
rect -3574 264218 -3338 264454
rect -3894 263898 -3658 264134
rect -3574 263898 -3338 264134
rect -3894 228218 -3658 228454
rect -3574 228218 -3338 228454
rect -3894 227898 -3658 228134
rect -3574 227898 -3338 228134
rect -3894 192218 -3658 192454
rect -3574 192218 -3338 192454
rect -3894 191898 -3658 192134
rect -3574 191898 -3338 192134
rect -3894 156218 -3658 156454
rect -3574 156218 -3338 156454
rect -3894 155898 -3658 156134
rect -3574 155898 -3338 156134
rect -3894 120218 -3658 120454
rect -3574 120218 -3338 120454
rect -3894 119898 -3658 120134
rect -3574 119898 -3338 120134
rect -3894 84218 -3658 84454
rect -3574 84218 -3338 84454
rect -3894 83898 -3658 84134
rect -3574 83898 -3338 84134
rect -3894 48218 -3658 48454
rect -3574 48218 -3338 48454
rect -3894 47898 -3658 48134
rect -3574 47898 -3338 48134
rect -3894 12218 -3658 12454
rect -3574 12218 -3338 12454
rect -3894 11898 -3658 12134
rect -3574 11898 -3338 12134
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 691718 -2698 691954
rect -2614 691718 -2378 691954
rect -2934 691398 -2698 691634
rect -2614 691398 -2378 691634
rect -2934 655718 -2698 655954
rect -2614 655718 -2378 655954
rect -2934 655398 -2698 655634
rect -2614 655398 -2378 655634
rect -2934 619718 -2698 619954
rect -2614 619718 -2378 619954
rect -2934 619398 -2698 619634
rect -2614 619398 -2378 619634
rect -2934 583718 -2698 583954
rect -2614 583718 -2378 583954
rect -2934 583398 -2698 583634
rect -2614 583398 -2378 583634
rect -2934 547718 -2698 547954
rect -2614 547718 -2378 547954
rect -2934 547398 -2698 547634
rect -2614 547398 -2378 547634
rect -2934 511718 -2698 511954
rect -2614 511718 -2378 511954
rect -2934 511398 -2698 511634
rect -2614 511398 -2378 511634
rect -2934 475718 -2698 475954
rect -2614 475718 -2378 475954
rect -2934 475398 -2698 475634
rect -2614 475398 -2378 475634
rect -2934 439718 -2698 439954
rect -2614 439718 -2378 439954
rect -2934 439398 -2698 439634
rect -2614 439398 -2378 439634
rect -2934 403718 -2698 403954
rect -2614 403718 -2378 403954
rect -2934 403398 -2698 403634
rect -2614 403398 -2378 403634
rect -2934 367718 -2698 367954
rect -2614 367718 -2378 367954
rect -2934 367398 -2698 367634
rect -2614 367398 -2378 367634
rect -2934 331718 -2698 331954
rect -2614 331718 -2378 331954
rect -2934 331398 -2698 331634
rect -2614 331398 -2378 331634
rect -2934 295718 -2698 295954
rect -2614 295718 -2378 295954
rect -2934 295398 -2698 295634
rect -2614 295398 -2378 295634
rect -2934 259718 -2698 259954
rect -2614 259718 -2378 259954
rect -2934 259398 -2698 259634
rect -2614 259398 -2378 259634
rect -2934 223718 -2698 223954
rect -2614 223718 -2378 223954
rect -2934 223398 -2698 223634
rect -2614 223398 -2378 223634
rect -2934 187718 -2698 187954
rect -2614 187718 -2378 187954
rect -2934 187398 -2698 187634
rect -2614 187398 -2378 187634
rect -2934 151718 -2698 151954
rect -2614 151718 -2378 151954
rect -2934 151398 -2698 151634
rect -2614 151398 -2378 151634
rect -2934 115718 -2698 115954
rect -2614 115718 -2378 115954
rect -2934 115398 -2698 115634
rect -2614 115398 -2378 115634
rect -2934 79718 -2698 79954
rect -2614 79718 -2378 79954
rect -2934 79398 -2698 79634
rect -2614 79398 -2378 79634
rect -2934 43718 -2698 43954
rect -2614 43718 -2378 43954
rect -2934 43398 -2698 43634
rect -2614 43398 -2378 43634
rect -2934 7718 -2698 7954
rect -2614 7718 -2378 7954
rect -2934 7398 -2698 7634
rect -2614 7398 -2378 7634
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 6326 705562 6562 705798
rect 6646 705562 6882 705798
rect 6326 705242 6562 705478
rect 6646 705242 6882 705478
rect 6326 691718 6562 691954
rect 6646 691718 6882 691954
rect 6326 691398 6562 691634
rect 6646 691398 6882 691634
rect 6326 655718 6562 655954
rect 6646 655718 6882 655954
rect 6326 655398 6562 655634
rect 6646 655398 6882 655634
rect 6326 619718 6562 619954
rect 6646 619718 6882 619954
rect 6326 619398 6562 619634
rect 6646 619398 6882 619634
rect 6326 583718 6562 583954
rect 6646 583718 6882 583954
rect 6326 583398 6562 583634
rect 6646 583398 6882 583634
rect 6326 547718 6562 547954
rect 6646 547718 6882 547954
rect 6326 547398 6562 547634
rect 6646 547398 6882 547634
rect 6326 511718 6562 511954
rect 6646 511718 6882 511954
rect 6326 511398 6562 511634
rect 6646 511398 6882 511634
rect 6326 475718 6562 475954
rect 6646 475718 6882 475954
rect 6326 475398 6562 475634
rect 6646 475398 6882 475634
rect 6326 439718 6562 439954
rect 6646 439718 6882 439954
rect 6326 439398 6562 439634
rect 6646 439398 6882 439634
rect 6326 403718 6562 403954
rect 6646 403718 6882 403954
rect 6326 403398 6562 403634
rect 6646 403398 6882 403634
rect 6326 367718 6562 367954
rect 6646 367718 6882 367954
rect 6326 367398 6562 367634
rect 6646 367398 6882 367634
rect 6326 331718 6562 331954
rect 6646 331718 6882 331954
rect 6326 331398 6562 331634
rect 6646 331398 6882 331634
rect 6326 295718 6562 295954
rect 6646 295718 6882 295954
rect 6326 295398 6562 295634
rect 6646 295398 6882 295634
rect 6326 259718 6562 259954
rect 6646 259718 6882 259954
rect 6326 259398 6562 259634
rect 6646 259398 6882 259634
rect 6326 223718 6562 223954
rect 6646 223718 6882 223954
rect 6326 223398 6562 223634
rect 6646 223398 6882 223634
rect 6326 187718 6562 187954
rect 6646 187718 6882 187954
rect 6326 187398 6562 187634
rect 6646 187398 6882 187634
rect 6326 151718 6562 151954
rect 6646 151718 6882 151954
rect 6326 151398 6562 151634
rect 6646 151398 6882 151634
rect 6326 115718 6562 115954
rect 6646 115718 6882 115954
rect 6326 115398 6562 115634
rect 6646 115398 6882 115634
rect 6326 79718 6562 79954
rect 6646 79718 6882 79954
rect 6326 79398 6562 79634
rect 6646 79398 6882 79634
rect 6326 43718 6562 43954
rect 6646 43718 6882 43954
rect 6326 43398 6562 43634
rect 6646 43398 6882 43634
rect 6326 7718 6562 7954
rect 6646 7718 6882 7954
rect 6326 7398 6562 7634
rect 6646 7398 6882 7634
rect 6326 -1542 6562 -1306
rect 6646 -1542 6882 -1306
rect 6326 -1862 6562 -1626
rect 6646 -1862 6882 -1626
rect 10826 706522 11062 706758
rect 11146 706522 11382 706758
rect 10826 706202 11062 706438
rect 11146 706202 11382 706438
rect 10826 696218 11062 696454
rect 11146 696218 11382 696454
rect 10826 695898 11062 696134
rect 11146 695898 11382 696134
rect 10826 660218 11062 660454
rect 11146 660218 11382 660454
rect 10826 659898 11062 660134
rect 11146 659898 11382 660134
rect 10826 624218 11062 624454
rect 11146 624218 11382 624454
rect 10826 623898 11062 624134
rect 11146 623898 11382 624134
rect 10826 588218 11062 588454
rect 11146 588218 11382 588454
rect 10826 587898 11062 588134
rect 11146 587898 11382 588134
rect 10826 552218 11062 552454
rect 11146 552218 11382 552454
rect 10826 551898 11062 552134
rect 11146 551898 11382 552134
rect 10826 516218 11062 516454
rect 11146 516218 11382 516454
rect 10826 515898 11062 516134
rect 11146 515898 11382 516134
rect 10826 480218 11062 480454
rect 11146 480218 11382 480454
rect 10826 479898 11062 480134
rect 11146 479898 11382 480134
rect 10826 444218 11062 444454
rect 11146 444218 11382 444454
rect 10826 443898 11062 444134
rect 11146 443898 11382 444134
rect 10826 408218 11062 408454
rect 11146 408218 11382 408454
rect 10826 407898 11062 408134
rect 11146 407898 11382 408134
rect 10826 372218 11062 372454
rect 11146 372218 11382 372454
rect 10826 371898 11062 372134
rect 11146 371898 11382 372134
rect 10826 336218 11062 336454
rect 11146 336218 11382 336454
rect 10826 335898 11062 336134
rect 11146 335898 11382 336134
rect 10826 300218 11062 300454
rect 11146 300218 11382 300454
rect 10826 299898 11062 300134
rect 11146 299898 11382 300134
rect 10826 264218 11062 264454
rect 11146 264218 11382 264454
rect 10826 263898 11062 264134
rect 11146 263898 11382 264134
rect 10826 228218 11062 228454
rect 11146 228218 11382 228454
rect 10826 227898 11062 228134
rect 11146 227898 11382 228134
rect 10826 192218 11062 192454
rect 11146 192218 11382 192454
rect 10826 191898 11062 192134
rect 11146 191898 11382 192134
rect 10826 156218 11062 156454
rect 11146 156218 11382 156454
rect 10826 155898 11062 156134
rect 11146 155898 11382 156134
rect 10826 120218 11062 120454
rect 11146 120218 11382 120454
rect 10826 119898 11062 120134
rect 11146 119898 11382 120134
rect 10826 84218 11062 84454
rect 11146 84218 11382 84454
rect 10826 83898 11062 84134
rect 11146 83898 11382 84134
rect 10826 48218 11062 48454
rect 11146 48218 11382 48454
rect 10826 47898 11062 48134
rect 11146 47898 11382 48134
rect 10826 12218 11062 12454
rect 11146 12218 11382 12454
rect 10826 11898 11062 12134
rect 11146 11898 11382 12134
rect 10826 -2502 11062 -2266
rect 11146 -2502 11382 -2266
rect 10826 -2822 11062 -2586
rect 11146 -2822 11382 -2586
rect 15326 707482 15562 707718
rect 15646 707482 15882 707718
rect 15326 707162 15562 707398
rect 15646 707162 15882 707398
rect 15326 700718 15562 700954
rect 15646 700718 15882 700954
rect 15326 700398 15562 700634
rect 15646 700398 15882 700634
rect 15326 664718 15562 664954
rect 15646 664718 15882 664954
rect 15326 664398 15562 664634
rect 15646 664398 15882 664634
rect 15326 628718 15562 628954
rect 15646 628718 15882 628954
rect 15326 628398 15562 628634
rect 15646 628398 15882 628634
rect 15326 592718 15562 592954
rect 15646 592718 15882 592954
rect 15326 592398 15562 592634
rect 15646 592398 15882 592634
rect 15326 556718 15562 556954
rect 15646 556718 15882 556954
rect 15326 556398 15562 556634
rect 15646 556398 15882 556634
rect 15326 520718 15562 520954
rect 15646 520718 15882 520954
rect 15326 520398 15562 520634
rect 15646 520398 15882 520634
rect 15326 484718 15562 484954
rect 15646 484718 15882 484954
rect 15326 484398 15562 484634
rect 15646 484398 15882 484634
rect 15326 448718 15562 448954
rect 15646 448718 15882 448954
rect 15326 448398 15562 448634
rect 15646 448398 15882 448634
rect 15326 412718 15562 412954
rect 15646 412718 15882 412954
rect 15326 412398 15562 412634
rect 15646 412398 15882 412634
rect 15326 376718 15562 376954
rect 15646 376718 15882 376954
rect 15326 376398 15562 376634
rect 15646 376398 15882 376634
rect 15326 340718 15562 340954
rect 15646 340718 15882 340954
rect 15326 340398 15562 340634
rect 15646 340398 15882 340634
rect 15326 304718 15562 304954
rect 15646 304718 15882 304954
rect 15326 304398 15562 304634
rect 15646 304398 15882 304634
rect 15326 268718 15562 268954
rect 15646 268718 15882 268954
rect 15326 268398 15562 268634
rect 15646 268398 15882 268634
rect 15326 232718 15562 232954
rect 15646 232718 15882 232954
rect 15326 232398 15562 232634
rect 15646 232398 15882 232634
rect 15326 196718 15562 196954
rect 15646 196718 15882 196954
rect 15326 196398 15562 196634
rect 15646 196398 15882 196634
rect 15326 160718 15562 160954
rect 15646 160718 15882 160954
rect 15326 160398 15562 160634
rect 15646 160398 15882 160634
rect 15326 124718 15562 124954
rect 15646 124718 15882 124954
rect 15326 124398 15562 124634
rect 15646 124398 15882 124634
rect 15326 88718 15562 88954
rect 15646 88718 15882 88954
rect 15326 88398 15562 88634
rect 15646 88398 15882 88634
rect 15326 52718 15562 52954
rect 15646 52718 15882 52954
rect 15326 52398 15562 52634
rect 15646 52398 15882 52634
rect 15326 16718 15562 16954
rect 15646 16718 15882 16954
rect 15326 16398 15562 16634
rect 15646 16398 15882 16634
rect 15326 -3462 15562 -3226
rect 15646 -3462 15882 -3226
rect 15326 -3782 15562 -3546
rect 15646 -3782 15882 -3546
rect 19826 708442 20062 708678
rect 20146 708442 20382 708678
rect 19826 708122 20062 708358
rect 20146 708122 20382 708358
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -4422 20062 -4186
rect 20146 -4422 20382 -4186
rect 19826 -4742 20062 -4506
rect 20146 -4742 20382 -4506
rect 24326 709402 24562 709638
rect 24646 709402 24882 709638
rect 24326 709082 24562 709318
rect 24646 709082 24882 709318
rect 24326 673718 24562 673954
rect 24646 673718 24882 673954
rect 24326 673398 24562 673634
rect 24646 673398 24882 673634
rect 24326 637718 24562 637954
rect 24646 637718 24882 637954
rect 24326 637398 24562 637634
rect 24646 637398 24882 637634
rect 24326 601718 24562 601954
rect 24646 601718 24882 601954
rect 24326 601398 24562 601634
rect 24646 601398 24882 601634
rect 24326 565718 24562 565954
rect 24646 565718 24882 565954
rect 24326 565398 24562 565634
rect 24646 565398 24882 565634
rect 24326 529718 24562 529954
rect 24646 529718 24882 529954
rect 24326 529398 24562 529634
rect 24646 529398 24882 529634
rect 24326 493718 24562 493954
rect 24646 493718 24882 493954
rect 24326 493398 24562 493634
rect 24646 493398 24882 493634
rect 24326 457718 24562 457954
rect 24646 457718 24882 457954
rect 24326 457398 24562 457634
rect 24646 457398 24882 457634
rect 24326 421718 24562 421954
rect 24646 421718 24882 421954
rect 24326 421398 24562 421634
rect 24646 421398 24882 421634
rect 24326 385718 24562 385954
rect 24646 385718 24882 385954
rect 24326 385398 24562 385634
rect 24646 385398 24882 385634
rect 24326 349718 24562 349954
rect 24646 349718 24882 349954
rect 24326 349398 24562 349634
rect 24646 349398 24882 349634
rect 24326 313718 24562 313954
rect 24646 313718 24882 313954
rect 24326 313398 24562 313634
rect 24646 313398 24882 313634
rect 24326 277718 24562 277954
rect 24646 277718 24882 277954
rect 24326 277398 24562 277634
rect 24646 277398 24882 277634
rect 24326 241718 24562 241954
rect 24646 241718 24882 241954
rect 24326 241398 24562 241634
rect 24646 241398 24882 241634
rect 24326 205718 24562 205954
rect 24646 205718 24882 205954
rect 24326 205398 24562 205634
rect 24646 205398 24882 205634
rect 24326 169718 24562 169954
rect 24646 169718 24882 169954
rect 24326 169398 24562 169634
rect 24646 169398 24882 169634
rect 24326 133718 24562 133954
rect 24646 133718 24882 133954
rect 24326 133398 24562 133634
rect 24646 133398 24882 133634
rect 24326 97718 24562 97954
rect 24646 97718 24882 97954
rect 24326 97398 24562 97634
rect 24646 97398 24882 97634
rect 24326 61718 24562 61954
rect 24646 61718 24882 61954
rect 24326 61398 24562 61634
rect 24646 61398 24882 61634
rect 24326 25718 24562 25954
rect 24646 25718 24882 25954
rect 24326 25398 24562 25634
rect 24646 25398 24882 25634
rect 24326 -5382 24562 -5146
rect 24646 -5382 24882 -5146
rect 24326 -5702 24562 -5466
rect 24646 -5702 24882 -5466
rect 28826 710362 29062 710598
rect 29146 710362 29382 710598
rect 28826 710042 29062 710278
rect 29146 710042 29382 710278
rect 28826 678218 29062 678454
rect 29146 678218 29382 678454
rect 28826 677898 29062 678134
rect 29146 677898 29382 678134
rect 28826 642218 29062 642454
rect 29146 642218 29382 642454
rect 28826 641898 29062 642134
rect 29146 641898 29382 642134
rect 28826 606218 29062 606454
rect 29146 606218 29382 606454
rect 28826 605898 29062 606134
rect 29146 605898 29382 606134
rect 28826 570218 29062 570454
rect 29146 570218 29382 570454
rect 28826 569898 29062 570134
rect 29146 569898 29382 570134
rect 28826 534218 29062 534454
rect 29146 534218 29382 534454
rect 28826 533898 29062 534134
rect 29146 533898 29382 534134
rect 28826 498218 29062 498454
rect 29146 498218 29382 498454
rect 28826 497898 29062 498134
rect 29146 497898 29382 498134
rect 28826 462218 29062 462454
rect 29146 462218 29382 462454
rect 28826 461898 29062 462134
rect 29146 461898 29382 462134
rect 28826 426218 29062 426454
rect 29146 426218 29382 426454
rect 28826 425898 29062 426134
rect 29146 425898 29382 426134
rect 28826 390218 29062 390454
rect 29146 390218 29382 390454
rect 28826 389898 29062 390134
rect 29146 389898 29382 390134
rect 28826 354218 29062 354454
rect 29146 354218 29382 354454
rect 28826 353898 29062 354134
rect 29146 353898 29382 354134
rect 28826 318218 29062 318454
rect 29146 318218 29382 318454
rect 28826 317898 29062 318134
rect 29146 317898 29382 318134
rect 28826 282218 29062 282454
rect 29146 282218 29382 282454
rect 28826 281898 29062 282134
rect 29146 281898 29382 282134
rect 28826 246218 29062 246454
rect 29146 246218 29382 246454
rect 28826 245898 29062 246134
rect 29146 245898 29382 246134
rect 28826 210218 29062 210454
rect 29146 210218 29382 210454
rect 28826 209898 29062 210134
rect 29146 209898 29382 210134
rect 28826 174218 29062 174454
rect 29146 174218 29382 174454
rect 28826 173898 29062 174134
rect 29146 173898 29382 174134
rect 28826 138218 29062 138454
rect 29146 138218 29382 138454
rect 28826 137898 29062 138134
rect 29146 137898 29382 138134
rect 28826 102218 29062 102454
rect 29146 102218 29382 102454
rect 28826 101898 29062 102134
rect 29146 101898 29382 102134
rect 28826 66218 29062 66454
rect 29146 66218 29382 66454
rect 28826 65898 29062 66134
rect 29146 65898 29382 66134
rect 28826 30218 29062 30454
rect 29146 30218 29382 30454
rect 28826 29898 29062 30134
rect 29146 29898 29382 30134
rect 28826 -6342 29062 -6106
rect 29146 -6342 29382 -6106
rect 28826 -6662 29062 -6426
rect 29146 -6662 29382 -6426
rect 33326 711322 33562 711558
rect 33646 711322 33882 711558
rect 33326 711002 33562 711238
rect 33646 711002 33882 711238
rect 33326 682718 33562 682954
rect 33646 682718 33882 682954
rect 33326 682398 33562 682634
rect 33646 682398 33882 682634
rect 33326 646718 33562 646954
rect 33646 646718 33882 646954
rect 33326 646398 33562 646634
rect 33646 646398 33882 646634
rect 33326 610718 33562 610954
rect 33646 610718 33882 610954
rect 33326 610398 33562 610634
rect 33646 610398 33882 610634
rect 33326 574718 33562 574954
rect 33646 574718 33882 574954
rect 33326 574398 33562 574634
rect 33646 574398 33882 574634
rect 33326 538718 33562 538954
rect 33646 538718 33882 538954
rect 33326 538398 33562 538634
rect 33646 538398 33882 538634
rect 33326 502718 33562 502954
rect 33646 502718 33882 502954
rect 33326 502398 33562 502634
rect 33646 502398 33882 502634
rect 33326 466718 33562 466954
rect 33646 466718 33882 466954
rect 33326 466398 33562 466634
rect 33646 466398 33882 466634
rect 33326 430718 33562 430954
rect 33646 430718 33882 430954
rect 33326 430398 33562 430634
rect 33646 430398 33882 430634
rect 33326 394718 33562 394954
rect 33646 394718 33882 394954
rect 33326 394398 33562 394634
rect 33646 394398 33882 394634
rect 33326 358718 33562 358954
rect 33646 358718 33882 358954
rect 33326 358398 33562 358634
rect 33646 358398 33882 358634
rect 33326 322718 33562 322954
rect 33646 322718 33882 322954
rect 33326 322398 33562 322634
rect 33646 322398 33882 322634
rect 33326 286718 33562 286954
rect 33646 286718 33882 286954
rect 33326 286398 33562 286634
rect 33646 286398 33882 286634
rect 33326 250718 33562 250954
rect 33646 250718 33882 250954
rect 33326 250398 33562 250634
rect 33646 250398 33882 250634
rect 33326 214718 33562 214954
rect 33646 214718 33882 214954
rect 33326 214398 33562 214634
rect 33646 214398 33882 214634
rect 33326 178718 33562 178954
rect 33646 178718 33882 178954
rect 33326 178398 33562 178634
rect 33646 178398 33882 178634
rect 33326 142718 33562 142954
rect 33646 142718 33882 142954
rect 33326 142398 33562 142634
rect 33646 142398 33882 142634
rect 33326 106718 33562 106954
rect 33646 106718 33882 106954
rect 33326 106398 33562 106634
rect 33646 106398 33882 106634
rect 33326 70718 33562 70954
rect 33646 70718 33882 70954
rect 33326 70398 33562 70634
rect 33646 70398 33882 70634
rect 33326 34718 33562 34954
rect 33646 34718 33882 34954
rect 33326 34398 33562 34634
rect 33646 34398 33882 34634
rect 33326 -7302 33562 -7066
rect 33646 -7302 33882 -7066
rect 33326 -7622 33562 -7386
rect 33646 -7622 33882 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 42326 705562 42562 705798
rect 42646 705562 42882 705798
rect 42326 705242 42562 705478
rect 42646 705242 42882 705478
rect 42326 691718 42562 691954
rect 42646 691718 42882 691954
rect 42326 691398 42562 691634
rect 42646 691398 42882 691634
rect 42326 655718 42562 655954
rect 42646 655718 42882 655954
rect 42326 655398 42562 655634
rect 42646 655398 42882 655634
rect 42326 619718 42562 619954
rect 42646 619718 42882 619954
rect 42326 619398 42562 619634
rect 42646 619398 42882 619634
rect 42326 583718 42562 583954
rect 42646 583718 42882 583954
rect 42326 583398 42562 583634
rect 42646 583398 42882 583634
rect 42326 547718 42562 547954
rect 42646 547718 42882 547954
rect 42326 547398 42562 547634
rect 42646 547398 42882 547634
rect 42326 511718 42562 511954
rect 42646 511718 42882 511954
rect 42326 511398 42562 511634
rect 42646 511398 42882 511634
rect 42326 475718 42562 475954
rect 42646 475718 42882 475954
rect 42326 475398 42562 475634
rect 42646 475398 42882 475634
rect 42326 439718 42562 439954
rect 42646 439718 42882 439954
rect 42326 439398 42562 439634
rect 42646 439398 42882 439634
rect 42326 403718 42562 403954
rect 42646 403718 42882 403954
rect 42326 403398 42562 403634
rect 42646 403398 42882 403634
rect 42326 367718 42562 367954
rect 42646 367718 42882 367954
rect 42326 367398 42562 367634
rect 42646 367398 42882 367634
rect 42326 331718 42562 331954
rect 42646 331718 42882 331954
rect 42326 331398 42562 331634
rect 42646 331398 42882 331634
rect 42326 295718 42562 295954
rect 42646 295718 42882 295954
rect 42326 295398 42562 295634
rect 42646 295398 42882 295634
rect 42326 259718 42562 259954
rect 42646 259718 42882 259954
rect 42326 259398 42562 259634
rect 42646 259398 42882 259634
rect 46826 706522 47062 706758
rect 47146 706522 47382 706758
rect 46826 706202 47062 706438
rect 47146 706202 47382 706438
rect 46826 696218 47062 696454
rect 47146 696218 47382 696454
rect 46826 695898 47062 696134
rect 47146 695898 47382 696134
rect 46826 660218 47062 660454
rect 47146 660218 47382 660454
rect 46826 659898 47062 660134
rect 47146 659898 47382 660134
rect 46826 624218 47062 624454
rect 47146 624218 47382 624454
rect 46826 623898 47062 624134
rect 47146 623898 47382 624134
rect 46826 588218 47062 588454
rect 47146 588218 47382 588454
rect 46826 587898 47062 588134
rect 47146 587898 47382 588134
rect 46826 552218 47062 552454
rect 47146 552218 47382 552454
rect 46826 551898 47062 552134
rect 47146 551898 47382 552134
rect 46826 516218 47062 516454
rect 47146 516218 47382 516454
rect 46826 515898 47062 516134
rect 47146 515898 47382 516134
rect 46826 480218 47062 480454
rect 47146 480218 47382 480454
rect 46826 479898 47062 480134
rect 47146 479898 47382 480134
rect 46826 444218 47062 444454
rect 47146 444218 47382 444454
rect 46826 443898 47062 444134
rect 47146 443898 47382 444134
rect 46826 408218 47062 408454
rect 47146 408218 47382 408454
rect 46826 407898 47062 408134
rect 47146 407898 47382 408134
rect 46826 372218 47062 372454
rect 47146 372218 47382 372454
rect 46826 371898 47062 372134
rect 47146 371898 47382 372134
rect 46826 336218 47062 336454
rect 47146 336218 47382 336454
rect 46826 335898 47062 336134
rect 47146 335898 47382 336134
rect 46826 300218 47062 300454
rect 47146 300218 47382 300454
rect 46826 299898 47062 300134
rect 47146 299898 47382 300134
rect 46826 264218 47062 264454
rect 47146 264218 47382 264454
rect 46826 263898 47062 264134
rect 47146 263898 47382 264134
rect 51326 707482 51562 707718
rect 51646 707482 51882 707718
rect 51326 707162 51562 707398
rect 51646 707162 51882 707398
rect 51326 700718 51562 700954
rect 51646 700718 51882 700954
rect 51326 700398 51562 700634
rect 51646 700398 51882 700634
rect 51326 664718 51562 664954
rect 51646 664718 51882 664954
rect 51326 664398 51562 664634
rect 51646 664398 51882 664634
rect 51326 628718 51562 628954
rect 51646 628718 51882 628954
rect 51326 628398 51562 628634
rect 51646 628398 51882 628634
rect 51326 592718 51562 592954
rect 51646 592718 51882 592954
rect 51326 592398 51562 592634
rect 51646 592398 51882 592634
rect 51326 556718 51562 556954
rect 51646 556718 51882 556954
rect 51326 556398 51562 556634
rect 51646 556398 51882 556634
rect 51326 520718 51562 520954
rect 51646 520718 51882 520954
rect 51326 520398 51562 520634
rect 51646 520398 51882 520634
rect 51326 484718 51562 484954
rect 51646 484718 51882 484954
rect 51326 484398 51562 484634
rect 51646 484398 51882 484634
rect 51326 448718 51562 448954
rect 51646 448718 51882 448954
rect 51326 448398 51562 448634
rect 51646 448398 51882 448634
rect 51326 412718 51562 412954
rect 51646 412718 51882 412954
rect 51326 412398 51562 412634
rect 51646 412398 51882 412634
rect 51326 376718 51562 376954
rect 51646 376718 51882 376954
rect 51326 376398 51562 376634
rect 51646 376398 51882 376634
rect 51326 340718 51562 340954
rect 51646 340718 51882 340954
rect 51326 340398 51562 340634
rect 51646 340398 51882 340634
rect 51326 304718 51562 304954
rect 51646 304718 51882 304954
rect 51326 304398 51562 304634
rect 51646 304398 51882 304634
rect 51326 268718 51562 268954
rect 51646 268718 51882 268954
rect 51326 268398 51562 268634
rect 51646 268398 51882 268634
rect 55826 708442 56062 708678
rect 56146 708442 56382 708678
rect 55826 708122 56062 708358
rect 56146 708122 56382 708358
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 60326 709402 60562 709638
rect 60646 709402 60882 709638
rect 60326 709082 60562 709318
rect 60646 709082 60882 709318
rect 60326 673718 60562 673954
rect 60646 673718 60882 673954
rect 60326 673398 60562 673634
rect 60646 673398 60882 673634
rect 60326 637718 60562 637954
rect 60646 637718 60882 637954
rect 60326 637398 60562 637634
rect 60646 637398 60882 637634
rect 60326 601718 60562 601954
rect 60646 601718 60882 601954
rect 60326 601398 60562 601634
rect 60646 601398 60882 601634
rect 60326 565718 60562 565954
rect 60646 565718 60882 565954
rect 60326 565398 60562 565634
rect 60646 565398 60882 565634
rect 60326 529718 60562 529954
rect 60646 529718 60882 529954
rect 60326 529398 60562 529634
rect 60646 529398 60882 529634
rect 60326 493718 60562 493954
rect 60646 493718 60882 493954
rect 60326 493398 60562 493634
rect 60646 493398 60882 493634
rect 60326 457718 60562 457954
rect 60646 457718 60882 457954
rect 60326 457398 60562 457634
rect 60646 457398 60882 457634
rect 60326 421718 60562 421954
rect 60646 421718 60882 421954
rect 60326 421398 60562 421634
rect 60646 421398 60882 421634
rect 60326 385718 60562 385954
rect 60646 385718 60882 385954
rect 60326 385398 60562 385634
rect 60646 385398 60882 385634
rect 60326 349718 60562 349954
rect 60646 349718 60882 349954
rect 60326 349398 60562 349634
rect 60646 349398 60882 349634
rect 60326 313718 60562 313954
rect 60646 313718 60882 313954
rect 60326 313398 60562 313634
rect 60646 313398 60882 313634
rect 60326 277718 60562 277954
rect 60646 277718 60882 277954
rect 60326 277398 60562 277634
rect 60646 277398 60882 277634
rect 64826 710362 65062 710598
rect 65146 710362 65382 710598
rect 64826 710042 65062 710278
rect 65146 710042 65382 710278
rect 64826 678218 65062 678454
rect 65146 678218 65382 678454
rect 64826 677898 65062 678134
rect 65146 677898 65382 678134
rect 64826 642218 65062 642454
rect 65146 642218 65382 642454
rect 64826 641898 65062 642134
rect 65146 641898 65382 642134
rect 64826 606218 65062 606454
rect 65146 606218 65382 606454
rect 64826 605898 65062 606134
rect 65146 605898 65382 606134
rect 64826 570218 65062 570454
rect 65146 570218 65382 570454
rect 64826 569898 65062 570134
rect 65146 569898 65382 570134
rect 64826 534218 65062 534454
rect 65146 534218 65382 534454
rect 64826 533898 65062 534134
rect 65146 533898 65382 534134
rect 64826 498218 65062 498454
rect 65146 498218 65382 498454
rect 64826 497898 65062 498134
rect 65146 497898 65382 498134
rect 64826 462218 65062 462454
rect 65146 462218 65382 462454
rect 64826 461898 65062 462134
rect 65146 461898 65382 462134
rect 64826 426218 65062 426454
rect 65146 426218 65382 426454
rect 64826 425898 65062 426134
rect 65146 425898 65382 426134
rect 64826 390218 65062 390454
rect 65146 390218 65382 390454
rect 64826 389898 65062 390134
rect 65146 389898 65382 390134
rect 64826 354218 65062 354454
rect 65146 354218 65382 354454
rect 64826 353898 65062 354134
rect 65146 353898 65382 354134
rect 64826 318218 65062 318454
rect 65146 318218 65382 318454
rect 64826 317898 65062 318134
rect 65146 317898 65382 318134
rect 64826 282218 65062 282454
rect 65146 282218 65382 282454
rect 64826 281898 65062 282134
rect 65146 281898 65382 282134
rect 64826 246218 65062 246454
rect 65146 246218 65382 246454
rect 64826 245898 65062 246134
rect 65146 245898 65382 246134
rect 69326 711322 69562 711558
rect 69646 711322 69882 711558
rect 69326 711002 69562 711238
rect 69646 711002 69882 711238
rect 69326 682718 69562 682954
rect 69646 682718 69882 682954
rect 69326 682398 69562 682634
rect 69646 682398 69882 682634
rect 69326 646718 69562 646954
rect 69646 646718 69882 646954
rect 69326 646398 69562 646634
rect 69646 646398 69882 646634
rect 69326 610718 69562 610954
rect 69646 610718 69882 610954
rect 69326 610398 69562 610634
rect 69646 610398 69882 610634
rect 69326 574718 69562 574954
rect 69646 574718 69882 574954
rect 69326 574398 69562 574634
rect 69646 574398 69882 574634
rect 69326 538718 69562 538954
rect 69646 538718 69882 538954
rect 69326 538398 69562 538634
rect 69646 538398 69882 538634
rect 69326 502718 69562 502954
rect 69646 502718 69882 502954
rect 69326 502398 69562 502634
rect 69646 502398 69882 502634
rect 69326 466718 69562 466954
rect 69646 466718 69882 466954
rect 69326 466398 69562 466634
rect 69646 466398 69882 466634
rect 69326 430718 69562 430954
rect 69646 430718 69882 430954
rect 69326 430398 69562 430634
rect 69646 430398 69882 430634
rect 69326 394718 69562 394954
rect 69646 394718 69882 394954
rect 69326 394398 69562 394634
rect 69646 394398 69882 394634
rect 69326 358718 69562 358954
rect 69646 358718 69882 358954
rect 69326 358398 69562 358634
rect 69646 358398 69882 358634
rect 69326 322718 69562 322954
rect 69646 322718 69882 322954
rect 69326 322398 69562 322634
rect 69646 322398 69882 322634
rect 69326 286718 69562 286954
rect 69646 286718 69882 286954
rect 69326 286398 69562 286634
rect 69646 286398 69882 286634
rect 69326 250718 69562 250954
rect 69646 250718 69882 250954
rect 69326 250398 69562 250634
rect 69646 250398 69882 250634
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 78326 705562 78562 705798
rect 78646 705562 78882 705798
rect 78326 705242 78562 705478
rect 78646 705242 78882 705478
rect 78326 691718 78562 691954
rect 78646 691718 78882 691954
rect 78326 691398 78562 691634
rect 78646 691398 78882 691634
rect 78326 655718 78562 655954
rect 78646 655718 78882 655954
rect 78326 655398 78562 655634
rect 78646 655398 78882 655634
rect 78326 619718 78562 619954
rect 78646 619718 78882 619954
rect 78326 619398 78562 619634
rect 78646 619398 78882 619634
rect 78326 583718 78562 583954
rect 78646 583718 78882 583954
rect 78326 583398 78562 583634
rect 78646 583398 78882 583634
rect 78326 547718 78562 547954
rect 78646 547718 78882 547954
rect 78326 547398 78562 547634
rect 78646 547398 78882 547634
rect 78326 511718 78562 511954
rect 78646 511718 78882 511954
rect 78326 511398 78562 511634
rect 78646 511398 78882 511634
rect 78326 475718 78562 475954
rect 78646 475718 78882 475954
rect 78326 475398 78562 475634
rect 78646 475398 78882 475634
rect 78326 439718 78562 439954
rect 78646 439718 78882 439954
rect 78326 439398 78562 439634
rect 78646 439398 78882 439634
rect 78326 403718 78562 403954
rect 78646 403718 78882 403954
rect 78326 403398 78562 403634
rect 78646 403398 78882 403634
rect 78326 367718 78562 367954
rect 78646 367718 78882 367954
rect 78326 367398 78562 367634
rect 78646 367398 78882 367634
rect 78326 331718 78562 331954
rect 78646 331718 78882 331954
rect 78326 331398 78562 331634
rect 78646 331398 78882 331634
rect 78326 295718 78562 295954
rect 78646 295718 78882 295954
rect 78326 295398 78562 295634
rect 78646 295398 78882 295634
rect 78326 259718 78562 259954
rect 78646 259718 78882 259954
rect 78326 259398 78562 259634
rect 78646 259398 78882 259634
rect 82826 706522 83062 706758
rect 83146 706522 83382 706758
rect 82826 706202 83062 706438
rect 83146 706202 83382 706438
rect 82826 696218 83062 696454
rect 83146 696218 83382 696454
rect 82826 695898 83062 696134
rect 83146 695898 83382 696134
rect 82826 660218 83062 660454
rect 83146 660218 83382 660454
rect 82826 659898 83062 660134
rect 83146 659898 83382 660134
rect 82826 624218 83062 624454
rect 83146 624218 83382 624454
rect 82826 623898 83062 624134
rect 83146 623898 83382 624134
rect 82826 588218 83062 588454
rect 83146 588218 83382 588454
rect 82826 587898 83062 588134
rect 83146 587898 83382 588134
rect 82826 552218 83062 552454
rect 83146 552218 83382 552454
rect 82826 551898 83062 552134
rect 83146 551898 83382 552134
rect 82826 516218 83062 516454
rect 83146 516218 83382 516454
rect 82826 515898 83062 516134
rect 83146 515898 83382 516134
rect 82826 480218 83062 480454
rect 83146 480218 83382 480454
rect 82826 479898 83062 480134
rect 83146 479898 83382 480134
rect 82826 444218 83062 444454
rect 83146 444218 83382 444454
rect 82826 443898 83062 444134
rect 83146 443898 83382 444134
rect 82826 408218 83062 408454
rect 83146 408218 83382 408454
rect 82826 407898 83062 408134
rect 83146 407898 83382 408134
rect 82826 372218 83062 372454
rect 83146 372218 83382 372454
rect 82826 371898 83062 372134
rect 83146 371898 83382 372134
rect 82826 336218 83062 336454
rect 83146 336218 83382 336454
rect 82826 335898 83062 336134
rect 83146 335898 83382 336134
rect 82826 300218 83062 300454
rect 83146 300218 83382 300454
rect 82826 299898 83062 300134
rect 83146 299898 83382 300134
rect 82826 264218 83062 264454
rect 83146 264218 83382 264454
rect 82826 263898 83062 264134
rect 83146 263898 83382 264134
rect 87326 707482 87562 707718
rect 87646 707482 87882 707718
rect 87326 707162 87562 707398
rect 87646 707162 87882 707398
rect 87326 700718 87562 700954
rect 87646 700718 87882 700954
rect 87326 700398 87562 700634
rect 87646 700398 87882 700634
rect 87326 664718 87562 664954
rect 87646 664718 87882 664954
rect 87326 664398 87562 664634
rect 87646 664398 87882 664634
rect 87326 628718 87562 628954
rect 87646 628718 87882 628954
rect 87326 628398 87562 628634
rect 87646 628398 87882 628634
rect 87326 592718 87562 592954
rect 87646 592718 87882 592954
rect 87326 592398 87562 592634
rect 87646 592398 87882 592634
rect 87326 556718 87562 556954
rect 87646 556718 87882 556954
rect 87326 556398 87562 556634
rect 87646 556398 87882 556634
rect 87326 520718 87562 520954
rect 87646 520718 87882 520954
rect 87326 520398 87562 520634
rect 87646 520398 87882 520634
rect 87326 484718 87562 484954
rect 87646 484718 87882 484954
rect 87326 484398 87562 484634
rect 87646 484398 87882 484634
rect 87326 448718 87562 448954
rect 87646 448718 87882 448954
rect 87326 448398 87562 448634
rect 87646 448398 87882 448634
rect 87326 412718 87562 412954
rect 87646 412718 87882 412954
rect 87326 412398 87562 412634
rect 87646 412398 87882 412634
rect 87326 376718 87562 376954
rect 87646 376718 87882 376954
rect 87326 376398 87562 376634
rect 87646 376398 87882 376634
rect 87326 340718 87562 340954
rect 87646 340718 87882 340954
rect 87326 340398 87562 340634
rect 87646 340398 87882 340634
rect 87326 304718 87562 304954
rect 87646 304718 87882 304954
rect 87326 304398 87562 304634
rect 87646 304398 87882 304634
rect 87326 268718 87562 268954
rect 87646 268718 87882 268954
rect 87326 268398 87562 268634
rect 87646 268398 87882 268634
rect 91826 708442 92062 708678
rect 92146 708442 92382 708678
rect 91826 708122 92062 708358
rect 92146 708122 92382 708358
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 96326 709402 96562 709638
rect 96646 709402 96882 709638
rect 96326 709082 96562 709318
rect 96646 709082 96882 709318
rect 96326 673718 96562 673954
rect 96646 673718 96882 673954
rect 96326 673398 96562 673634
rect 96646 673398 96882 673634
rect 96326 637718 96562 637954
rect 96646 637718 96882 637954
rect 96326 637398 96562 637634
rect 96646 637398 96882 637634
rect 96326 601718 96562 601954
rect 96646 601718 96882 601954
rect 96326 601398 96562 601634
rect 96646 601398 96882 601634
rect 96326 565718 96562 565954
rect 96646 565718 96882 565954
rect 96326 565398 96562 565634
rect 96646 565398 96882 565634
rect 96326 529718 96562 529954
rect 96646 529718 96882 529954
rect 96326 529398 96562 529634
rect 96646 529398 96882 529634
rect 96326 493718 96562 493954
rect 96646 493718 96882 493954
rect 96326 493398 96562 493634
rect 96646 493398 96882 493634
rect 96326 457718 96562 457954
rect 96646 457718 96882 457954
rect 96326 457398 96562 457634
rect 96646 457398 96882 457634
rect 96326 421718 96562 421954
rect 96646 421718 96882 421954
rect 96326 421398 96562 421634
rect 96646 421398 96882 421634
rect 96326 385718 96562 385954
rect 96646 385718 96882 385954
rect 96326 385398 96562 385634
rect 96646 385398 96882 385634
rect 96326 349718 96562 349954
rect 96646 349718 96882 349954
rect 96326 349398 96562 349634
rect 96646 349398 96882 349634
rect 96326 313718 96562 313954
rect 96646 313718 96882 313954
rect 96326 313398 96562 313634
rect 96646 313398 96882 313634
rect 96326 277718 96562 277954
rect 96646 277718 96882 277954
rect 96326 277398 96562 277634
rect 96646 277398 96882 277634
rect 100826 710362 101062 710598
rect 101146 710362 101382 710598
rect 100826 710042 101062 710278
rect 101146 710042 101382 710278
rect 100826 678218 101062 678454
rect 101146 678218 101382 678454
rect 100826 677898 101062 678134
rect 101146 677898 101382 678134
rect 100826 642218 101062 642454
rect 101146 642218 101382 642454
rect 100826 641898 101062 642134
rect 101146 641898 101382 642134
rect 100826 606218 101062 606454
rect 101146 606218 101382 606454
rect 100826 605898 101062 606134
rect 101146 605898 101382 606134
rect 100826 570218 101062 570454
rect 101146 570218 101382 570454
rect 100826 569898 101062 570134
rect 101146 569898 101382 570134
rect 100826 534218 101062 534454
rect 101146 534218 101382 534454
rect 100826 533898 101062 534134
rect 101146 533898 101382 534134
rect 100826 498218 101062 498454
rect 101146 498218 101382 498454
rect 100826 497898 101062 498134
rect 101146 497898 101382 498134
rect 100826 462218 101062 462454
rect 101146 462218 101382 462454
rect 100826 461898 101062 462134
rect 101146 461898 101382 462134
rect 100826 426218 101062 426454
rect 101146 426218 101382 426454
rect 100826 425898 101062 426134
rect 101146 425898 101382 426134
rect 100826 390218 101062 390454
rect 101146 390218 101382 390454
rect 100826 389898 101062 390134
rect 101146 389898 101382 390134
rect 100826 354218 101062 354454
rect 101146 354218 101382 354454
rect 100826 353898 101062 354134
rect 101146 353898 101382 354134
rect 100826 318218 101062 318454
rect 101146 318218 101382 318454
rect 100826 317898 101062 318134
rect 101146 317898 101382 318134
rect 100826 282218 101062 282454
rect 101146 282218 101382 282454
rect 100826 281898 101062 282134
rect 101146 281898 101382 282134
rect 100826 246218 101062 246454
rect 101146 246218 101382 246454
rect 100826 245898 101062 246134
rect 101146 245898 101382 246134
rect 105326 711322 105562 711558
rect 105646 711322 105882 711558
rect 105326 711002 105562 711238
rect 105646 711002 105882 711238
rect 105326 682718 105562 682954
rect 105646 682718 105882 682954
rect 105326 682398 105562 682634
rect 105646 682398 105882 682634
rect 105326 646718 105562 646954
rect 105646 646718 105882 646954
rect 105326 646398 105562 646634
rect 105646 646398 105882 646634
rect 105326 610718 105562 610954
rect 105646 610718 105882 610954
rect 105326 610398 105562 610634
rect 105646 610398 105882 610634
rect 105326 574718 105562 574954
rect 105646 574718 105882 574954
rect 105326 574398 105562 574634
rect 105646 574398 105882 574634
rect 105326 538718 105562 538954
rect 105646 538718 105882 538954
rect 105326 538398 105562 538634
rect 105646 538398 105882 538634
rect 105326 502718 105562 502954
rect 105646 502718 105882 502954
rect 105326 502398 105562 502634
rect 105646 502398 105882 502634
rect 105326 466718 105562 466954
rect 105646 466718 105882 466954
rect 105326 466398 105562 466634
rect 105646 466398 105882 466634
rect 105326 430718 105562 430954
rect 105646 430718 105882 430954
rect 105326 430398 105562 430634
rect 105646 430398 105882 430634
rect 105326 394718 105562 394954
rect 105646 394718 105882 394954
rect 105326 394398 105562 394634
rect 105646 394398 105882 394634
rect 105326 358718 105562 358954
rect 105646 358718 105882 358954
rect 105326 358398 105562 358634
rect 105646 358398 105882 358634
rect 105326 322718 105562 322954
rect 105646 322718 105882 322954
rect 105326 322398 105562 322634
rect 105646 322398 105882 322634
rect 105326 286718 105562 286954
rect 105646 286718 105882 286954
rect 105326 286398 105562 286634
rect 105646 286398 105882 286634
rect 105326 250718 105562 250954
rect 105646 250718 105882 250954
rect 105326 250398 105562 250634
rect 105646 250398 105882 250634
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 114326 705562 114562 705798
rect 114646 705562 114882 705798
rect 114326 705242 114562 705478
rect 114646 705242 114882 705478
rect 114326 691718 114562 691954
rect 114646 691718 114882 691954
rect 114326 691398 114562 691634
rect 114646 691398 114882 691634
rect 114326 655718 114562 655954
rect 114646 655718 114882 655954
rect 114326 655398 114562 655634
rect 114646 655398 114882 655634
rect 114326 619718 114562 619954
rect 114646 619718 114882 619954
rect 114326 619398 114562 619634
rect 114646 619398 114882 619634
rect 114326 583718 114562 583954
rect 114646 583718 114882 583954
rect 114326 583398 114562 583634
rect 114646 583398 114882 583634
rect 114326 547718 114562 547954
rect 114646 547718 114882 547954
rect 114326 547398 114562 547634
rect 114646 547398 114882 547634
rect 114326 511718 114562 511954
rect 114646 511718 114882 511954
rect 114326 511398 114562 511634
rect 114646 511398 114882 511634
rect 114326 475718 114562 475954
rect 114646 475718 114882 475954
rect 114326 475398 114562 475634
rect 114646 475398 114882 475634
rect 114326 439718 114562 439954
rect 114646 439718 114882 439954
rect 114326 439398 114562 439634
rect 114646 439398 114882 439634
rect 114326 403718 114562 403954
rect 114646 403718 114882 403954
rect 114326 403398 114562 403634
rect 114646 403398 114882 403634
rect 114326 367718 114562 367954
rect 114646 367718 114882 367954
rect 114326 367398 114562 367634
rect 114646 367398 114882 367634
rect 114326 331718 114562 331954
rect 114646 331718 114882 331954
rect 114326 331398 114562 331634
rect 114646 331398 114882 331634
rect 114326 295718 114562 295954
rect 114646 295718 114882 295954
rect 114326 295398 114562 295634
rect 114646 295398 114882 295634
rect 114326 259718 114562 259954
rect 114646 259718 114882 259954
rect 114326 259398 114562 259634
rect 114646 259398 114882 259634
rect 118826 706522 119062 706758
rect 119146 706522 119382 706758
rect 118826 706202 119062 706438
rect 119146 706202 119382 706438
rect 118826 696218 119062 696454
rect 119146 696218 119382 696454
rect 118826 695898 119062 696134
rect 119146 695898 119382 696134
rect 118826 660218 119062 660454
rect 119146 660218 119382 660454
rect 118826 659898 119062 660134
rect 119146 659898 119382 660134
rect 118826 624218 119062 624454
rect 119146 624218 119382 624454
rect 118826 623898 119062 624134
rect 119146 623898 119382 624134
rect 118826 588218 119062 588454
rect 119146 588218 119382 588454
rect 118826 587898 119062 588134
rect 119146 587898 119382 588134
rect 118826 552218 119062 552454
rect 119146 552218 119382 552454
rect 118826 551898 119062 552134
rect 119146 551898 119382 552134
rect 118826 516218 119062 516454
rect 119146 516218 119382 516454
rect 118826 515898 119062 516134
rect 119146 515898 119382 516134
rect 118826 480218 119062 480454
rect 119146 480218 119382 480454
rect 118826 479898 119062 480134
rect 119146 479898 119382 480134
rect 118826 444218 119062 444454
rect 119146 444218 119382 444454
rect 118826 443898 119062 444134
rect 119146 443898 119382 444134
rect 118826 408218 119062 408454
rect 119146 408218 119382 408454
rect 118826 407898 119062 408134
rect 119146 407898 119382 408134
rect 118826 372218 119062 372454
rect 119146 372218 119382 372454
rect 118826 371898 119062 372134
rect 119146 371898 119382 372134
rect 118826 336218 119062 336454
rect 119146 336218 119382 336454
rect 118826 335898 119062 336134
rect 119146 335898 119382 336134
rect 118826 300218 119062 300454
rect 119146 300218 119382 300454
rect 118826 299898 119062 300134
rect 119146 299898 119382 300134
rect 118826 264218 119062 264454
rect 119146 264218 119382 264454
rect 118826 263898 119062 264134
rect 119146 263898 119382 264134
rect 123326 707482 123562 707718
rect 123646 707482 123882 707718
rect 123326 707162 123562 707398
rect 123646 707162 123882 707398
rect 123326 700718 123562 700954
rect 123646 700718 123882 700954
rect 123326 700398 123562 700634
rect 123646 700398 123882 700634
rect 123326 664718 123562 664954
rect 123646 664718 123882 664954
rect 123326 664398 123562 664634
rect 123646 664398 123882 664634
rect 123326 628718 123562 628954
rect 123646 628718 123882 628954
rect 123326 628398 123562 628634
rect 123646 628398 123882 628634
rect 123326 592718 123562 592954
rect 123646 592718 123882 592954
rect 123326 592398 123562 592634
rect 123646 592398 123882 592634
rect 123326 556718 123562 556954
rect 123646 556718 123882 556954
rect 123326 556398 123562 556634
rect 123646 556398 123882 556634
rect 123326 520718 123562 520954
rect 123646 520718 123882 520954
rect 123326 520398 123562 520634
rect 123646 520398 123882 520634
rect 123326 484718 123562 484954
rect 123646 484718 123882 484954
rect 123326 484398 123562 484634
rect 123646 484398 123882 484634
rect 123326 448718 123562 448954
rect 123646 448718 123882 448954
rect 123326 448398 123562 448634
rect 123646 448398 123882 448634
rect 123326 412718 123562 412954
rect 123646 412718 123882 412954
rect 123326 412398 123562 412634
rect 123646 412398 123882 412634
rect 123326 376718 123562 376954
rect 123646 376718 123882 376954
rect 123326 376398 123562 376634
rect 123646 376398 123882 376634
rect 123326 340718 123562 340954
rect 123646 340718 123882 340954
rect 123326 340398 123562 340634
rect 123646 340398 123882 340634
rect 123326 304718 123562 304954
rect 123646 304718 123882 304954
rect 123326 304398 123562 304634
rect 123646 304398 123882 304634
rect 123326 268718 123562 268954
rect 123646 268718 123882 268954
rect 123326 268398 123562 268634
rect 123646 268398 123882 268634
rect 127826 708442 128062 708678
rect 128146 708442 128382 708678
rect 127826 708122 128062 708358
rect 128146 708122 128382 708358
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 132326 709402 132562 709638
rect 132646 709402 132882 709638
rect 132326 709082 132562 709318
rect 132646 709082 132882 709318
rect 132326 673718 132562 673954
rect 132646 673718 132882 673954
rect 132326 673398 132562 673634
rect 132646 673398 132882 673634
rect 132326 637718 132562 637954
rect 132646 637718 132882 637954
rect 132326 637398 132562 637634
rect 132646 637398 132882 637634
rect 132326 601718 132562 601954
rect 132646 601718 132882 601954
rect 132326 601398 132562 601634
rect 132646 601398 132882 601634
rect 132326 565718 132562 565954
rect 132646 565718 132882 565954
rect 132326 565398 132562 565634
rect 132646 565398 132882 565634
rect 132326 529718 132562 529954
rect 132646 529718 132882 529954
rect 132326 529398 132562 529634
rect 132646 529398 132882 529634
rect 132326 493718 132562 493954
rect 132646 493718 132882 493954
rect 132326 493398 132562 493634
rect 132646 493398 132882 493634
rect 132326 457718 132562 457954
rect 132646 457718 132882 457954
rect 132326 457398 132562 457634
rect 132646 457398 132882 457634
rect 132326 421718 132562 421954
rect 132646 421718 132882 421954
rect 132326 421398 132562 421634
rect 132646 421398 132882 421634
rect 132326 385718 132562 385954
rect 132646 385718 132882 385954
rect 132326 385398 132562 385634
rect 132646 385398 132882 385634
rect 132326 349718 132562 349954
rect 132646 349718 132882 349954
rect 132326 349398 132562 349634
rect 132646 349398 132882 349634
rect 132326 313718 132562 313954
rect 132646 313718 132882 313954
rect 132326 313398 132562 313634
rect 132646 313398 132882 313634
rect 132326 277718 132562 277954
rect 132646 277718 132882 277954
rect 132326 277398 132562 277634
rect 132646 277398 132882 277634
rect 136826 710362 137062 710598
rect 137146 710362 137382 710598
rect 136826 710042 137062 710278
rect 137146 710042 137382 710278
rect 136826 678218 137062 678454
rect 137146 678218 137382 678454
rect 136826 677898 137062 678134
rect 137146 677898 137382 678134
rect 136826 642218 137062 642454
rect 137146 642218 137382 642454
rect 136826 641898 137062 642134
rect 137146 641898 137382 642134
rect 136826 606218 137062 606454
rect 137146 606218 137382 606454
rect 136826 605898 137062 606134
rect 137146 605898 137382 606134
rect 136826 570218 137062 570454
rect 137146 570218 137382 570454
rect 136826 569898 137062 570134
rect 137146 569898 137382 570134
rect 136826 534218 137062 534454
rect 137146 534218 137382 534454
rect 136826 533898 137062 534134
rect 137146 533898 137382 534134
rect 136826 498218 137062 498454
rect 137146 498218 137382 498454
rect 136826 497898 137062 498134
rect 137146 497898 137382 498134
rect 136826 462218 137062 462454
rect 137146 462218 137382 462454
rect 136826 461898 137062 462134
rect 137146 461898 137382 462134
rect 136826 426218 137062 426454
rect 137146 426218 137382 426454
rect 136826 425898 137062 426134
rect 137146 425898 137382 426134
rect 136826 390218 137062 390454
rect 137146 390218 137382 390454
rect 136826 389898 137062 390134
rect 137146 389898 137382 390134
rect 136826 354218 137062 354454
rect 137146 354218 137382 354454
rect 136826 353898 137062 354134
rect 137146 353898 137382 354134
rect 136826 318218 137062 318454
rect 137146 318218 137382 318454
rect 136826 317898 137062 318134
rect 137146 317898 137382 318134
rect 136826 282218 137062 282454
rect 137146 282218 137382 282454
rect 136826 281898 137062 282134
rect 137146 281898 137382 282134
rect 136826 246218 137062 246454
rect 137146 246218 137382 246454
rect 136826 245898 137062 246134
rect 137146 245898 137382 246134
rect 141326 711322 141562 711558
rect 141646 711322 141882 711558
rect 141326 711002 141562 711238
rect 141646 711002 141882 711238
rect 141326 682718 141562 682954
rect 141646 682718 141882 682954
rect 141326 682398 141562 682634
rect 141646 682398 141882 682634
rect 141326 646718 141562 646954
rect 141646 646718 141882 646954
rect 141326 646398 141562 646634
rect 141646 646398 141882 646634
rect 141326 610718 141562 610954
rect 141646 610718 141882 610954
rect 141326 610398 141562 610634
rect 141646 610398 141882 610634
rect 141326 574718 141562 574954
rect 141646 574718 141882 574954
rect 141326 574398 141562 574634
rect 141646 574398 141882 574634
rect 141326 538718 141562 538954
rect 141646 538718 141882 538954
rect 141326 538398 141562 538634
rect 141646 538398 141882 538634
rect 141326 502718 141562 502954
rect 141646 502718 141882 502954
rect 141326 502398 141562 502634
rect 141646 502398 141882 502634
rect 141326 466718 141562 466954
rect 141646 466718 141882 466954
rect 141326 466398 141562 466634
rect 141646 466398 141882 466634
rect 141326 430718 141562 430954
rect 141646 430718 141882 430954
rect 141326 430398 141562 430634
rect 141646 430398 141882 430634
rect 141326 394718 141562 394954
rect 141646 394718 141882 394954
rect 141326 394398 141562 394634
rect 141646 394398 141882 394634
rect 141326 358718 141562 358954
rect 141646 358718 141882 358954
rect 141326 358398 141562 358634
rect 141646 358398 141882 358634
rect 141326 322718 141562 322954
rect 141646 322718 141882 322954
rect 141326 322398 141562 322634
rect 141646 322398 141882 322634
rect 141326 286718 141562 286954
rect 141646 286718 141882 286954
rect 141326 286398 141562 286634
rect 141646 286398 141882 286634
rect 141326 250718 141562 250954
rect 141646 250718 141882 250954
rect 141326 250398 141562 250634
rect 141646 250398 141882 250634
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 150326 705562 150562 705798
rect 150646 705562 150882 705798
rect 150326 705242 150562 705478
rect 150646 705242 150882 705478
rect 150326 691718 150562 691954
rect 150646 691718 150882 691954
rect 150326 691398 150562 691634
rect 150646 691398 150882 691634
rect 150326 655718 150562 655954
rect 150646 655718 150882 655954
rect 150326 655398 150562 655634
rect 150646 655398 150882 655634
rect 150326 619718 150562 619954
rect 150646 619718 150882 619954
rect 150326 619398 150562 619634
rect 150646 619398 150882 619634
rect 150326 583718 150562 583954
rect 150646 583718 150882 583954
rect 150326 583398 150562 583634
rect 150646 583398 150882 583634
rect 150326 547718 150562 547954
rect 150646 547718 150882 547954
rect 150326 547398 150562 547634
rect 150646 547398 150882 547634
rect 150326 511718 150562 511954
rect 150646 511718 150882 511954
rect 150326 511398 150562 511634
rect 150646 511398 150882 511634
rect 150326 475718 150562 475954
rect 150646 475718 150882 475954
rect 150326 475398 150562 475634
rect 150646 475398 150882 475634
rect 150326 439718 150562 439954
rect 150646 439718 150882 439954
rect 150326 439398 150562 439634
rect 150646 439398 150882 439634
rect 150326 403718 150562 403954
rect 150646 403718 150882 403954
rect 150326 403398 150562 403634
rect 150646 403398 150882 403634
rect 150326 367718 150562 367954
rect 150646 367718 150882 367954
rect 150326 367398 150562 367634
rect 150646 367398 150882 367634
rect 150326 331718 150562 331954
rect 150646 331718 150882 331954
rect 150326 331398 150562 331634
rect 150646 331398 150882 331634
rect 150326 295718 150562 295954
rect 150646 295718 150882 295954
rect 150326 295398 150562 295634
rect 150646 295398 150882 295634
rect 150326 259718 150562 259954
rect 150646 259718 150882 259954
rect 150326 259398 150562 259634
rect 150646 259398 150882 259634
rect 154826 706522 155062 706758
rect 155146 706522 155382 706758
rect 154826 706202 155062 706438
rect 155146 706202 155382 706438
rect 154826 696218 155062 696454
rect 155146 696218 155382 696454
rect 154826 695898 155062 696134
rect 155146 695898 155382 696134
rect 154826 660218 155062 660454
rect 155146 660218 155382 660454
rect 154826 659898 155062 660134
rect 155146 659898 155382 660134
rect 154826 624218 155062 624454
rect 155146 624218 155382 624454
rect 154826 623898 155062 624134
rect 155146 623898 155382 624134
rect 154826 588218 155062 588454
rect 155146 588218 155382 588454
rect 154826 587898 155062 588134
rect 155146 587898 155382 588134
rect 154826 552218 155062 552454
rect 155146 552218 155382 552454
rect 154826 551898 155062 552134
rect 155146 551898 155382 552134
rect 154826 516218 155062 516454
rect 155146 516218 155382 516454
rect 154826 515898 155062 516134
rect 155146 515898 155382 516134
rect 154826 480218 155062 480454
rect 155146 480218 155382 480454
rect 154826 479898 155062 480134
rect 155146 479898 155382 480134
rect 154826 444218 155062 444454
rect 155146 444218 155382 444454
rect 154826 443898 155062 444134
rect 155146 443898 155382 444134
rect 154826 408218 155062 408454
rect 155146 408218 155382 408454
rect 154826 407898 155062 408134
rect 155146 407898 155382 408134
rect 154826 372218 155062 372454
rect 155146 372218 155382 372454
rect 154826 371898 155062 372134
rect 155146 371898 155382 372134
rect 154826 336218 155062 336454
rect 155146 336218 155382 336454
rect 154826 335898 155062 336134
rect 155146 335898 155382 336134
rect 154826 300218 155062 300454
rect 155146 300218 155382 300454
rect 154826 299898 155062 300134
rect 155146 299898 155382 300134
rect 154826 264218 155062 264454
rect 155146 264218 155382 264454
rect 154826 263898 155062 264134
rect 155146 263898 155382 264134
rect 159326 707482 159562 707718
rect 159646 707482 159882 707718
rect 159326 707162 159562 707398
rect 159646 707162 159882 707398
rect 159326 700718 159562 700954
rect 159646 700718 159882 700954
rect 159326 700398 159562 700634
rect 159646 700398 159882 700634
rect 159326 664718 159562 664954
rect 159646 664718 159882 664954
rect 159326 664398 159562 664634
rect 159646 664398 159882 664634
rect 159326 628718 159562 628954
rect 159646 628718 159882 628954
rect 159326 628398 159562 628634
rect 159646 628398 159882 628634
rect 159326 592718 159562 592954
rect 159646 592718 159882 592954
rect 159326 592398 159562 592634
rect 159646 592398 159882 592634
rect 159326 556718 159562 556954
rect 159646 556718 159882 556954
rect 159326 556398 159562 556634
rect 159646 556398 159882 556634
rect 159326 520718 159562 520954
rect 159646 520718 159882 520954
rect 159326 520398 159562 520634
rect 159646 520398 159882 520634
rect 159326 484718 159562 484954
rect 159646 484718 159882 484954
rect 159326 484398 159562 484634
rect 159646 484398 159882 484634
rect 159326 448718 159562 448954
rect 159646 448718 159882 448954
rect 159326 448398 159562 448634
rect 159646 448398 159882 448634
rect 159326 412718 159562 412954
rect 159646 412718 159882 412954
rect 159326 412398 159562 412634
rect 159646 412398 159882 412634
rect 159326 376718 159562 376954
rect 159646 376718 159882 376954
rect 159326 376398 159562 376634
rect 159646 376398 159882 376634
rect 159326 340718 159562 340954
rect 159646 340718 159882 340954
rect 159326 340398 159562 340634
rect 159646 340398 159882 340634
rect 159326 304718 159562 304954
rect 159646 304718 159882 304954
rect 159326 304398 159562 304634
rect 159646 304398 159882 304634
rect 159326 268718 159562 268954
rect 159646 268718 159882 268954
rect 159326 268398 159562 268634
rect 159646 268398 159882 268634
rect 163826 708442 164062 708678
rect 164146 708442 164382 708678
rect 163826 708122 164062 708358
rect 164146 708122 164382 708358
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 168326 709402 168562 709638
rect 168646 709402 168882 709638
rect 168326 709082 168562 709318
rect 168646 709082 168882 709318
rect 168326 673718 168562 673954
rect 168646 673718 168882 673954
rect 168326 673398 168562 673634
rect 168646 673398 168882 673634
rect 168326 637718 168562 637954
rect 168646 637718 168882 637954
rect 168326 637398 168562 637634
rect 168646 637398 168882 637634
rect 168326 601718 168562 601954
rect 168646 601718 168882 601954
rect 168326 601398 168562 601634
rect 168646 601398 168882 601634
rect 168326 565718 168562 565954
rect 168646 565718 168882 565954
rect 168326 565398 168562 565634
rect 168646 565398 168882 565634
rect 168326 529718 168562 529954
rect 168646 529718 168882 529954
rect 168326 529398 168562 529634
rect 168646 529398 168882 529634
rect 168326 493718 168562 493954
rect 168646 493718 168882 493954
rect 168326 493398 168562 493634
rect 168646 493398 168882 493634
rect 168326 457718 168562 457954
rect 168646 457718 168882 457954
rect 168326 457398 168562 457634
rect 168646 457398 168882 457634
rect 168326 421718 168562 421954
rect 168646 421718 168882 421954
rect 168326 421398 168562 421634
rect 168646 421398 168882 421634
rect 168326 385718 168562 385954
rect 168646 385718 168882 385954
rect 168326 385398 168562 385634
rect 168646 385398 168882 385634
rect 168326 349718 168562 349954
rect 168646 349718 168882 349954
rect 168326 349398 168562 349634
rect 168646 349398 168882 349634
rect 168326 313718 168562 313954
rect 168646 313718 168882 313954
rect 168326 313398 168562 313634
rect 168646 313398 168882 313634
rect 168326 277718 168562 277954
rect 168646 277718 168882 277954
rect 168326 277398 168562 277634
rect 168646 277398 168882 277634
rect 172826 710362 173062 710598
rect 173146 710362 173382 710598
rect 172826 710042 173062 710278
rect 173146 710042 173382 710278
rect 172826 678218 173062 678454
rect 173146 678218 173382 678454
rect 172826 677898 173062 678134
rect 173146 677898 173382 678134
rect 172826 642218 173062 642454
rect 173146 642218 173382 642454
rect 172826 641898 173062 642134
rect 173146 641898 173382 642134
rect 172826 606218 173062 606454
rect 173146 606218 173382 606454
rect 172826 605898 173062 606134
rect 173146 605898 173382 606134
rect 172826 570218 173062 570454
rect 173146 570218 173382 570454
rect 172826 569898 173062 570134
rect 173146 569898 173382 570134
rect 172826 534218 173062 534454
rect 173146 534218 173382 534454
rect 172826 533898 173062 534134
rect 173146 533898 173382 534134
rect 172826 498218 173062 498454
rect 173146 498218 173382 498454
rect 172826 497898 173062 498134
rect 173146 497898 173382 498134
rect 172826 462218 173062 462454
rect 173146 462218 173382 462454
rect 172826 461898 173062 462134
rect 173146 461898 173382 462134
rect 172826 426218 173062 426454
rect 173146 426218 173382 426454
rect 172826 425898 173062 426134
rect 173146 425898 173382 426134
rect 172826 390218 173062 390454
rect 173146 390218 173382 390454
rect 172826 389898 173062 390134
rect 173146 389898 173382 390134
rect 172826 354218 173062 354454
rect 173146 354218 173382 354454
rect 172826 353898 173062 354134
rect 173146 353898 173382 354134
rect 172826 318218 173062 318454
rect 173146 318218 173382 318454
rect 172826 317898 173062 318134
rect 173146 317898 173382 318134
rect 172826 282218 173062 282454
rect 173146 282218 173382 282454
rect 172826 281898 173062 282134
rect 173146 281898 173382 282134
rect 172826 246218 173062 246454
rect 173146 246218 173382 246454
rect 172826 245898 173062 246134
rect 173146 245898 173382 246134
rect 177326 711322 177562 711558
rect 177646 711322 177882 711558
rect 177326 711002 177562 711238
rect 177646 711002 177882 711238
rect 177326 682718 177562 682954
rect 177646 682718 177882 682954
rect 177326 682398 177562 682634
rect 177646 682398 177882 682634
rect 177326 646718 177562 646954
rect 177646 646718 177882 646954
rect 177326 646398 177562 646634
rect 177646 646398 177882 646634
rect 177326 610718 177562 610954
rect 177646 610718 177882 610954
rect 177326 610398 177562 610634
rect 177646 610398 177882 610634
rect 177326 574718 177562 574954
rect 177646 574718 177882 574954
rect 177326 574398 177562 574634
rect 177646 574398 177882 574634
rect 177326 538718 177562 538954
rect 177646 538718 177882 538954
rect 177326 538398 177562 538634
rect 177646 538398 177882 538634
rect 177326 502718 177562 502954
rect 177646 502718 177882 502954
rect 177326 502398 177562 502634
rect 177646 502398 177882 502634
rect 177326 466718 177562 466954
rect 177646 466718 177882 466954
rect 177326 466398 177562 466634
rect 177646 466398 177882 466634
rect 177326 430718 177562 430954
rect 177646 430718 177882 430954
rect 177326 430398 177562 430634
rect 177646 430398 177882 430634
rect 177326 394718 177562 394954
rect 177646 394718 177882 394954
rect 177326 394398 177562 394634
rect 177646 394398 177882 394634
rect 177326 358718 177562 358954
rect 177646 358718 177882 358954
rect 177326 358398 177562 358634
rect 177646 358398 177882 358634
rect 177326 322718 177562 322954
rect 177646 322718 177882 322954
rect 177326 322398 177562 322634
rect 177646 322398 177882 322634
rect 177326 286718 177562 286954
rect 177646 286718 177882 286954
rect 177326 286398 177562 286634
rect 177646 286398 177882 286634
rect 177326 250718 177562 250954
rect 177646 250718 177882 250954
rect 177326 250398 177562 250634
rect 177646 250398 177882 250634
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 186326 705562 186562 705798
rect 186646 705562 186882 705798
rect 186326 705242 186562 705478
rect 186646 705242 186882 705478
rect 186326 691718 186562 691954
rect 186646 691718 186882 691954
rect 186326 691398 186562 691634
rect 186646 691398 186882 691634
rect 186326 655718 186562 655954
rect 186646 655718 186882 655954
rect 186326 655398 186562 655634
rect 186646 655398 186882 655634
rect 186326 619718 186562 619954
rect 186646 619718 186882 619954
rect 186326 619398 186562 619634
rect 186646 619398 186882 619634
rect 186326 583718 186562 583954
rect 186646 583718 186882 583954
rect 186326 583398 186562 583634
rect 186646 583398 186882 583634
rect 186326 547718 186562 547954
rect 186646 547718 186882 547954
rect 186326 547398 186562 547634
rect 186646 547398 186882 547634
rect 186326 511718 186562 511954
rect 186646 511718 186882 511954
rect 186326 511398 186562 511634
rect 186646 511398 186882 511634
rect 186326 475718 186562 475954
rect 186646 475718 186882 475954
rect 186326 475398 186562 475634
rect 186646 475398 186882 475634
rect 186326 439718 186562 439954
rect 186646 439718 186882 439954
rect 186326 439398 186562 439634
rect 186646 439398 186882 439634
rect 186326 403718 186562 403954
rect 186646 403718 186882 403954
rect 186326 403398 186562 403634
rect 186646 403398 186882 403634
rect 186326 367718 186562 367954
rect 186646 367718 186882 367954
rect 186326 367398 186562 367634
rect 186646 367398 186882 367634
rect 186326 331718 186562 331954
rect 186646 331718 186882 331954
rect 186326 331398 186562 331634
rect 186646 331398 186882 331634
rect 186326 295718 186562 295954
rect 186646 295718 186882 295954
rect 186326 295398 186562 295634
rect 186646 295398 186882 295634
rect 186326 259718 186562 259954
rect 186646 259718 186882 259954
rect 186326 259398 186562 259634
rect 186646 259398 186882 259634
rect 190826 706522 191062 706758
rect 191146 706522 191382 706758
rect 190826 706202 191062 706438
rect 191146 706202 191382 706438
rect 190826 696218 191062 696454
rect 191146 696218 191382 696454
rect 190826 695898 191062 696134
rect 191146 695898 191382 696134
rect 190826 660218 191062 660454
rect 191146 660218 191382 660454
rect 190826 659898 191062 660134
rect 191146 659898 191382 660134
rect 190826 624218 191062 624454
rect 191146 624218 191382 624454
rect 190826 623898 191062 624134
rect 191146 623898 191382 624134
rect 190826 588218 191062 588454
rect 191146 588218 191382 588454
rect 190826 587898 191062 588134
rect 191146 587898 191382 588134
rect 190826 552218 191062 552454
rect 191146 552218 191382 552454
rect 190826 551898 191062 552134
rect 191146 551898 191382 552134
rect 190826 516218 191062 516454
rect 191146 516218 191382 516454
rect 190826 515898 191062 516134
rect 191146 515898 191382 516134
rect 190826 480218 191062 480454
rect 191146 480218 191382 480454
rect 190826 479898 191062 480134
rect 191146 479898 191382 480134
rect 190826 444218 191062 444454
rect 191146 444218 191382 444454
rect 190826 443898 191062 444134
rect 191146 443898 191382 444134
rect 190826 408218 191062 408454
rect 191146 408218 191382 408454
rect 190826 407898 191062 408134
rect 191146 407898 191382 408134
rect 190826 372218 191062 372454
rect 191146 372218 191382 372454
rect 190826 371898 191062 372134
rect 191146 371898 191382 372134
rect 190826 336218 191062 336454
rect 191146 336218 191382 336454
rect 190826 335898 191062 336134
rect 191146 335898 191382 336134
rect 190826 300218 191062 300454
rect 191146 300218 191382 300454
rect 190826 299898 191062 300134
rect 191146 299898 191382 300134
rect 190826 264218 191062 264454
rect 191146 264218 191382 264454
rect 190826 263898 191062 264134
rect 191146 263898 191382 264134
rect 195326 707482 195562 707718
rect 195646 707482 195882 707718
rect 195326 707162 195562 707398
rect 195646 707162 195882 707398
rect 195326 700718 195562 700954
rect 195646 700718 195882 700954
rect 195326 700398 195562 700634
rect 195646 700398 195882 700634
rect 195326 664718 195562 664954
rect 195646 664718 195882 664954
rect 195326 664398 195562 664634
rect 195646 664398 195882 664634
rect 195326 628718 195562 628954
rect 195646 628718 195882 628954
rect 195326 628398 195562 628634
rect 195646 628398 195882 628634
rect 195326 592718 195562 592954
rect 195646 592718 195882 592954
rect 195326 592398 195562 592634
rect 195646 592398 195882 592634
rect 195326 556718 195562 556954
rect 195646 556718 195882 556954
rect 195326 556398 195562 556634
rect 195646 556398 195882 556634
rect 195326 520718 195562 520954
rect 195646 520718 195882 520954
rect 195326 520398 195562 520634
rect 195646 520398 195882 520634
rect 195326 484718 195562 484954
rect 195646 484718 195882 484954
rect 195326 484398 195562 484634
rect 195646 484398 195882 484634
rect 195326 448718 195562 448954
rect 195646 448718 195882 448954
rect 195326 448398 195562 448634
rect 195646 448398 195882 448634
rect 195326 412718 195562 412954
rect 195646 412718 195882 412954
rect 195326 412398 195562 412634
rect 195646 412398 195882 412634
rect 195326 376718 195562 376954
rect 195646 376718 195882 376954
rect 195326 376398 195562 376634
rect 195646 376398 195882 376634
rect 195326 340718 195562 340954
rect 195646 340718 195882 340954
rect 195326 340398 195562 340634
rect 195646 340398 195882 340634
rect 195326 304718 195562 304954
rect 195646 304718 195882 304954
rect 195326 304398 195562 304634
rect 195646 304398 195882 304634
rect 195326 268718 195562 268954
rect 195646 268718 195882 268954
rect 195326 268398 195562 268634
rect 195646 268398 195882 268634
rect 199826 708442 200062 708678
rect 200146 708442 200382 708678
rect 199826 708122 200062 708358
rect 200146 708122 200382 708358
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 204326 709402 204562 709638
rect 204646 709402 204882 709638
rect 204326 709082 204562 709318
rect 204646 709082 204882 709318
rect 204326 673718 204562 673954
rect 204646 673718 204882 673954
rect 204326 673398 204562 673634
rect 204646 673398 204882 673634
rect 204326 637718 204562 637954
rect 204646 637718 204882 637954
rect 204326 637398 204562 637634
rect 204646 637398 204882 637634
rect 204326 601718 204562 601954
rect 204646 601718 204882 601954
rect 204326 601398 204562 601634
rect 204646 601398 204882 601634
rect 204326 565718 204562 565954
rect 204646 565718 204882 565954
rect 204326 565398 204562 565634
rect 204646 565398 204882 565634
rect 204326 529718 204562 529954
rect 204646 529718 204882 529954
rect 204326 529398 204562 529634
rect 204646 529398 204882 529634
rect 204326 493718 204562 493954
rect 204646 493718 204882 493954
rect 204326 493398 204562 493634
rect 204646 493398 204882 493634
rect 204326 457718 204562 457954
rect 204646 457718 204882 457954
rect 204326 457398 204562 457634
rect 204646 457398 204882 457634
rect 204326 421718 204562 421954
rect 204646 421718 204882 421954
rect 204326 421398 204562 421634
rect 204646 421398 204882 421634
rect 204326 385718 204562 385954
rect 204646 385718 204882 385954
rect 204326 385398 204562 385634
rect 204646 385398 204882 385634
rect 204326 349718 204562 349954
rect 204646 349718 204882 349954
rect 204326 349398 204562 349634
rect 204646 349398 204882 349634
rect 204326 313718 204562 313954
rect 204646 313718 204882 313954
rect 204326 313398 204562 313634
rect 204646 313398 204882 313634
rect 204326 277718 204562 277954
rect 204646 277718 204882 277954
rect 204326 277398 204562 277634
rect 204646 277398 204882 277634
rect 208826 710362 209062 710598
rect 209146 710362 209382 710598
rect 208826 710042 209062 710278
rect 209146 710042 209382 710278
rect 208826 678218 209062 678454
rect 209146 678218 209382 678454
rect 208826 677898 209062 678134
rect 209146 677898 209382 678134
rect 208826 642218 209062 642454
rect 209146 642218 209382 642454
rect 208826 641898 209062 642134
rect 209146 641898 209382 642134
rect 208826 606218 209062 606454
rect 209146 606218 209382 606454
rect 208826 605898 209062 606134
rect 209146 605898 209382 606134
rect 208826 570218 209062 570454
rect 209146 570218 209382 570454
rect 208826 569898 209062 570134
rect 209146 569898 209382 570134
rect 208826 534218 209062 534454
rect 209146 534218 209382 534454
rect 208826 533898 209062 534134
rect 209146 533898 209382 534134
rect 208826 498218 209062 498454
rect 209146 498218 209382 498454
rect 208826 497898 209062 498134
rect 209146 497898 209382 498134
rect 208826 462218 209062 462454
rect 209146 462218 209382 462454
rect 208826 461898 209062 462134
rect 209146 461898 209382 462134
rect 208826 426218 209062 426454
rect 209146 426218 209382 426454
rect 208826 425898 209062 426134
rect 209146 425898 209382 426134
rect 208826 390218 209062 390454
rect 209146 390218 209382 390454
rect 208826 389898 209062 390134
rect 209146 389898 209382 390134
rect 208826 354218 209062 354454
rect 209146 354218 209382 354454
rect 208826 353898 209062 354134
rect 209146 353898 209382 354134
rect 208826 318218 209062 318454
rect 209146 318218 209382 318454
rect 208826 317898 209062 318134
rect 209146 317898 209382 318134
rect 208826 282218 209062 282454
rect 209146 282218 209382 282454
rect 208826 281898 209062 282134
rect 209146 281898 209382 282134
rect 208826 246218 209062 246454
rect 209146 246218 209382 246454
rect 208826 245898 209062 246134
rect 209146 245898 209382 246134
rect 213326 711322 213562 711558
rect 213646 711322 213882 711558
rect 213326 711002 213562 711238
rect 213646 711002 213882 711238
rect 213326 682718 213562 682954
rect 213646 682718 213882 682954
rect 213326 682398 213562 682634
rect 213646 682398 213882 682634
rect 213326 646718 213562 646954
rect 213646 646718 213882 646954
rect 213326 646398 213562 646634
rect 213646 646398 213882 646634
rect 213326 610718 213562 610954
rect 213646 610718 213882 610954
rect 213326 610398 213562 610634
rect 213646 610398 213882 610634
rect 213326 574718 213562 574954
rect 213646 574718 213882 574954
rect 213326 574398 213562 574634
rect 213646 574398 213882 574634
rect 213326 538718 213562 538954
rect 213646 538718 213882 538954
rect 213326 538398 213562 538634
rect 213646 538398 213882 538634
rect 213326 502718 213562 502954
rect 213646 502718 213882 502954
rect 213326 502398 213562 502634
rect 213646 502398 213882 502634
rect 213326 466718 213562 466954
rect 213646 466718 213882 466954
rect 213326 466398 213562 466634
rect 213646 466398 213882 466634
rect 213326 430718 213562 430954
rect 213646 430718 213882 430954
rect 213326 430398 213562 430634
rect 213646 430398 213882 430634
rect 213326 394718 213562 394954
rect 213646 394718 213882 394954
rect 213326 394398 213562 394634
rect 213646 394398 213882 394634
rect 213326 358718 213562 358954
rect 213646 358718 213882 358954
rect 213326 358398 213562 358634
rect 213646 358398 213882 358634
rect 213326 322718 213562 322954
rect 213646 322718 213882 322954
rect 213326 322398 213562 322634
rect 213646 322398 213882 322634
rect 213326 286718 213562 286954
rect 213646 286718 213882 286954
rect 213326 286398 213562 286634
rect 213646 286398 213882 286634
rect 213326 250718 213562 250954
rect 213646 250718 213882 250954
rect 213326 250398 213562 250634
rect 213646 250398 213882 250634
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 222326 705562 222562 705798
rect 222646 705562 222882 705798
rect 222326 705242 222562 705478
rect 222646 705242 222882 705478
rect 222326 691718 222562 691954
rect 222646 691718 222882 691954
rect 222326 691398 222562 691634
rect 222646 691398 222882 691634
rect 222326 655718 222562 655954
rect 222646 655718 222882 655954
rect 222326 655398 222562 655634
rect 222646 655398 222882 655634
rect 222326 619718 222562 619954
rect 222646 619718 222882 619954
rect 222326 619398 222562 619634
rect 222646 619398 222882 619634
rect 222326 583718 222562 583954
rect 222646 583718 222882 583954
rect 222326 583398 222562 583634
rect 222646 583398 222882 583634
rect 222326 547718 222562 547954
rect 222646 547718 222882 547954
rect 222326 547398 222562 547634
rect 222646 547398 222882 547634
rect 222326 511718 222562 511954
rect 222646 511718 222882 511954
rect 222326 511398 222562 511634
rect 222646 511398 222882 511634
rect 222326 475718 222562 475954
rect 222646 475718 222882 475954
rect 222326 475398 222562 475634
rect 222646 475398 222882 475634
rect 222326 439718 222562 439954
rect 222646 439718 222882 439954
rect 222326 439398 222562 439634
rect 222646 439398 222882 439634
rect 222326 403718 222562 403954
rect 222646 403718 222882 403954
rect 222326 403398 222562 403634
rect 222646 403398 222882 403634
rect 222326 367718 222562 367954
rect 222646 367718 222882 367954
rect 222326 367398 222562 367634
rect 222646 367398 222882 367634
rect 222326 331718 222562 331954
rect 222646 331718 222882 331954
rect 222326 331398 222562 331634
rect 222646 331398 222882 331634
rect 222326 295718 222562 295954
rect 222646 295718 222882 295954
rect 222326 295398 222562 295634
rect 222646 295398 222882 295634
rect 222326 259718 222562 259954
rect 222646 259718 222882 259954
rect 222326 259398 222562 259634
rect 222646 259398 222882 259634
rect 226826 706522 227062 706758
rect 227146 706522 227382 706758
rect 226826 706202 227062 706438
rect 227146 706202 227382 706438
rect 226826 696218 227062 696454
rect 227146 696218 227382 696454
rect 226826 695898 227062 696134
rect 227146 695898 227382 696134
rect 226826 660218 227062 660454
rect 227146 660218 227382 660454
rect 226826 659898 227062 660134
rect 227146 659898 227382 660134
rect 226826 624218 227062 624454
rect 227146 624218 227382 624454
rect 226826 623898 227062 624134
rect 227146 623898 227382 624134
rect 226826 588218 227062 588454
rect 227146 588218 227382 588454
rect 226826 587898 227062 588134
rect 227146 587898 227382 588134
rect 226826 552218 227062 552454
rect 227146 552218 227382 552454
rect 226826 551898 227062 552134
rect 227146 551898 227382 552134
rect 226826 516218 227062 516454
rect 227146 516218 227382 516454
rect 226826 515898 227062 516134
rect 227146 515898 227382 516134
rect 226826 480218 227062 480454
rect 227146 480218 227382 480454
rect 226826 479898 227062 480134
rect 227146 479898 227382 480134
rect 226826 444218 227062 444454
rect 227146 444218 227382 444454
rect 226826 443898 227062 444134
rect 227146 443898 227382 444134
rect 226826 408218 227062 408454
rect 227146 408218 227382 408454
rect 226826 407898 227062 408134
rect 227146 407898 227382 408134
rect 226826 372218 227062 372454
rect 227146 372218 227382 372454
rect 226826 371898 227062 372134
rect 227146 371898 227382 372134
rect 226826 336218 227062 336454
rect 227146 336218 227382 336454
rect 226826 335898 227062 336134
rect 227146 335898 227382 336134
rect 226826 300218 227062 300454
rect 227146 300218 227382 300454
rect 226826 299898 227062 300134
rect 227146 299898 227382 300134
rect 226826 264218 227062 264454
rect 227146 264218 227382 264454
rect 226826 263898 227062 264134
rect 227146 263898 227382 264134
rect 231326 707482 231562 707718
rect 231646 707482 231882 707718
rect 231326 707162 231562 707398
rect 231646 707162 231882 707398
rect 231326 700718 231562 700954
rect 231646 700718 231882 700954
rect 231326 700398 231562 700634
rect 231646 700398 231882 700634
rect 231326 664718 231562 664954
rect 231646 664718 231882 664954
rect 231326 664398 231562 664634
rect 231646 664398 231882 664634
rect 231326 628718 231562 628954
rect 231646 628718 231882 628954
rect 231326 628398 231562 628634
rect 231646 628398 231882 628634
rect 231326 592718 231562 592954
rect 231646 592718 231882 592954
rect 231326 592398 231562 592634
rect 231646 592398 231882 592634
rect 231326 556718 231562 556954
rect 231646 556718 231882 556954
rect 231326 556398 231562 556634
rect 231646 556398 231882 556634
rect 231326 520718 231562 520954
rect 231646 520718 231882 520954
rect 231326 520398 231562 520634
rect 231646 520398 231882 520634
rect 231326 484718 231562 484954
rect 231646 484718 231882 484954
rect 231326 484398 231562 484634
rect 231646 484398 231882 484634
rect 231326 448718 231562 448954
rect 231646 448718 231882 448954
rect 231326 448398 231562 448634
rect 231646 448398 231882 448634
rect 231326 412718 231562 412954
rect 231646 412718 231882 412954
rect 231326 412398 231562 412634
rect 231646 412398 231882 412634
rect 231326 376718 231562 376954
rect 231646 376718 231882 376954
rect 231326 376398 231562 376634
rect 231646 376398 231882 376634
rect 231326 340718 231562 340954
rect 231646 340718 231882 340954
rect 231326 340398 231562 340634
rect 231646 340398 231882 340634
rect 231326 304718 231562 304954
rect 231646 304718 231882 304954
rect 231326 304398 231562 304634
rect 231646 304398 231882 304634
rect 231326 268718 231562 268954
rect 231646 268718 231882 268954
rect 231326 268398 231562 268634
rect 231646 268398 231882 268634
rect 235826 708442 236062 708678
rect 236146 708442 236382 708678
rect 235826 708122 236062 708358
rect 236146 708122 236382 708358
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 235826 273218 236062 273454
rect 236146 273218 236382 273454
rect 235826 272898 236062 273134
rect 236146 272898 236382 273134
rect 240326 709402 240562 709638
rect 240646 709402 240882 709638
rect 240326 709082 240562 709318
rect 240646 709082 240882 709318
rect 240326 673718 240562 673954
rect 240646 673718 240882 673954
rect 240326 673398 240562 673634
rect 240646 673398 240882 673634
rect 240326 637718 240562 637954
rect 240646 637718 240882 637954
rect 240326 637398 240562 637634
rect 240646 637398 240882 637634
rect 240326 601718 240562 601954
rect 240646 601718 240882 601954
rect 240326 601398 240562 601634
rect 240646 601398 240882 601634
rect 240326 565718 240562 565954
rect 240646 565718 240882 565954
rect 240326 565398 240562 565634
rect 240646 565398 240882 565634
rect 240326 529718 240562 529954
rect 240646 529718 240882 529954
rect 240326 529398 240562 529634
rect 240646 529398 240882 529634
rect 240326 493718 240562 493954
rect 240646 493718 240882 493954
rect 240326 493398 240562 493634
rect 240646 493398 240882 493634
rect 240326 457718 240562 457954
rect 240646 457718 240882 457954
rect 240326 457398 240562 457634
rect 240646 457398 240882 457634
rect 240326 421718 240562 421954
rect 240646 421718 240882 421954
rect 240326 421398 240562 421634
rect 240646 421398 240882 421634
rect 240326 385718 240562 385954
rect 240646 385718 240882 385954
rect 240326 385398 240562 385634
rect 240646 385398 240882 385634
rect 240326 349718 240562 349954
rect 240646 349718 240882 349954
rect 240326 349398 240562 349634
rect 240646 349398 240882 349634
rect 240326 313718 240562 313954
rect 240646 313718 240882 313954
rect 240326 313398 240562 313634
rect 240646 313398 240882 313634
rect 240326 277718 240562 277954
rect 240646 277718 240882 277954
rect 240326 277398 240562 277634
rect 240646 277398 240882 277634
rect 244826 710362 245062 710598
rect 245146 710362 245382 710598
rect 244826 710042 245062 710278
rect 245146 710042 245382 710278
rect 244826 678218 245062 678454
rect 245146 678218 245382 678454
rect 244826 677898 245062 678134
rect 245146 677898 245382 678134
rect 244826 642218 245062 642454
rect 245146 642218 245382 642454
rect 244826 641898 245062 642134
rect 245146 641898 245382 642134
rect 244826 606218 245062 606454
rect 245146 606218 245382 606454
rect 244826 605898 245062 606134
rect 245146 605898 245382 606134
rect 244826 570218 245062 570454
rect 245146 570218 245382 570454
rect 244826 569898 245062 570134
rect 245146 569898 245382 570134
rect 244826 534218 245062 534454
rect 245146 534218 245382 534454
rect 244826 533898 245062 534134
rect 245146 533898 245382 534134
rect 244826 498218 245062 498454
rect 245146 498218 245382 498454
rect 244826 497898 245062 498134
rect 245146 497898 245382 498134
rect 244826 462218 245062 462454
rect 245146 462218 245382 462454
rect 244826 461898 245062 462134
rect 245146 461898 245382 462134
rect 244826 426218 245062 426454
rect 245146 426218 245382 426454
rect 244826 425898 245062 426134
rect 245146 425898 245382 426134
rect 244826 390218 245062 390454
rect 245146 390218 245382 390454
rect 244826 389898 245062 390134
rect 245146 389898 245382 390134
rect 244826 354218 245062 354454
rect 245146 354218 245382 354454
rect 244826 353898 245062 354134
rect 245146 353898 245382 354134
rect 244826 318218 245062 318454
rect 245146 318218 245382 318454
rect 244826 317898 245062 318134
rect 245146 317898 245382 318134
rect 244826 282218 245062 282454
rect 245146 282218 245382 282454
rect 244826 281898 245062 282134
rect 245146 281898 245382 282134
rect 244826 246218 245062 246454
rect 245146 246218 245382 246454
rect 244826 245898 245062 246134
rect 245146 245898 245382 246134
rect 249326 711322 249562 711558
rect 249646 711322 249882 711558
rect 249326 711002 249562 711238
rect 249646 711002 249882 711238
rect 249326 682718 249562 682954
rect 249646 682718 249882 682954
rect 249326 682398 249562 682634
rect 249646 682398 249882 682634
rect 249326 646718 249562 646954
rect 249646 646718 249882 646954
rect 249326 646398 249562 646634
rect 249646 646398 249882 646634
rect 249326 610718 249562 610954
rect 249646 610718 249882 610954
rect 249326 610398 249562 610634
rect 249646 610398 249882 610634
rect 249326 574718 249562 574954
rect 249646 574718 249882 574954
rect 249326 574398 249562 574634
rect 249646 574398 249882 574634
rect 249326 538718 249562 538954
rect 249646 538718 249882 538954
rect 249326 538398 249562 538634
rect 249646 538398 249882 538634
rect 249326 502718 249562 502954
rect 249646 502718 249882 502954
rect 249326 502398 249562 502634
rect 249646 502398 249882 502634
rect 249326 466718 249562 466954
rect 249646 466718 249882 466954
rect 249326 466398 249562 466634
rect 249646 466398 249882 466634
rect 249326 430718 249562 430954
rect 249646 430718 249882 430954
rect 249326 430398 249562 430634
rect 249646 430398 249882 430634
rect 249326 394718 249562 394954
rect 249646 394718 249882 394954
rect 249326 394398 249562 394634
rect 249646 394398 249882 394634
rect 249326 358718 249562 358954
rect 249646 358718 249882 358954
rect 249326 358398 249562 358634
rect 249646 358398 249882 358634
rect 249326 322718 249562 322954
rect 249646 322718 249882 322954
rect 249326 322398 249562 322634
rect 249646 322398 249882 322634
rect 249326 286718 249562 286954
rect 249646 286718 249882 286954
rect 249326 286398 249562 286634
rect 249646 286398 249882 286634
rect 249326 250718 249562 250954
rect 249646 250718 249882 250954
rect 249326 250398 249562 250634
rect 249646 250398 249882 250634
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 258326 705562 258562 705798
rect 258646 705562 258882 705798
rect 258326 705242 258562 705478
rect 258646 705242 258882 705478
rect 258326 691718 258562 691954
rect 258646 691718 258882 691954
rect 258326 691398 258562 691634
rect 258646 691398 258882 691634
rect 258326 655718 258562 655954
rect 258646 655718 258882 655954
rect 258326 655398 258562 655634
rect 258646 655398 258882 655634
rect 258326 619718 258562 619954
rect 258646 619718 258882 619954
rect 258326 619398 258562 619634
rect 258646 619398 258882 619634
rect 258326 583718 258562 583954
rect 258646 583718 258882 583954
rect 258326 583398 258562 583634
rect 258646 583398 258882 583634
rect 258326 547718 258562 547954
rect 258646 547718 258882 547954
rect 258326 547398 258562 547634
rect 258646 547398 258882 547634
rect 258326 511718 258562 511954
rect 258646 511718 258882 511954
rect 258326 511398 258562 511634
rect 258646 511398 258882 511634
rect 258326 475718 258562 475954
rect 258646 475718 258882 475954
rect 258326 475398 258562 475634
rect 258646 475398 258882 475634
rect 258326 439718 258562 439954
rect 258646 439718 258882 439954
rect 258326 439398 258562 439634
rect 258646 439398 258882 439634
rect 258326 403718 258562 403954
rect 258646 403718 258882 403954
rect 258326 403398 258562 403634
rect 258646 403398 258882 403634
rect 258326 367718 258562 367954
rect 258646 367718 258882 367954
rect 258326 367398 258562 367634
rect 258646 367398 258882 367634
rect 258326 331718 258562 331954
rect 258646 331718 258882 331954
rect 258326 331398 258562 331634
rect 258646 331398 258882 331634
rect 258326 295718 258562 295954
rect 258646 295718 258882 295954
rect 258326 295398 258562 295634
rect 258646 295398 258882 295634
rect 258326 259718 258562 259954
rect 258646 259718 258882 259954
rect 258326 259398 258562 259634
rect 258646 259398 258882 259634
rect 262826 706522 263062 706758
rect 263146 706522 263382 706758
rect 262826 706202 263062 706438
rect 263146 706202 263382 706438
rect 262826 696218 263062 696454
rect 263146 696218 263382 696454
rect 262826 695898 263062 696134
rect 263146 695898 263382 696134
rect 262826 660218 263062 660454
rect 263146 660218 263382 660454
rect 262826 659898 263062 660134
rect 263146 659898 263382 660134
rect 262826 624218 263062 624454
rect 263146 624218 263382 624454
rect 262826 623898 263062 624134
rect 263146 623898 263382 624134
rect 262826 588218 263062 588454
rect 263146 588218 263382 588454
rect 262826 587898 263062 588134
rect 263146 587898 263382 588134
rect 262826 552218 263062 552454
rect 263146 552218 263382 552454
rect 262826 551898 263062 552134
rect 263146 551898 263382 552134
rect 262826 516218 263062 516454
rect 263146 516218 263382 516454
rect 262826 515898 263062 516134
rect 263146 515898 263382 516134
rect 262826 480218 263062 480454
rect 263146 480218 263382 480454
rect 262826 479898 263062 480134
rect 263146 479898 263382 480134
rect 262826 444218 263062 444454
rect 263146 444218 263382 444454
rect 262826 443898 263062 444134
rect 263146 443898 263382 444134
rect 262826 408218 263062 408454
rect 263146 408218 263382 408454
rect 262826 407898 263062 408134
rect 263146 407898 263382 408134
rect 262826 372218 263062 372454
rect 263146 372218 263382 372454
rect 262826 371898 263062 372134
rect 263146 371898 263382 372134
rect 262826 336218 263062 336454
rect 263146 336218 263382 336454
rect 262826 335898 263062 336134
rect 263146 335898 263382 336134
rect 262826 300218 263062 300454
rect 263146 300218 263382 300454
rect 262826 299898 263062 300134
rect 263146 299898 263382 300134
rect 262826 264218 263062 264454
rect 263146 264218 263382 264454
rect 262826 263898 263062 264134
rect 263146 263898 263382 264134
rect 267326 707482 267562 707718
rect 267646 707482 267882 707718
rect 267326 707162 267562 707398
rect 267646 707162 267882 707398
rect 267326 700718 267562 700954
rect 267646 700718 267882 700954
rect 267326 700398 267562 700634
rect 267646 700398 267882 700634
rect 267326 664718 267562 664954
rect 267646 664718 267882 664954
rect 267326 664398 267562 664634
rect 267646 664398 267882 664634
rect 267326 628718 267562 628954
rect 267646 628718 267882 628954
rect 267326 628398 267562 628634
rect 267646 628398 267882 628634
rect 267326 592718 267562 592954
rect 267646 592718 267882 592954
rect 267326 592398 267562 592634
rect 267646 592398 267882 592634
rect 267326 556718 267562 556954
rect 267646 556718 267882 556954
rect 267326 556398 267562 556634
rect 267646 556398 267882 556634
rect 267326 520718 267562 520954
rect 267646 520718 267882 520954
rect 267326 520398 267562 520634
rect 267646 520398 267882 520634
rect 267326 484718 267562 484954
rect 267646 484718 267882 484954
rect 267326 484398 267562 484634
rect 267646 484398 267882 484634
rect 267326 448718 267562 448954
rect 267646 448718 267882 448954
rect 267326 448398 267562 448634
rect 267646 448398 267882 448634
rect 267326 412718 267562 412954
rect 267646 412718 267882 412954
rect 267326 412398 267562 412634
rect 267646 412398 267882 412634
rect 267326 376718 267562 376954
rect 267646 376718 267882 376954
rect 267326 376398 267562 376634
rect 267646 376398 267882 376634
rect 267326 340718 267562 340954
rect 267646 340718 267882 340954
rect 267326 340398 267562 340634
rect 267646 340398 267882 340634
rect 267326 304718 267562 304954
rect 267646 304718 267882 304954
rect 267326 304398 267562 304634
rect 267646 304398 267882 304634
rect 267326 268718 267562 268954
rect 267646 268718 267882 268954
rect 267326 268398 267562 268634
rect 267646 268398 267882 268634
rect 271826 708442 272062 708678
rect 272146 708442 272382 708678
rect 271826 708122 272062 708358
rect 272146 708122 272382 708358
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 276326 709402 276562 709638
rect 276646 709402 276882 709638
rect 276326 709082 276562 709318
rect 276646 709082 276882 709318
rect 276326 673718 276562 673954
rect 276646 673718 276882 673954
rect 276326 673398 276562 673634
rect 276646 673398 276882 673634
rect 276326 637718 276562 637954
rect 276646 637718 276882 637954
rect 276326 637398 276562 637634
rect 276646 637398 276882 637634
rect 276326 601718 276562 601954
rect 276646 601718 276882 601954
rect 276326 601398 276562 601634
rect 276646 601398 276882 601634
rect 276326 565718 276562 565954
rect 276646 565718 276882 565954
rect 276326 565398 276562 565634
rect 276646 565398 276882 565634
rect 276326 529718 276562 529954
rect 276646 529718 276882 529954
rect 276326 529398 276562 529634
rect 276646 529398 276882 529634
rect 276326 493718 276562 493954
rect 276646 493718 276882 493954
rect 276326 493398 276562 493634
rect 276646 493398 276882 493634
rect 276326 457718 276562 457954
rect 276646 457718 276882 457954
rect 276326 457398 276562 457634
rect 276646 457398 276882 457634
rect 276326 421718 276562 421954
rect 276646 421718 276882 421954
rect 276326 421398 276562 421634
rect 276646 421398 276882 421634
rect 276326 385718 276562 385954
rect 276646 385718 276882 385954
rect 276326 385398 276562 385634
rect 276646 385398 276882 385634
rect 276326 349718 276562 349954
rect 276646 349718 276882 349954
rect 276326 349398 276562 349634
rect 276646 349398 276882 349634
rect 276326 313718 276562 313954
rect 276646 313718 276882 313954
rect 276326 313398 276562 313634
rect 276646 313398 276882 313634
rect 276326 277718 276562 277954
rect 276646 277718 276882 277954
rect 276326 277398 276562 277634
rect 276646 277398 276882 277634
rect 280826 710362 281062 710598
rect 281146 710362 281382 710598
rect 280826 710042 281062 710278
rect 281146 710042 281382 710278
rect 280826 678218 281062 678454
rect 281146 678218 281382 678454
rect 280826 677898 281062 678134
rect 281146 677898 281382 678134
rect 280826 642218 281062 642454
rect 281146 642218 281382 642454
rect 280826 641898 281062 642134
rect 281146 641898 281382 642134
rect 280826 606218 281062 606454
rect 281146 606218 281382 606454
rect 280826 605898 281062 606134
rect 281146 605898 281382 606134
rect 280826 570218 281062 570454
rect 281146 570218 281382 570454
rect 280826 569898 281062 570134
rect 281146 569898 281382 570134
rect 280826 534218 281062 534454
rect 281146 534218 281382 534454
rect 280826 533898 281062 534134
rect 281146 533898 281382 534134
rect 280826 498218 281062 498454
rect 281146 498218 281382 498454
rect 280826 497898 281062 498134
rect 281146 497898 281382 498134
rect 280826 462218 281062 462454
rect 281146 462218 281382 462454
rect 280826 461898 281062 462134
rect 281146 461898 281382 462134
rect 280826 426218 281062 426454
rect 281146 426218 281382 426454
rect 280826 425898 281062 426134
rect 281146 425898 281382 426134
rect 280826 390218 281062 390454
rect 281146 390218 281382 390454
rect 280826 389898 281062 390134
rect 281146 389898 281382 390134
rect 280826 354218 281062 354454
rect 281146 354218 281382 354454
rect 280826 353898 281062 354134
rect 281146 353898 281382 354134
rect 280826 318218 281062 318454
rect 281146 318218 281382 318454
rect 280826 317898 281062 318134
rect 281146 317898 281382 318134
rect 280826 282218 281062 282454
rect 281146 282218 281382 282454
rect 280826 281898 281062 282134
rect 281146 281898 281382 282134
rect 280826 246218 281062 246454
rect 281146 246218 281382 246454
rect 280826 245898 281062 246134
rect 281146 245898 281382 246134
rect 285326 711322 285562 711558
rect 285646 711322 285882 711558
rect 285326 711002 285562 711238
rect 285646 711002 285882 711238
rect 285326 682718 285562 682954
rect 285646 682718 285882 682954
rect 285326 682398 285562 682634
rect 285646 682398 285882 682634
rect 285326 646718 285562 646954
rect 285646 646718 285882 646954
rect 285326 646398 285562 646634
rect 285646 646398 285882 646634
rect 285326 610718 285562 610954
rect 285646 610718 285882 610954
rect 285326 610398 285562 610634
rect 285646 610398 285882 610634
rect 285326 574718 285562 574954
rect 285646 574718 285882 574954
rect 285326 574398 285562 574634
rect 285646 574398 285882 574634
rect 285326 538718 285562 538954
rect 285646 538718 285882 538954
rect 285326 538398 285562 538634
rect 285646 538398 285882 538634
rect 285326 502718 285562 502954
rect 285646 502718 285882 502954
rect 285326 502398 285562 502634
rect 285646 502398 285882 502634
rect 285326 466718 285562 466954
rect 285646 466718 285882 466954
rect 285326 466398 285562 466634
rect 285646 466398 285882 466634
rect 285326 430718 285562 430954
rect 285646 430718 285882 430954
rect 285326 430398 285562 430634
rect 285646 430398 285882 430634
rect 285326 394718 285562 394954
rect 285646 394718 285882 394954
rect 285326 394398 285562 394634
rect 285646 394398 285882 394634
rect 285326 358718 285562 358954
rect 285646 358718 285882 358954
rect 285326 358398 285562 358634
rect 285646 358398 285882 358634
rect 285326 322718 285562 322954
rect 285646 322718 285882 322954
rect 285326 322398 285562 322634
rect 285646 322398 285882 322634
rect 285326 286718 285562 286954
rect 285646 286718 285882 286954
rect 285326 286398 285562 286634
rect 285646 286398 285882 286634
rect 285326 250718 285562 250954
rect 285646 250718 285882 250954
rect 285326 250398 285562 250634
rect 285646 250398 285882 250634
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 294326 705562 294562 705798
rect 294646 705562 294882 705798
rect 294326 705242 294562 705478
rect 294646 705242 294882 705478
rect 294326 691718 294562 691954
rect 294646 691718 294882 691954
rect 294326 691398 294562 691634
rect 294646 691398 294882 691634
rect 294326 655718 294562 655954
rect 294646 655718 294882 655954
rect 294326 655398 294562 655634
rect 294646 655398 294882 655634
rect 294326 619718 294562 619954
rect 294646 619718 294882 619954
rect 294326 619398 294562 619634
rect 294646 619398 294882 619634
rect 294326 583718 294562 583954
rect 294646 583718 294882 583954
rect 294326 583398 294562 583634
rect 294646 583398 294882 583634
rect 294326 547718 294562 547954
rect 294646 547718 294882 547954
rect 294326 547398 294562 547634
rect 294646 547398 294882 547634
rect 294326 511718 294562 511954
rect 294646 511718 294882 511954
rect 294326 511398 294562 511634
rect 294646 511398 294882 511634
rect 294326 475718 294562 475954
rect 294646 475718 294882 475954
rect 294326 475398 294562 475634
rect 294646 475398 294882 475634
rect 294326 439718 294562 439954
rect 294646 439718 294882 439954
rect 294326 439398 294562 439634
rect 294646 439398 294882 439634
rect 294326 403718 294562 403954
rect 294646 403718 294882 403954
rect 294326 403398 294562 403634
rect 294646 403398 294882 403634
rect 294326 367718 294562 367954
rect 294646 367718 294882 367954
rect 294326 367398 294562 367634
rect 294646 367398 294882 367634
rect 294326 331718 294562 331954
rect 294646 331718 294882 331954
rect 294326 331398 294562 331634
rect 294646 331398 294882 331634
rect 294326 295718 294562 295954
rect 294646 295718 294882 295954
rect 294326 295398 294562 295634
rect 294646 295398 294882 295634
rect 294326 259718 294562 259954
rect 294646 259718 294882 259954
rect 294326 259398 294562 259634
rect 294646 259398 294882 259634
rect 298826 706522 299062 706758
rect 299146 706522 299382 706758
rect 298826 706202 299062 706438
rect 299146 706202 299382 706438
rect 298826 696218 299062 696454
rect 299146 696218 299382 696454
rect 298826 695898 299062 696134
rect 299146 695898 299382 696134
rect 298826 660218 299062 660454
rect 299146 660218 299382 660454
rect 298826 659898 299062 660134
rect 299146 659898 299382 660134
rect 298826 624218 299062 624454
rect 299146 624218 299382 624454
rect 298826 623898 299062 624134
rect 299146 623898 299382 624134
rect 298826 588218 299062 588454
rect 299146 588218 299382 588454
rect 298826 587898 299062 588134
rect 299146 587898 299382 588134
rect 298826 552218 299062 552454
rect 299146 552218 299382 552454
rect 298826 551898 299062 552134
rect 299146 551898 299382 552134
rect 298826 516218 299062 516454
rect 299146 516218 299382 516454
rect 298826 515898 299062 516134
rect 299146 515898 299382 516134
rect 298826 480218 299062 480454
rect 299146 480218 299382 480454
rect 298826 479898 299062 480134
rect 299146 479898 299382 480134
rect 298826 444218 299062 444454
rect 299146 444218 299382 444454
rect 298826 443898 299062 444134
rect 299146 443898 299382 444134
rect 298826 408218 299062 408454
rect 299146 408218 299382 408454
rect 298826 407898 299062 408134
rect 299146 407898 299382 408134
rect 298826 372218 299062 372454
rect 299146 372218 299382 372454
rect 298826 371898 299062 372134
rect 299146 371898 299382 372134
rect 298826 336218 299062 336454
rect 299146 336218 299382 336454
rect 298826 335898 299062 336134
rect 299146 335898 299382 336134
rect 298826 300218 299062 300454
rect 299146 300218 299382 300454
rect 298826 299898 299062 300134
rect 299146 299898 299382 300134
rect 298826 264218 299062 264454
rect 299146 264218 299382 264454
rect 298826 263898 299062 264134
rect 299146 263898 299382 264134
rect 303326 707482 303562 707718
rect 303646 707482 303882 707718
rect 303326 707162 303562 707398
rect 303646 707162 303882 707398
rect 303326 700718 303562 700954
rect 303646 700718 303882 700954
rect 303326 700398 303562 700634
rect 303646 700398 303882 700634
rect 303326 664718 303562 664954
rect 303646 664718 303882 664954
rect 303326 664398 303562 664634
rect 303646 664398 303882 664634
rect 303326 628718 303562 628954
rect 303646 628718 303882 628954
rect 303326 628398 303562 628634
rect 303646 628398 303882 628634
rect 303326 592718 303562 592954
rect 303646 592718 303882 592954
rect 303326 592398 303562 592634
rect 303646 592398 303882 592634
rect 303326 556718 303562 556954
rect 303646 556718 303882 556954
rect 303326 556398 303562 556634
rect 303646 556398 303882 556634
rect 303326 520718 303562 520954
rect 303646 520718 303882 520954
rect 303326 520398 303562 520634
rect 303646 520398 303882 520634
rect 303326 484718 303562 484954
rect 303646 484718 303882 484954
rect 303326 484398 303562 484634
rect 303646 484398 303882 484634
rect 303326 448718 303562 448954
rect 303646 448718 303882 448954
rect 303326 448398 303562 448634
rect 303646 448398 303882 448634
rect 303326 412718 303562 412954
rect 303646 412718 303882 412954
rect 303326 412398 303562 412634
rect 303646 412398 303882 412634
rect 303326 376718 303562 376954
rect 303646 376718 303882 376954
rect 303326 376398 303562 376634
rect 303646 376398 303882 376634
rect 303326 340718 303562 340954
rect 303646 340718 303882 340954
rect 303326 340398 303562 340634
rect 303646 340398 303882 340634
rect 303326 304718 303562 304954
rect 303646 304718 303882 304954
rect 303326 304398 303562 304634
rect 303646 304398 303882 304634
rect 303326 268718 303562 268954
rect 303646 268718 303882 268954
rect 303326 268398 303562 268634
rect 303646 268398 303882 268634
rect 307826 708442 308062 708678
rect 308146 708442 308382 708678
rect 307826 708122 308062 708358
rect 308146 708122 308382 708358
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 312326 709402 312562 709638
rect 312646 709402 312882 709638
rect 312326 709082 312562 709318
rect 312646 709082 312882 709318
rect 312326 673718 312562 673954
rect 312646 673718 312882 673954
rect 312326 673398 312562 673634
rect 312646 673398 312882 673634
rect 312326 637718 312562 637954
rect 312646 637718 312882 637954
rect 312326 637398 312562 637634
rect 312646 637398 312882 637634
rect 312326 601718 312562 601954
rect 312646 601718 312882 601954
rect 312326 601398 312562 601634
rect 312646 601398 312882 601634
rect 312326 565718 312562 565954
rect 312646 565718 312882 565954
rect 312326 565398 312562 565634
rect 312646 565398 312882 565634
rect 312326 529718 312562 529954
rect 312646 529718 312882 529954
rect 312326 529398 312562 529634
rect 312646 529398 312882 529634
rect 312326 493718 312562 493954
rect 312646 493718 312882 493954
rect 312326 493398 312562 493634
rect 312646 493398 312882 493634
rect 312326 457718 312562 457954
rect 312646 457718 312882 457954
rect 312326 457398 312562 457634
rect 312646 457398 312882 457634
rect 312326 421718 312562 421954
rect 312646 421718 312882 421954
rect 312326 421398 312562 421634
rect 312646 421398 312882 421634
rect 312326 385718 312562 385954
rect 312646 385718 312882 385954
rect 312326 385398 312562 385634
rect 312646 385398 312882 385634
rect 312326 349718 312562 349954
rect 312646 349718 312882 349954
rect 312326 349398 312562 349634
rect 312646 349398 312882 349634
rect 312326 313718 312562 313954
rect 312646 313718 312882 313954
rect 312326 313398 312562 313634
rect 312646 313398 312882 313634
rect 312326 277718 312562 277954
rect 312646 277718 312882 277954
rect 312326 277398 312562 277634
rect 312646 277398 312882 277634
rect 316826 710362 317062 710598
rect 317146 710362 317382 710598
rect 316826 710042 317062 710278
rect 317146 710042 317382 710278
rect 316826 678218 317062 678454
rect 317146 678218 317382 678454
rect 316826 677898 317062 678134
rect 317146 677898 317382 678134
rect 316826 642218 317062 642454
rect 317146 642218 317382 642454
rect 316826 641898 317062 642134
rect 317146 641898 317382 642134
rect 316826 606218 317062 606454
rect 317146 606218 317382 606454
rect 316826 605898 317062 606134
rect 317146 605898 317382 606134
rect 316826 570218 317062 570454
rect 317146 570218 317382 570454
rect 316826 569898 317062 570134
rect 317146 569898 317382 570134
rect 316826 534218 317062 534454
rect 317146 534218 317382 534454
rect 316826 533898 317062 534134
rect 317146 533898 317382 534134
rect 316826 498218 317062 498454
rect 317146 498218 317382 498454
rect 316826 497898 317062 498134
rect 317146 497898 317382 498134
rect 316826 462218 317062 462454
rect 317146 462218 317382 462454
rect 316826 461898 317062 462134
rect 317146 461898 317382 462134
rect 316826 426218 317062 426454
rect 317146 426218 317382 426454
rect 316826 425898 317062 426134
rect 317146 425898 317382 426134
rect 316826 390218 317062 390454
rect 317146 390218 317382 390454
rect 316826 389898 317062 390134
rect 317146 389898 317382 390134
rect 316826 354218 317062 354454
rect 317146 354218 317382 354454
rect 316826 353898 317062 354134
rect 317146 353898 317382 354134
rect 316826 318218 317062 318454
rect 317146 318218 317382 318454
rect 316826 317898 317062 318134
rect 317146 317898 317382 318134
rect 316826 282218 317062 282454
rect 317146 282218 317382 282454
rect 316826 281898 317062 282134
rect 317146 281898 317382 282134
rect 316826 246218 317062 246454
rect 317146 246218 317382 246454
rect 316826 245898 317062 246134
rect 317146 245898 317382 246134
rect 321326 711322 321562 711558
rect 321646 711322 321882 711558
rect 321326 711002 321562 711238
rect 321646 711002 321882 711238
rect 321326 682718 321562 682954
rect 321646 682718 321882 682954
rect 321326 682398 321562 682634
rect 321646 682398 321882 682634
rect 321326 646718 321562 646954
rect 321646 646718 321882 646954
rect 321326 646398 321562 646634
rect 321646 646398 321882 646634
rect 321326 610718 321562 610954
rect 321646 610718 321882 610954
rect 321326 610398 321562 610634
rect 321646 610398 321882 610634
rect 321326 574718 321562 574954
rect 321646 574718 321882 574954
rect 321326 574398 321562 574634
rect 321646 574398 321882 574634
rect 321326 538718 321562 538954
rect 321646 538718 321882 538954
rect 321326 538398 321562 538634
rect 321646 538398 321882 538634
rect 321326 502718 321562 502954
rect 321646 502718 321882 502954
rect 321326 502398 321562 502634
rect 321646 502398 321882 502634
rect 321326 466718 321562 466954
rect 321646 466718 321882 466954
rect 321326 466398 321562 466634
rect 321646 466398 321882 466634
rect 321326 430718 321562 430954
rect 321646 430718 321882 430954
rect 321326 430398 321562 430634
rect 321646 430398 321882 430634
rect 321326 394718 321562 394954
rect 321646 394718 321882 394954
rect 321326 394398 321562 394634
rect 321646 394398 321882 394634
rect 321326 358718 321562 358954
rect 321646 358718 321882 358954
rect 321326 358398 321562 358634
rect 321646 358398 321882 358634
rect 321326 322718 321562 322954
rect 321646 322718 321882 322954
rect 321326 322398 321562 322634
rect 321646 322398 321882 322634
rect 321326 286718 321562 286954
rect 321646 286718 321882 286954
rect 321326 286398 321562 286634
rect 321646 286398 321882 286634
rect 321326 250718 321562 250954
rect 321646 250718 321882 250954
rect 321326 250398 321562 250634
rect 321646 250398 321882 250634
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 330326 705562 330562 705798
rect 330646 705562 330882 705798
rect 330326 705242 330562 705478
rect 330646 705242 330882 705478
rect 330326 691718 330562 691954
rect 330646 691718 330882 691954
rect 330326 691398 330562 691634
rect 330646 691398 330882 691634
rect 330326 655718 330562 655954
rect 330646 655718 330882 655954
rect 330326 655398 330562 655634
rect 330646 655398 330882 655634
rect 330326 619718 330562 619954
rect 330646 619718 330882 619954
rect 330326 619398 330562 619634
rect 330646 619398 330882 619634
rect 330326 583718 330562 583954
rect 330646 583718 330882 583954
rect 330326 583398 330562 583634
rect 330646 583398 330882 583634
rect 330326 547718 330562 547954
rect 330646 547718 330882 547954
rect 330326 547398 330562 547634
rect 330646 547398 330882 547634
rect 330326 511718 330562 511954
rect 330646 511718 330882 511954
rect 330326 511398 330562 511634
rect 330646 511398 330882 511634
rect 330326 475718 330562 475954
rect 330646 475718 330882 475954
rect 330326 475398 330562 475634
rect 330646 475398 330882 475634
rect 330326 439718 330562 439954
rect 330646 439718 330882 439954
rect 330326 439398 330562 439634
rect 330646 439398 330882 439634
rect 330326 403718 330562 403954
rect 330646 403718 330882 403954
rect 330326 403398 330562 403634
rect 330646 403398 330882 403634
rect 330326 367718 330562 367954
rect 330646 367718 330882 367954
rect 330326 367398 330562 367634
rect 330646 367398 330882 367634
rect 330326 331718 330562 331954
rect 330646 331718 330882 331954
rect 330326 331398 330562 331634
rect 330646 331398 330882 331634
rect 330326 295718 330562 295954
rect 330646 295718 330882 295954
rect 330326 295398 330562 295634
rect 330646 295398 330882 295634
rect 330326 259718 330562 259954
rect 330646 259718 330882 259954
rect 330326 259398 330562 259634
rect 330646 259398 330882 259634
rect 334826 706522 335062 706758
rect 335146 706522 335382 706758
rect 334826 706202 335062 706438
rect 335146 706202 335382 706438
rect 334826 696218 335062 696454
rect 335146 696218 335382 696454
rect 334826 695898 335062 696134
rect 335146 695898 335382 696134
rect 334826 660218 335062 660454
rect 335146 660218 335382 660454
rect 334826 659898 335062 660134
rect 335146 659898 335382 660134
rect 334826 624218 335062 624454
rect 335146 624218 335382 624454
rect 334826 623898 335062 624134
rect 335146 623898 335382 624134
rect 334826 588218 335062 588454
rect 335146 588218 335382 588454
rect 334826 587898 335062 588134
rect 335146 587898 335382 588134
rect 334826 552218 335062 552454
rect 335146 552218 335382 552454
rect 334826 551898 335062 552134
rect 335146 551898 335382 552134
rect 334826 516218 335062 516454
rect 335146 516218 335382 516454
rect 334826 515898 335062 516134
rect 335146 515898 335382 516134
rect 334826 480218 335062 480454
rect 335146 480218 335382 480454
rect 334826 479898 335062 480134
rect 335146 479898 335382 480134
rect 334826 444218 335062 444454
rect 335146 444218 335382 444454
rect 334826 443898 335062 444134
rect 335146 443898 335382 444134
rect 334826 408218 335062 408454
rect 335146 408218 335382 408454
rect 334826 407898 335062 408134
rect 335146 407898 335382 408134
rect 334826 372218 335062 372454
rect 335146 372218 335382 372454
rect 334826 371898 335062 372134
rect 335146 371898 335382 372134
rect 334826 336218 335062 336454
rect 335146 336218 335382 336454
rect 334826 335898 335062 336134
rect 335146 335898 335382 336134
rect 334826 300218 335062 300454
rect 335146 300218 335382 300454
rect 334826 299898 335062 300134
rect 335146 299898 335382 300134
rect 334826 264218 335062 264454
rect 335146 264218 335382 264454
rect 334826 263898 335062 264134
rect 335146 263898 335382 264134
rect 339326 707482 339562 707718
rect 339646 707482 339882 707718
rect 339326 707162 339562 707398
rect 339646 707162 339882 707398
rect 339326 700718 339562 700954
rect 339646 700718 339882 700954
rect 339326 700398 339562 700634
rect 339646 700398 339882 700634
rect 339326 664718 339562 664954
rect 339646 664718 339882 664954
rect 339326 664398 339562 664634
rect 339646 664398 339882 664634
rect 339326 628718 339562 628954
rect 339646 628718 339882 628954
rect 339326 628398 339562 628634
rect 339646 628398 339882 628634
rect 339326 592718 339562 592954
rect 339646 592718 339882 592954
rect 339326 592398 339562 592634
rect 339646 592398 339882 592634
rect 339326 556718 339562 556954
rect 339646 556718 339882 556954
rect 339326 556398 339562 556634
rect 339646 556398 339882 556634
rect 339326 520718 339562 520954
rect 339646 520718 339882 520954
rect 339326 520398 339562 520634
rect 339646 520398 339882 520634
rect 339326 484718 339562 484954
rect 339646 484718 339882 484954
rect 339326 484398 339562 484634
rect 339646 484398 339882 484634
rect 339326 448718 339562 448954
rect 339646 448718 339882 448954
rect 339326 448398 339562 448634
rect 339646 448398 339882 448634
rect 339326 412718 339562 412954
rect 339646 412718 339882 412954
rect 339326 412398 339562 412634
rect 339646 412398 339882 412634
rect 339326 376718 339562 376954
rect 339646 376718 339882 376954
rect 339326 376398 339562 376634
rect 339646 376398 339882 376634
rect 339326 340718 339562 340954
rect 339646 340718 339882 340954
rect 339326 340398 339562 340634
rect 339646 340398 339882 340634
rect 339326 304718 339562 304954
rect 339646 304718 339882 304954
rect 339326 304398 339562 304634
rect 339646 304398 339882 304634
rect 339326 268718 339562 268954
rect 339646 268718 339882 268954
rect 339326 268398 339562 268634
rect 339646 268398 339882 268634
rect 343826 708442 344062 708678
rect 344146 708442 344382 708678
rect 343826 708122 344062 708358
rect 344146 708122 344382 708358
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 348326 709402 348562 709638
rect 348646 709402 348882 709638
rect 348326 709082 348562 709318
rect 348646 709082 348882 709318
rect 348326 673718 348562 673954
rect 348646 673718 348882 673954
rect 348326 673398 348562 673634
rect 348646 673398 348882 673634
rect 348326 637718 348562 637954
rect 348646 637718 348882 637954
rect 348326 637398 348562 637634
rect 348646 637398 348882 637634
rect 348326 601718 348562 601954
rect 348646 601718 348882 601954
rect 348326 601398 348562 601634
rect 348646 601398 348882 601634
rect 348326 565718 348562 565954
rect 348646 565718 348882 565954
rect 348326 565398 348562 565634
rect 348646 565398 348882 565634
rect 348326 529718 348562 529954
rect 348646 529718 348882 529954
rect 348326 529398 348562 529634
rect 348646 529398 348882 529634
rect 348326 493718 348562 493954
rect 348646 493718 348882 493954
rect 348326 493398 348562 493634
rect 348646 493398 348882 493634
rect 348326 457718 348562 457954
rect 348646 457718 348882 457954
rect 348326 457398 348562 457634
rect 348646 457398 348882 457634
rect 348326 421718 348562 421954
rect 348646 421718 348882 421954
rect 348326 421398 348562 421634
rect 348646 421398 348882 421634
rect 348326 385718 348562 385954
rect 348646 385718 348882 385954
rect 348326 385398 348562 385634
rect 348646 385398 348882 385634
rect 348326 349718 348562 349954
rect 348646 349718 348882 349954
rect 348326 349398 348562 349634
rect 348646 349398 348882 349634
rect 348326 313718 348562 313954
rect 348646 313718 348882 313954
rect 348326 313398 348562 313634
rect 348646 313398 348882 313634
rect 348326 277718 348562 277954
rect 348646 277718 348882 277954
rect 348326 277398 348562 277634
rect 348646 277398 348882 277634
rect 352826 710362 353062 710598
rect 353146 710362 353382 710598
rect 352826 710042 353062 710278
rect 353146 710042 353382 710278
rect 352826 678218 353062 678454
rect 353146 678218 353382 678454
rect 352826 677898 353062 678134
rect 353146 677898 353382 678134
rect 352826 642218 353062 642454
rect 353146 642218 353382 642454
rect 352826 641898 353062 642134
rect 353146 641898 353382 642134
rect 352826 606218 353062 606454
rect 353146 606218 353382 606454
rect 352826 605898 353062 606134
rect 353146 605898 353382 606134
rect 352826 570218 353062 570454
rect 353146 570218 353382 570454
rect 352826 569898 353062 570134
rect 353146 569898 353382 570134
rect 352826 534218 353062 534454
rect 353146 534218 353382 534454
rect 352826 533898 353062 534134
rect 353146 533898 353382 534134
rect 352826 498218 353062 498454
rect 353146 498218 353382 498454
rect 352826 497898 353062 498134
rect 353146 497898 353382 498134
rect 352826 462218 353062 462454
rect 353146 462218 353382 462454
rect 352826 461898 353062 462134
rect 353146 461898 353382 462134
rect 352826 426218 353062 426454
rect 353146 426218 353382 426454
rect 352826 425898 353062 426134
rect 353146 425898 353382 426134
rect 352826 390218 353062 390454
rect 353146 390218 353382 390454
rect 352826 389898 353062 390134
rect 353146 389898 353382 390134
rect 352826 354218 353062 354454
rect 353146 354218 353382 354454
rect 352826 353898 353062 354134
rect 353146 353898 353382 354134
rect 352826 318218 353062 318454
rect 353146 318218 353382 318454
rect 352826 317898 353062 318134
rect 353146 317898 353382 318134
rect 352826 282218 353062 282454
rect 353146 282218 353382 282454
rect 352826 281898 353062 282134
rect 353146 281898 353382 282134
rect 352826 246218 353062 246454
rect 353146 246218 353382 246454
rect 352826 245898 353062 246134
rect 353146 245898 353382 246134
rect 357326 711322 357562 711558
rect 357646 711322 357882 711558
rect 357326 711002 357562 711238
rect 357646 711002 357882 711238
rect 357326 682718 357562 682954
rect 357646 682718 357882 682954
rect 357326 682398 357562 682634
rect 357646 682398 357882 682634
rect 357326 646718 357562 646954
rect 357646 646718 357882 646954
rect 357326 646398 357562 646634
rect 357646 646398 357882 646634
rect 357326 610718 357562 610954
rect 357646 610718 357882 610954
rect 357326 610398 357562 610634
rect 357646 610398 357882 610634
rect 357326 574718 357562 574954
rect 357646 574718 357882 574954
rect 357326 574398 357562 574634
rect 357646 574398 357882 574634
rect 357326 538718 357562 538954
rect 357646 538718 357882 538954
rect 357326 538398 357562 538634
rect 357646 538398 357882 538634
rect 357326 502718 357562 502954
rect 357646 502718 357882 502954
rect 357326 502398 357562 502634
rect 357646 502398 357882 502634
rect 357326 466718 357562 466954
rect 357646 466718 357882 466954
rect 357326 466398 357562 466634
rect 357646 466398 357882 466634
rect 357326 430718 357562 430954
rect 357646 430718 357882 430954
rect 357326 430398 357562 430634
rect 357646 430398 357882 430634
rect 357326 394718 357562 394954
rect 357646 394718 357882 394954
rect 357326 394398 357562 394634
rect 357646 394398 357882 394634
rect 357326 358718 357562 358954
rect 357646 358718 357882 358954
rect 357326 358398 357562 358634
rect 357646 358398 357882 358634
rect 357326 322718 357562 322954
rect 357646 322718 357882 322954
rect 357326 322398 357562 322634
rect 357646 322398 357882 322634
rect 357326 286718 357562 286954
rect 357646 286718 357882 286954
rect 357326 286398 357562 286634
rect 357646 286398 357882 286634
rect 357326 250718 357562 250954
rect 357646 250718 357882 250954
rect 357326 250398 357562 250634
rect 357646 250398 357882 250634
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 366326 705562 366562 705798
rect 366646 705562 366882 705798
rect 366326 705242 366562 705478
rect 366646 705242 366882 705478
rect 366326 691718 366562 691954
rect 366646 691718 366882 691954
rect 366326 691398 366562 691634
rect 366646 691398 366882 691634
rect 366326 655718 366562 655954
rect 366646 655718 366882 655954
rect 366326 655398 366562 655634
rect 366646 655398 366882 655634
rect 366326 619718 366562 619954
rect 366646 619718 366882 619954
rect 366326 619398 366562 619634
rect 366646 619398 366882 619634
rect 366326 583718 366562 583954
rect 366646 583718 366882 583954
rect 366326 583398 366562 583634
rect 366646 583398 366882 583634
rect 366326 547718 366562 547954
rect 366646 547718 366882 547954
rect 366326 547398 366562 547634
rect 366646 547398 366882 547634
rect 366326 511718 366562 511954
rect 366646 511718 366882 511954
rect 366326 511398 366562 511634
rect 366646 511398 366882 511634
rect 366326 475718 366562 475954
rect 366646 475718 366882 475954
rect 366326 475398 366562 475634
rect 366646 475398 366882 475634
rect 366326 439718 366562 439954
rect 366646 439718 366882 439954
rect 366326 439398 366562 439634
rect 366646 439398 366882 439634
rect 366326 403718 366562 403954
rect 366646 403718 366882 403954
rect 366326 403398 366562 403634
rect 366646 403398 366882 403634
rect 366326 367718 366562 367954
rect 366646 367718 366882 367954
rect 366326 367398 366562 367634
rect 366646 367398 366882 367634
rect 366326 331718 366562 331954
rect 366646 331718 366882 331954
rect 366326 331398 366562 331634
rect 366646 331398 366882 331634
rect 366326 295718 366562 295954
rect 366646 295718 366882 295954
rect 366326 295398 366562 295634
rect 366646 295398 366882 295634
rect 366326 259718 366562 259954
rect 366646 259718 366882 259954
rect 366326 259398 366562 259634
rect 366646 259398 366882 259634
rect 370826 706522 371062 706758
rect 371146 706522 371382 706758
rect 370826 706202 371062 706438
rect 371146 706202 371382 706438
rect 370826 696218 371062 696454
rect 371146 696218 371382 696454
rect 370826 695898 371062 696134
rect 371146 695898 371382 696134
rect 370826 660218 371062 660454
rect 371146 660218 371382 660454
rect 370826 659898 371062 660134
rect 371146 659898 371382 660134
rect 370826 624218 371062 624454
rect 371146 624218 371382 624454
rect 370826 623898 371062 624134
rect 371146 623898 371382 624134
rect 370826 588218 371062 588454
rect 371146 588218 371382 588454
rect 370826 587898 371062 588134
rect 371146 587898 371382 588134
rect 370826 552218 371062 552454
rect 371146 552218 371382 552454
rect 370826 551898 371062 552134
rect 371146 551898 371382 552134
rect 370826 516218 371062 516454
rect 371146 516218 371382 516454
rect 370826 515898 371062 516134
rect 371146 515898 371382 516134
rect 370826 480218 371062 480454
rect 371146 480218 371382 480454
rect 370826 479898 371062 480134
rect 371146 479898 371382 480134
rect 370826 444218 371062 444454
rect 371146 444218 371382 444454
rect 370826 443898 371062 444134
rect 371146 443898 371382 444134
rect 370826 408218 371062 408454
rect 371146 408218 371382 408454
rect 370826 407898 371062 408134
rect 371146 407898 371382 408134
rect 370826 372218 371062 372454
rect 371146 372218 371382 372454
rect 370826 371898 371062 372134
rect 371146 371898 371382 372134
rect 370826 336218 371062 336454
rect 371146 336218 371382 336454
rect 370826 335898 371062 336134
rect 371146 335898 371382 336134
rect 370826 300218 371062 300454
rect 371146 300218 371382 300454
rect 370826 299898 371062 300134
rect 371146 299898 371382 300134
rect 370826 264218 371062 264454
rect 371146 264218 371382 264454
rect 370826 263898 371062 264134
rect 371146 263898 371382 264134
rect 375326 707482 375562 707718
rect 375646 707482 375882 707718
rect 375326 707162 375562 707398
rect 375646 707162 375882 707398
rect 375326 700718 375562 700954
rect 375646 700718 375882 700954
rect 375326 700398 375562 700634
rect 375646 700398 375882 700634
rect 375326 664718 375562 664954
rect 375646 664718 375882 664954
rect 375326 664398 375562 664634
rect 375646 664398 375882 664634
rect 375326 628718 375562 628954
rect 375646 628718 375882 628954
rect 375326 628398 375562 628634
rect 375646 628398 375882 628634
rect 375326 592718 375562 592954
rect 375646 592718 375882 592954
rect 375326 592398 375562 592634
rect 375646 592398 375882 592634
rect 375326 556718 375562 556954
rect 375646 556718 375882 556954
rect 375326 556398 375562 556634
rect 375646 556398 375882 556634
rect 375326 520718 375562 520954
rect 375646 520718 375882 520954
rect 375326 520398 375562 520634
rect 375646 520398 375882 520634
rect 375326 484718 375562 484954
rect 375646 484718 375882 484954
rect 375326 484398 375562 484634
rect 375646 484398 375882 484634
rect 375326 448718 375562 448954
rect 375646 448718 375882 448954
rect 375326 448398 375562 448634
rect 375646 448398 375882 448634
rect 375326 412718 375562 412954
rect 375646 412718 375882 412954
rect 375326 412398 375562 412634
rect 375646 412398 375882 412634
rect 375326 376718 375562 376954
rect 375646 376718 375882 376954
rect 375326 376398 375562 376634
rect 375646 376398 375882 376634
rect 375326 340718 375562 340954
rect 375646 340718 375882 340954
rect 375326 340398 375562 340634
rect 375646 340398 375882 340634
rect 375326 304718 375562 304954
rect 375646 304718 375882 304954
rect 375326 304398 375562 304634
rect 375646 304398 375882 304634
rect 375326 268718 375562 268954
rect 375646 268718 375882 268954
rect 375326 268398 375562 268634
rect 375646 268398 375882 268634
rect 379826 708442 380062 708678
rect 380146 708442 380382 708678
rect 379826 708122 380062 708358
rect 380146 708122 380382 708358
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 384326 709402 384562 709638
rect 384646 709402 384882 709638
rect 384326 709082 384562 709318
rect 384646 709082 384882 709318
rect 384326 673718 384562 673954
rect 384646 673718 384882 673954
rect 384326 673398 384562 673634
rect 384646 673398 384882 673634
rect 384326 637718 384562 637954
rect 384646 637718 384882 637954
rect 384326 637398 384562 637634
rect 384646 637398 384882 637634
rect 384326 601718 384562 601954
rect 384646 601718 384882 601954
rect 384326 601398 384562 601634
rect 384646 601398 384882 601634
rect 384326 565718 384562 565954
rect 384646 565718 384882 565954
rect 384326 565398 384562 565634
rect 384646 565398 384882 565634
rect 384326 529718 384562 529954
rect 384646 529718 384882 529954
rect 384326 529398 384562 529634
rect 384646 529398 384882 529634
rect 384326 493718 384562 493954
rect 384646 493718 384882 493954
rect 384326 493398 384562 493634
rect 384646 493398 384882 493634
rect 384326 457718 384562 457954
rect 384646 457718 384882 457954
rect 384326 457398 384562 457634
rect 384646 457398 384882 457634
rect 384326 421718 384562 421954
rect 384646 421718 384882 421954
rect 384326 421398 384562 421634
rect 384646 421398 384882 421634
rect 384326 385718 384562 385954
rect 384646 385718 384882 385954
rect 384326 385398 384562 385634
rect 384646 385398 384882 385634
rect 384326 349718 384562 349954
rect 384646 349718 384882 349954
rect 384326 349398 384562 349634
rect 384646 349398 384882 349634
rect 384326 313718 384562 313954
rect 384646 313718 384882 313954
rect 384326 313398 384562 313634
rect 384646 313398 384882 313634
rect 384326 277718 384562 277954
rect 384646 277718 384882 277954
rect 384326 277398 384562 277634
rect 384646 277398 384882 277634
rect 388826 710362 389062 710598
rect 389146 710362 389382 710598
rect 388826 710042 389062 710278
rect 389146 710042 389382 710278
rect 388826 678218 389062 678454
rect 389146 678218 389382 678454
rect 388826 677898 389062 678134
rect 389146 677898 389382 678134
rect 388826 642218 389062 642454
rect 389146 642218 389382 642454
rect 388826 641898 389062 642134
rect 389146 641898 389382 642134
rect 388826 606218 389062 606454
rect 389146 606218 389382 606454
rect 388826 605898 389062 606134
rect 389146 605898 389382 606134
rect 388826 570218 389062 570454
rect 389146 570218 389382 570454
rect 388826 569898 389062 570134
rect 389146 569898 389382 570134
rect 388826 534218 389062 534454
rect 389146 534218 389382 534454
rect 388826 533898 389062 534134
rect 389146 533898 389382 534134
rect 388826 498218 389062 498454
rect 389146 498218 389382 498454
rect 388826 497898 389062 498134
rect 389146 497898 389382 498134
rect 388826 462218 389062 462454
rect 389146 462218 389382 462454
rect 388826 461898 389062 462134
rect 389146 461898 389382 462134
rect 388826 426218 389062 426454
rect 389146 426218 389382 426454
rect 388826 425898 389062 426134
rect 389146 425898 389382 426134
rect 388826 390218 389062 390454
rect 389146 390218 389382 390454
rect 388826 389898 389062 390134
rect 389146 389898 389382 390134
rect 388826 354218 389062 354454
rect 389146 354218 389382 354454
rect 388826 353898 389062 354134
rect 389146 353898 389382 354134
rect 388826 318218 389062 318454
rect 389146 318218 389382 318454
rect 388826 317898 389062 318134
rect 389146 317898 389382 318134
rect 388826 282218 389062 282454
rect 389146 282218 389382 282454
rect 388826 281898 389062 282134
rect 389146 281898 389382 282134
rect 388826 246218 389062 246454
rect 389146 246218 389382 246454
rect 388826 245898 389062 246134
rect 389146 245898 389382 246134
rect 393326 711322 393562 711558
rect 393646 711322 393882 711558
rect 393326 711002 393562 711238
rect 393646 711002 393882 711238
rect 393326 682718 393562 682954
rect 393646 682718 393882 682954
rect 393326 682398 393562 682634
rect 393646 682398 393882 682634
rect 393326 646718 393562 646954
rect 393646 646718 393882 646954
rect 393326 646398 393562 646634
rect 393646 646398 393882 646634
rect 393326 610718 393562 610954
rect 393646 610718 393882 610954
rect 393326 610398 393562 610634
rect 393646 610398 393882 610634
rect 393326 574718 393562 574954
rect 393646 574718 393882 574954
rect 393326 574398 393562 574634
rect 393646 574398 393882 574634
rect 393326 538718 393562 538954
rect 393646 538718 393882 538954
rect 393326 538398 393562 538634
rect 393646 538398 393882 538634
rect 393326 502718 393562 502954
rect 393646 502718 393882 502954
rect 393326 502398 393562 502634
rect 393646 502398 393882 502634
rect 393326 466718 393562 466954
rect 393646 466718 393882 466954
rect 393326 466398 393562 466634
rect 393646 466398 393882 466634
rect 393326 430718 393562 430954
rect 393646 430718 393882 430954
rect 393326 430398 393562 430634
rect 393646 430398 393882 430634
rect 393326 394718 393562 394954
rect 393646 394718 393882 394954
rect 393326 394398 393562 394634
rect 393646 394398 393882 394634
rect 393326 358718 393562 358954
rect 393646 358718 393882 358954
rect 393326 358398 393562 358634
rect 393646 358398 393882 358634
rect 393326 322718 393562 322954
rect 393646 322718 393882 322954
rect 393326 322398 393562 322634
rect 393646 322398 393882 322634
rect 393326 286718 393562 286954
rect 393646 286718 393882 286954
rect 393326 286398 393562 286634
rect 393646 286398 393882 286634
rect 393326 250718 393562 250954
rect 393646 250718 393882 250954
rect 393326 250398 393562 250634
rect 393646 250398 393882 250634
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 402326 705562 402562 705798
rect 402646 705562 402882 705798
rect 402326 705242 402562 705478
rect 402646 705242 402882 705478
rect 402326 691718 402562 691954
rect 402646 691718 402882 691954
rect 402326 691398 402562 691634
rect 402646 691398 402882 691634
rect 402326 655718 402562 655954
rect 402646 655718 402882 655954
rect 402326 655398 402562 655634
rect 402646 655398 402882 655634
rect 402326 619718 402562 619954
rect 402646 619718 402882 619954
rect 402326 619398 402562 619634
rect 402646 619398 402882 619634
rect 402326 583718 402562 583954
rect 402646 583718 402882 583954
rect 402326 583398 402562 583634
rect 402646 583398 402882 583634
rect 402326 547718 402562 547954
rect 402646 547718 402882 547954
rect 402326 547398 402562 547634
rect 402646 547398 402882 547634
rect 402326 511718 402562 511954
rect 402646 511718 402882 511954
rect 402326 511398 402562 511634
rect 402646 511398 402882 511634
rect 402326 475718 402562 475954
rect 402646 475718 402882 475954
rect 402326 475398 402562 475634
rect 402646 475398 402882 475634
rect 402326 439718 402562 439954
rect 402646 439718 402882 439954
rect 402326 439398 402562 439634
rect 402646 439398 402882 439634
rect 402326 403718 402562 403954
rect 402646 403718 402882 403954
rect 402326 403398 402562 403634
rect 402646 403398 402882 403634
rect 402326 367718 402562 367954
rect 402646 367718 402882 367954
rect 402326 367398 402562 367634
rect 402646 367398 402882 367634
rect 402326 331718 402562 331954
rect 402646 331718 402882 331954
rect 402326 331398 402562 331634
rect 402646 331398 402882 331634
rect 402326 295718 402562 295954
rect 402646 295718 402882 295954
rect 402326 295398 402562 295634
rect 402646 295398 402882 295634
rect 402326 259718 402562 259954
rect 402646 259718 402882 259954
rect 402326 259398 402562 259634
rect 402646 259398 402882 259634
rect 406826 706522 407062 706758
rect 407146 706522 407382 706758
rect 406826 706202 407062 706438
rect 407146 706202 407382 706438
rect 406826 696218 407062 696454
rect 407146 696218 407382 696454
rect 406826 695898 407062 696134
rect 407146 695898 407382 696134
rect 406826 660218 407062 660454
rect 407146 660218 407382 660454
rect 406826 659898 407062 660134
rect 407146 659898 407382 660134
rect 406826 624218 407062 624454
rect 407146 624218 407382 624454
rect 406826 623898 407062 624134
rect 407146 623898 407382 624134
rect 406826 588218 407062 588454
rect 407146 588218 407382 588454
rect 406826 587898 407062 588134
rect 407146 587898 407382 588134
rect 406826 552218 407062 552454
rect 407146 552218 407382 552454
rect 406826 551898 407062 552134
rect 407146 551898 407382 552134
rect 406826 516218 407062 516454
rect 407146 516218 407382 516454
rect 406826 515898 407062 516134
rect 407146 515898 407382 516134
rect 406826 480218 407062 480454
rect 407146 480218 407382 480454
rect 406826 479898 407062 480134
rect 407146 479898 407382 480134
rect 406826 444218 407062 444454
rect 407146 444218 407382 444454
rect 406826 443898 407062 444134
rect 407146 443898 407382 444134
rect 406826 408218 407062 408454
rect 407146 408218 407382 408454
rect 406826 407898 407062 408134
rect 407146 407898 407382 408134
rect 406826 372218 407062 372454
rect 407146 372218 407382 372454
rect 406826 371898 407062 372134
rect 407146 371898 407382 372134
rect 406826 336218 407062 336454
rect 407146 336218 407382 336454
rect 406826 335898 407062 336134
rect 407146 335898 407382 336134
rect 406826 300218 407062 300454
rect 407146 300218 407382 300454
rect 406826 299898 407062 300134
rect 407146 299898 407382 300134
rect 406826 264218 407062 264454
rect 407146 264218 407382 264454
rect 406826 263898 407062 264134
rect 407146 263898 407382 264134
rect 71462 241717 71698 241953
rect 71782 241717 72018 241953
rect 72102 241717 72338 241953
rect 72422 241717 72658 241953
rect 72742 241717 72978 241953
rect 73062 241717 73298 241953
rect 73382 241717 73618 241953
rect 73702 241717 73938 241953
rect 74022 241717 74258 241953
rect 74342 241717 74578 241953
rect 74662 241717 74898 241953
rect 74982 241717 75218 241953
rect 75302 241717 75538 241953
rect 75622 241717 75858 241953
rect 75942 241717 76178 241953
rect 76262 241717 76498 241953
rect 76582 241717 76818 241953
rect 76902 241717 77138 241953
rect 71462 241397 71698 241633
rect 71782 241397 72018 241633
rect 72102 241397 72338 241633
rect 72422 241397 72658 241633
rect 72742 241397 72978 241633
rect 73062 241397 73298 241633
rect 73382 241397 73618 241633
rect 73702 241397 73938 241633
rect 74022 241397 74258 241633
rect 74342 241397 74578 241633
rect 74662 241397 74898 241633
rect 74982 241397 75218 241633
rect 75302 241397 75538 241633
rect 75622 241397 75858 241633
rect 75942 241397 76178 241633
rect 76262 241397 76498 241633
rect 76582 241397 76818 241633
rect 76902 241397 77138 241633
rect 46039 237217 46275 237453
rect 46359 237217 46595 237453
rect 46679 237217 46915 237453
rect 46999 237217 47235 237453
rect 47319 237217 47555 237453
rect 47639 237217 47875 237453
rect 47959 237217 48195 237453
rect 48279 237217 48515 237453
rect 48599 237217 48835 237453
rect 48919 237217 49155 237453
rect 49239 237217 49475 237453
rect 49559 237217 49795 237453
rect 49879 237217 50115 237453
rect 50199 237217 50435 237453
rect 50519 237217 50755 237453
rect 46039 236897 46275 237133
rect 46359 236897 46595 237133
rect 46679 236897 46915 237133
rect 46999 236897 47235 237133
rect 47319 236897 47555 237133
rect 47639 236897 47875 237133
rect 47959 236897 48195 237133
rect 48279 236897 48515 237133
rect 48599 236897 48835 237133
rect 48919 236897 49155 237133
rect 49239 236897 49475 237133
rect 49559 236897 49795 237133
rect 49879 236897 50115 237133
rect 50199 236897 50435 237133
rect 50519 236897 50755 237133
rect 42326 223718 42562 223954
rect 42646 223718 42882 223954
rect 42326 223398 42562 223634
rect 42646 223398 42882 223634
rect 42326 187718 42562 187954
rect 42646 187718 42882 187954
rect 42326 187398 42562 187634
rect 42646 187398 42882 187634
rect 42326 151718 42562 151954
rect 42646 151718 42882 151954
rect 42326 151398 42562 151634
rect 42646 151398 42882 151634
rect 42326 115718 42562 115954
rect 42646 115718 42882 115954
rect 42326 115398 42562 115634
rect 42646 115398 42882 115634
rect 42326 79718 42562 79954
rect 42646 79718 42882 79954
rect 42326 79398 42562 79634
rect 42646 79398 42882 79634
rect 42326 43718 42562 43954
rect 42646 43718 42882 43954
rect 42326 43398 42562 43634
rect 42646 43398 42882 43634
rect 42326 7718 42562 7954
rect 42646 7718 42882 7954
rect 42326 7398 42562 7634
rect 42646 7398 42882 7634
rect 42326 -1542 42562 -1306
rect 42646 -1542 42882 -1306
rect 42326 -1862 42562 -1626
rect 42646 -1862 42882 -1626
rect 46826 228217 47062 228453
rect 47146 228217 47382 228453
rect 46826 227897 47062 228133
rect 47146 227897 47382 228133
rect 46826 192218 47062 192454
rect 47146 192218 47382 192454
rect 46826 191898 47062 192134
rect 47146 191898 47382 192134
rect 46826 156218 47062 156454
rect 47146 156218 47382 156454
rect 46826 155898 47062 156134
rect 47146 155898 47382 156134
rect 46826 120218 47062 120454
rect 47146 120218 47382 120454
rect 46826 119898 47062 120134
rect 47146 119898 47382 120134
rect 46826 84218 47062 84454
rect 47146 84218 47382 84454
rect 46826 83898 47062 84134
rect 47146 83898 47382 84134
rect 46826 48218 47062 48454
rect 47146 48218 47382 48454
rect 46826 47898 47062 48134
rect 47146 47898 47382 48134
rect 46826 12218 47062 12454
rect 47146 12218 47382 12454
rect 46826 11898 47062 12134
rect 47146 11898 47382 12134
rect 46826 -2502 47062 -2266
rect 47146 -2502 47382 -2266
rect 46826 -2822 47062 -2586
rect 47146 -2822 47382 -2586
rect 51326 196718 51562 196954
rect 51646 196718 51882 196954
rect 51326 196398 51562 196634
rect 51646 196398 51882 196634
rect 51326 160718 51562 160954
rect 51646 160718 51882 160954
rect 51326 160398 51562 160634
rect 51646 160398 51882 160634
rect 51326 124718 51562 124954
rect 51646 124718 51882 124954
rect 51326 124398 51562 124634
rect 51646 124398 51882 124634
rect 51326 88718 51562 88954
rect 51646 88718 51882 88954
rect 51326 88398 51562 88634
rect 51646 88398 51882 88634
rect 51326 52718 51562 52954
rect 51646 52718 51882 52954
rect 51326 52398 51562 52634
rect 51646 52398 51882 52634
rect 51326 16718 51562 16954
rect 51646 16718 51882 16954
rect 51326 16398 51562 16634
rect 51646 16398 51882 16634
rect 51326 -3462 51562 -3226
rect 51646 -3462 51882 -3226
rect 51326 -3782 51562 -3546
rect 51646 -3782 51882 -3546
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -4422 56062 -4186
rect 56146 -4422 56382 -4186
rect 55826 -4742 56062 -4506
rect 56146 -4742 56382 -4506
rect 60326 205718 60562 205954
rect 60646 205718 60882 205954
rect 60326 205398 60562 205634
rect 60646 205398 60882 205634
rect 60326 169718 60562 169954
rect 60646 169718 60882 169954
rect 60326 169398 60562 169634
rect 60646 169398 60882 169634
rect 60326 133718 60562 133954
rect 60646 133718 60882 133954
rect 60326 133398 60562 133634
rect 60646 133398 60882 133634
rect 60326 97718 60562 97954
rect 60646 97718 60882 97954
rect 60326 97398 60562 97634
rect 60646 97398 60882 97634
rect 60326 61718 60562 61954
rect 60646 61718 60882 61954
rect 60326 61398 60562 61634
rect 60646 61398 60882 61634
rect 60326 25718 60562 25954
rect 60646 25718 60882 25954
rect 60326 25398 60562 25634
rect 60646 25398 60882 25634
rect 60326 -5382 60562 -5146
rect 60646 -5382 60882 -5146
rect 60326 -5702 60562 -5466
rect 60646 -5702 60882 -5466
rect 64826 210218 65062 210454
rect 65146 210218 65382 210454
rect 64826 209898 65062 210134
rect 65146 209898 65382 210134
rect 64826 174218 65062 174454
rect 65146 174218 65382 174454
rect 64826 173898 65062 174134
rect 65146 173898 65382 174134
rect 64826 138218 65062 138454
rect 65146 138218 65382 138454
rect 64826 137898 65062 138134
rect 65146 137898 65382 138134
rect 64826 102218 65062 102454
rect 65146 102218 65382 102454
rect 64826 101898 65062 102134
rect 65146 101898 65382 102134
rect 64826 66218 65062 66454
rect 65146 66218 65382 66454
rect 64826 65898 65062 66134
rect 65146 65898 65382 66134
rect 64826 30218 65062 30454
rect 65146 30218 65382 30454
rect 64826 29898 65062 30134
rect 65146 29898 65382 30134
rect 64826 -6342 65062 -6106
rect 65146 -6342 65382 -6106
rect 64826 -6662 65062 -6426
rect 65146 -6662 65382 -6426
rect 69326 214718 69562 214954
rect 69646 214718 69882 214954
rect 69326 214398 69562 214634
rect 69646 214398 69882 214634
rect 69326 178718 69562 178954
rect 69646 178718 69882 178954
rect 69326 178398 69562 178634
rect 69646 178398 69882 178634
rect 69326 142718 69562 142954
rect 69646 142718 69882 142954
rect 69326 142398 69562 142634
rect 69646 142398 69882 142634
rect 69326 106718 69562 106954
rect 69646 106718 69882 106954
rect 69326 106398 69562 106634
rect 69646 106398 69882 106634
rect 69326 70718 69562 70954
rect 69646 70718 69882 70954
rect 69326 70398 69562 70634
rect 69646 70398 69882 70634
rect 69326 34718 69562 34954
rect 69646 34718 69882 34954
rect 69326 34398 69562 34634
rect 69646 34398 69882 34634
rect 69326 -7302 69562 -7066
rect 69646 -7302 69882 -7066
rect 69326 -7622 69562 -7386
rect 69646 -7622 69882 -7386
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 78326 223718 78562 223954
rect 78646 223718 78882 223954
rect 78326 223398 78562 223634
rect 78646 223398 78882 223634
rect 78326 187718 78562 187954
rect 78646 187718 78882 187954
rect 78326 187398 78562 187634
rect 78646 187398 78882 187634
rect 78326 151718 78562 151954
rect 78646 151718 78882 151954
rect 78326 151398 78562 151634
rect 78646 151398 78882 151634
rect 78326 115718 78562 115954
rect 78646 115718 78882 115954
rect 78326 115398 78562 115634
rect 78646 115398 78882 115634
rect 78326 79718 78562 79954
rect 78646 79718 78882 79954
rect 78326 79398 78562 79634
rect 78646 79398 78882 79634
rect 78326 43718 78562 43954
rect 78646 43718 78882 43954
rect 78326 43398 78562 43634
rect 78646 43398 78882 43634
rect 78326 7718 78562 7954
rect 78646 7718 78882 7954
rect 78326 7398 78562 7634
rect 78646 7398 78882 7634
rect 78326 -1542 78562 -1306
rect 78646 -1542 78882 -1306
rect 78326 -1862 78562 -1626
rect 78646 -1862 78882 -1626
rect 82826 228217 83062 228453
rect 83146 228217 83382 228453
rect 82826 227897 83062 228133
rect 83146 227897 83382 228133
rect 82826 192218 83062 192454
rect 83146 192218 83382 192454
rect 82826 191898 83062 192134
rect 83146 191898 83382 192134
rect 82826 156218 83062 156454
rect 83146 156218 83382 156454
rect 82826 155898 83062 156134
rect 83146 155898 83382 156134
rect 82826 120218 83062 120454
rect 83146 120218 83382 120454
rect 82826 119898 83062 120134
rect 83146 119898 83382 120134
rect 82826 84218 83062 84454
rect 83146 84218 83382 84454
rect 82826 83898 83062 84134
rect 83146 83898 83382 84134
rect 82826 48218 83062 48454
rect 83146 48218 83382 48454
rect 82826 47898 83062 48134
rect 83146 47898 83382 48134
rect 82826 12218 83062 12454
rect 83146 12218 83382 12454
rect 82826 11898 83062 12134
rect 83146 11898 83382 12134
rect 82826 -2502 83062 -2266
rect 83146 -2502 83382 -2266
rect 82826 -2822 83062 -2586
rect 83146 -2822 83382 -2586
rect 87326 196718 87562 196954
rect 87646 196718 87882 196954
rect 87326 196398 87562 196634
rect 87646 196398 87882 196634
rect 87326 160718 87562 160954
rect 87646 160718 87882 160954
rect 87326 160398 87562 160634
rect 87646 160398 87882 160634
rect 87326 124718 87562 124954
rect 87646 124718 87882 124954
rect 87326 124398 87562 124634
rect 87646 124398 87882 124634
rect 87326 88718 87562 88954
rect 87646 88718 87882 88954
rect 87326 88398 87562 88634
rect 87646 88398 87882 88634
rect 87326 52718 87562 52954
rect 87646 52718 87882 52954
rect 87326 52398 87562 52634
rect 87646 52398 87882 52634
rect 87326 16718 87562 16954
rect 87646 16718 87882 16954
rect 87326 16398 87562 16634
rect 87646 16398 87882 16634
rect 87326 -3462 87562 -3226
rect 87646 -3462 87882 -3226
rect 87326 -3782 87562 -3546
rect 87646 -3782 87882 -3546
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 91826 129218 92062 129454
rect 92146 129218 92382 129454
rect 91826 128898 92062 129134
rect 92146 128898 92382 129134
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -4422 92062 -4186
rect 92146 -4422 92382 -4186
rect 91826 -4742 92062 -4506
rect 92146 -4742 92382 -4506
rect 96326 205718 96562 205954
rect 96646 205718 96882 205954
rect 96326 205398 96562 205634
rect 96646 205398 96882 205634
rect 96326 169718 96562 169954
rect 96646 169718 96882 169954
rect 96326 169398 96562 169634
rect 96646 169398 96882 169634
rect 96326 133718 96562 133954
rect 96646 133718 96882 133954
rect 96326 133398 96562 133634
rect 96646 133398 96882 133634
rect 96326 97718 96562 97954
rect 96646 97718 96882 97954
rect 96326 97398 96562 97634
rect 96646 97398 96882 97634
rect 96326 61718 96562 61954
rect 96646 61718 96882 61954
rect 96326 61398 96562 61634
rect 96646 61398 96882 61634
rect 96326 25718 96562 25954
rect 96646 25718 96882 25954
rect 96326 25398 96562 25634
rect 96646 25398 96882 25634
rect 96326 -5382 96562 -5146
rect 96646 -5382 96882 -5146
rect 96326 -5702 96562 -5466
rect 96646 -5702 96882 -5466
rect 100826 210218 101062 210454
rect 101146 210218 101382 210454
rect 100826 209898 101062 210134
rect 101146 209898 101382 210134
rect 100826 174218 101062 174454
rect 101146 174218 101382 174454
rect 100826 173898 101062 174134
rect 101146 173898 101382 174134
rect 100826 138218 101062 138454
rect 101146 138218 101382 138454
rect 100826 137898 101062 138134
rect 101146 137898 101382 138134
rect 100826 102218 101062 102454
rect 101146 102218 101382 102454
rect 100826 101898 101062 102134
rect 101146 101898 101382 102134
rect 100826 66218 101062 66454
rect 101146 66218 101382 66454
rect 100826 65898 101062 66134
rect 101146 65898 101382 66134
rect 100826 30218 101062 30454
rect 101146 30218 101382 30454
rect 100826 29898 101062 30134
rect 101146 29898 101382 30134
rect 100826 -6342 101062 -6106
rect 101146 -6342 101382 -6106
rect 100826 -6662 101062 -6426
rect 101146 -6662 101382 -6426
rect 105326 214718 105562 214954
rect 105646 214718 105882 214954
rect 105326 214398 105562 214634
rect 105646 214398 105882 214634
rect 105326 178718 105562 178954
rect 105646 178718 105882 178954
rect 105326 178398 105562 178634
rect 105646 178398 105882 178634
rect 105326 142718 105562 142954
rect 105646 142718 105882 142954
rect 105326 142398 105562 142634
rect 105646 142398 105882 142634
rect 105326 106718 105562 106954
rect 105646 106718 105882 106954
rect 105326 106398 105562 106634
rect 105646 106398 105882 106634
rect 105326 70718 105562 70954
rect 105646 70718 105882 70954
rect 105326 70398 105562 70634
rect 105646 70398 105882 70634
rect 105326 34718 105562 34954
rect 105646 34718 105882 34954
rect 105326 34398 105562 34634
rect 105646 34398 105882 34634
rect 105326 -7302 105562 -7066
rect 105646 -7302 105882 -7066
rect 105326 -7622 105562 -7386
rect 105646 -7622 105882 -7386
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 114326 223718 114562 223954
rect 114646 223718 114882 223954
rect 114326 223398 114562 223634
rect 114646 223398 114882 223634
rect 114326 187718 114562 187954
rect 114646 187718 114882 187954
rect 114326 187398 114562 187634
rect 114646 187398 114882 187634
rect 114326 151718 114562 151954
rect 114646 151718 114882 151954
rect 114326 151398 114562 151634
rect 114646 151398 114882 151634
rect 118826 228217 119062 228453
rect 119146 228217 119382 228453
rect 118826 227897 119062 228133
rect 119146 227897 119382 228133
rect 118826 192218 119062 192454
rect 119146 192218 119382 192454
rect 118826 191898 119062 192134
rect 119146 191898 119382 192134
rect 118826 156218 119062 156454
rect 119146 156218 119382 156454
rect 118826 155898 119062 156134
rect 119146 155898 119382 156134
rect 123326 196718 123562 196954
rect 123646 196718 123882 196954
rect 123326 196398 123562 196634
rect 123646 196398 123882 196634
rect 123326 160718 123562 160954
rect 123646 160718 123882 160954
rect 123326 160398 123562 160634
rect 123646 160398 123882 160634
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 127826 165218 128062 165454
rect 128146 165218 128382 165454
rect 127826 164898 128062 165134
rect 128146 164898 128382 165134
rect 132326 205718 132562 205954
rect 132646 205718 132882 205954
rect 132326 205398 132562 205634
rect 132646 205398 132882 205634
rect 136036 205718 136272 205954
rect 136356 205718 136592 205954
rect 136676 205718 136912 205954
rect 136996 205718 137232 205954
rect 137316 205718 137552 205954
rect 137636 205718 137872 205954
rect 137956 205718 138192 205954
rect 138276 205718 138512 205954
rect 138596 205718 138832 205954
rect 138916 205718 139152 205954
rect 139236 205718 139472 205954
rect 139556 205718 139792 205954
rect 139876 205718 140112 205954
rect 140196 205718 140432 205954
rect 140516 205718 140752 205954
rect 140836 205718 141072 205954
rect 141156 205718 141392 205954
rect 141476 205718 141712 205954
rect 141796 205718 142032 205954
rect 142116 205718 142352 205954
rect 142436 205718 142672 205954
rect 142756 205718 142992 205954
rect 143076 205718 143312 205954
rect 143396 205718 143632 205954
rect 143716 205718 143952 205954
rect 144036 205718 144272 205954
rect 144356 205718 144592 205954
rect 144676 205718 144912 205954
rect 144996 205718 145232 205954
rect 145316 205718 145552 205954
rect 145636 205718 145872 205954
rect 145956 205718 146192 205954
rect 146276 205718 146512 205954
rect 146596 205718 146832 205954
rect 146916 205718 147152 205954
rect 147236 205718 147472 205954
rect 147556 205718 147792 205954
rect 147876 205718 148112 205954
rect 148196 205718 148432 205954
rect 148516 205718 148752 205954
rect 148836 205718 149072 205954
rect 149156 205718 149392 205954
rect 149476 205718 149712 205954
rect 149796 205718 150032 205954
rect 150116 205718 150352 205954
rect 150436 205718 150672 205954
rect 150756 205718 150992 205954
rect 151076 205718 151312 205954
rect 151396 205718 151632 205954
rect 151716 205718 151952 205954
rect 152036 205718 152272 205954
rect 152356 205718 152592 205954
rect 152676 205718 152912 205954
rect 152996 205718 153232 205954
rect 153316 205718 153552 205954
rect 153636 205718 153872 205954
rect 153956 205718 154192 205954
rect 154276 205718 154512 205954
rect 154596 205718 154832 205954
rect 154916 205718 155152 205954
rect 155236 205718 155472 205954
rect 155556 205718 155792 205954
rect 155876 205718 156112 205954
rect 156196 205718 156432 205954
rect 156516 205718 156752 205954
rect 156836 205718 157072 205954
rect 157156 205718 157392 205954
rect 157476 205718 157712 205954
rect 157796 205718 158032 205954
rect 158116 205718 158352 205954
rect 158436 205718 158672 205954
rect 158756 205718 158992 205954
rect 159076 205718 159312 205954
rect 159396 205718 159632 205954
rect 159716 205718 159952 205954
rect 160036 205718 160272 205954
rect 160356 205718 160592 205954
rect 160676 205718 160912 205954
rect 160996 205718 161232 205954
rect 161316 205718 161552 205954
rect 161636 205718 161872 205954
rect 161956 205718 162192 205954
rect 162276 205718 162512 205954
rect 162596 205718 162832 205954
rect 162916 205718 163152 205954
rect 163236 205718 163472 205954
rect 163556 205718 163792 205954
rect 163876 205718 164112 205954
rect 164196 205718 164432 205954
rect 164516 205718 164752 205954
rect 164836 205718 165072 205954
rect 165156 205718 165392 205954
rect 136036 205398 136272 205634
rect 136356 205398 136592 205634
rect 136676 205398 136912 205634
rect 136996 205398 137232 205634
rect 137316 205398 137552 205634
rect 137636 205398 137872 205634
rect 137956 205398 138192 205634
rect 138276 205398 138512 205634
rect 138596 205398 138832 205634
rect 138916 205398 139152 205634
rect 139236 205398 139472 205634
rect 139556 205398 139792 205634
rect 139876 205398 140112 205634
rect 140196 205398 140432 205634
rect 140516 205398 140752 205634
rect 140836 205398 141072 205634
rect 141156 205398 141392 205634
rect 141476 205398 141712 205634
rect 141796 205398 142032 205634
rect 142116 205398 142352 205634
rect 142436 205398 142672 205634
rect 142756 205398 142992 205634
rect 143076 205398 143312 205634
rect 143396 205398 143632 205634
rect 143716 205398 143952 205634
rect 144036 205398 144272 205634
rect 144356 205398 144592 205634
rect 144676 205398 144912 205634
rect 144996 205398 145232 205634
rect 145316 205398 145552 205634
rect 145636 205398 145872 205634
rect 145956 205398 146192 205634
rect 146276 205398 146512 205634
rect 146596 205398 146832 205634
rect 146916 205398 147152 205634
rect 147236 205398 147472 205634
rect 147556 205398 147792 205634
rect 147876 205398 148112 205634
rect 148196 205398 148432 205634
rect 148516 205398 148752 205634
rect 148836 205398 149072 205634
rect 149156 205398 149392 205634
rect 149476 205398 149712 205634
rect 149796 205398 150032 205634
rect 150116 205398 150352 205634
rect 150436 205398 150672 205634
rect 150756 205398 150992 205634
rect 151076 205398 151312 205634
rect 151396 205398 151632 205634
rect 151716 205398 151952 205634
rect 152036 205398 152272 205634
rect 152356 205398 152592 205634
rect 152676 205398 152912 205634
rect 152996 205398 153232 205634
rect 153316 205398 153552 205634
rect 153636 205398 153872 205634
rect 153956 205398 154192 205634
rect 154276 205398 154512 205634
rect 154596 205398 154832 205634
rect 154916 205398 155152 205634
rect 155236 205398 155472 205634
rect 155556 205398 155792 205634
rect 155876 205398 156112 205634
rect 156196 205398 156432 205634
rect 156516 205398 156752 205634
rect 156836 205398 157072 205634
rect 157156 205398 157392 205634
rect 157476 205398 157712 205634
rect 157796 205398 158032 205634
rect 158116 205398 158352 205634
rect 158436 205398 158672 205634
rect 158756 205398 158992 205634
rect 159076 205398 159312 205634
rect 159396 205398 159632 205634
rect 159716 205398 159952 205634
rect 160036 205398 160272 205634
rect 160356 205398 160592 205634
rect 160676 205398 160912 205634
rect 160996 205398 161232 205634
rect 161316 205398 161552 205634
rect 161636 205398 161872 205634
rect 161956 205398 162192 205634
rect 162276 205398 162512 205634
rect 162596 205398 162832 205634
rect 162916 205398 163152 205634
rect 163236 205398 163472 205634
rect 163556 205398 163792 205634
rect 163876 205398 164112 205634
rect 164196 205398 164432 205634
rect 164516 205398 164752 205634
rect 164836 205398 165072 205634
rect 165156 205398 165392 205634
rect 168326 205718 168562 205954
rect 168646 205718 168882 205954
rect 168326 205398 168562 205634
rect 168646 205398 168882 205634
rect 137376 201218 137612 201454
rect 137696 201218 137932 201454
rect 138016 201218 138252 201454
rect 138336 201218 138572 201454
rect 138656 201218 138892 201454
rect 138976 201218 139212 201454
rect 139296 201218 139532 201454
rect 139616 201218 139852 201454
rect 139936 201218 140172 201454
rect 140256 201218 140492 201454
rect 140576 201218 140812 201454
rect 140896 201218 141132 201454
rect 141216 201218 141452 201454
rect 141536 201218 141772 201454
rect 141856 201218 142092 201454
rect 142176 201218 142412 201454
rect 142496 201218 142732 201454
rect 142816 201218 143052 201454
rect 143136 201218 143372 201454
rect 143456 201218 143692 201454
rect 143776 201218 144012 201454
rect 144096 201218 144332 201454
rect 144416 201218 144652 201454
rect 144736 201218 144972 201454
rect 145056 201218 145292 201454
rect 145376 201218 145612 201454
rect 145696 201218 145932 201454
rect 146016 201218 146252 201454
rect 146336 201218 146572 201454
rect 146656 201218 146892 201454
rect 146976 201218 147212 201454
rect 147296 201218 147532 201454
rect 147616 201218 147852 201454
rect 147936 201218 148172 201454
rect 148256 201218 148492 201454
rect 148576 201218 148812 201454
rect 148896 201218 149132 201454
rect 149216 201218 149452 201454
rect 149536 201218 149772 201454
rect 149856 201218 150092 201454
rect 150176 201218 150412 201454
rect 150496 201218 150732 201454
rect 150816 201218 151052 201454
rect 151136 201218 151372 201454
rect 151456 201218 151692 201454
rect 151776 201218 152012 201454
rect 152096 201218 152332 201454
rect 152416 201218 152652 201454
rect 152736 201218 152972 201454
rect 153056 201218 153292 201454
rect 153376 201218 153612 201454
rect 153696 201218 153932 201454
rect 154016 201218 154252 201454
rect 154336 201218 154572 201454
rect 154656 201218 154892 201454
rect 154976 201218 155212 201454
rect 155296 201218 155532 201454
rect 155616 201218 155852 201454
rect 155936 201218 156172 201454
rect 156256 201218 156492 201454
rect 156576 201218 156812 201454
rect 156896 201218 157132 201454
rect 157216 201218 157452 201454
rect 157536 201218 157772 201454
rect 157856 201218 158092 201454
rect 158176 201218 158412 201454
rect 158496 201218 158732 201454
rect 158816 201218 159052 201454
rect 159136 201218 159372 201454
rect 159456 201218 159692 201454
rect 159776 201218 160012 201454
rect 160096 201218 160332 201454
rect 160416 201218 160652 201454
rect 160736 201218 160972 201454
rect 161056 201218 161292 201454
rect 161376 201218 161612 201454
rect 161696 201218 161932 201454
rect 162016 201218 162252 201454
rect 162336 201218 162572 201454
rect 162656 201218 162892 201454
rect 162976 201218 163212 201454
rect 163296 201218 163532 201454
rect 163616 201218 163852 201454
rect 163936 201218 164172 201454
rect 164256 201218 164492 201454
rect 164576 201218 164812 201454
rect 164896 201218 165132 201454
rect 165216 201218 165452 201454
rect 137376 200898 137612 201134
rect 137696 200898 137932 201134
rect 138016 200898 138252 201134
rect 138336 200898 138572 201134
rect 138656 200898 138892 201134
rect 138976 200898 139212 201134
rect 139296 200898 139532 201134
rect 139616 200898 139852 201134
rect 139936 200898 140172 201134
rect 140256 200898 140492 201134
rect 140576 200898 140812 201134
rect 140896 200898 141132 201134
rect 141216 200898 141452 201134
rect 141536 200898 141772 201134
rect 141856 200898 142092 201134
rect 142176 200898 142412 201134
rect 142496 200898 142732 201134
rect 142816 200898 143052 201134
rect 143136 200898 143372 201134
rect 143456 200898 143692 201134
rect 143776 200898 144012 201134
rect 144096 200898 144332 201134
rect 144416 200898 144652 201134
rect 144736 200898 144972 201134
rect 145056 200898 145292 201134
rect 145376 200898 145612 201134
rect 145696 200898 145932 201134
rect 146016 200898 146252 201134
rect 146336 200898 146572 201134
rect 146656 200898 146892 201134
rect 146976 200898 147212 201134
rect 147296 200898 147532 201134
rect 147616 200898 147852 201134
rect 147936 200898 148172 201134
rect 148256 200898 148492 201134
rect 148576 200898 148812 201134
rect 148896 200898 149132 201134
rect 149216 200898 149452 201134
rect 149536 200898 149772 201134
rect 149856 200898 150092 201134
rect 150176 200898 150412 201134
rect 150496 200898 150732 201134
rect 150816 200898 151052 201134
rect 151136 200898 151372 201134
rect 151456 200898 151692 201134
rect 151776 200898 152012 201134
rect 152096 200898 152332 201134
rect 152416 200898 152652 201134
rect 152736 200898 152972 201134
rect 153056 200898 153292 201134
rect 153376 200898 153612 201134
rect 153696 200898 153932 201134
rect 154016 200898 154252 201134
rect 154336 200898 154572 201134
rect 154656 200898 154892 201134
rect 154976 200898 155212 201134
rect 155296 200898 155532 201134
rect 155616 200898 155852 201134
rect 155936 200898 156172 201134
rect 156256 200898 156492 201134
rect 156576 200898 156812 201134
rect 156896 200898 157132 201134
rect 157216 200898 157452 201134
rect 157536 200898 157772 201134
rect 157856 200898 158092 201134
rect 158176 200898 158412 201134
rect 158496 200898 158732 201134
rect 158816 200898 159052 201134
rect 159136 200898 159372 201134
rect 159456 200898 159692 201134
rect 159776 200898 160012 201134
rect 160096 200898 160332 201134
rect 160416 200898 160652 201134
rect 160736 200898 160972 201134
rect 161056 200898 161292 201134
rect 161376 200898 161612 201134
rect 161696 200898 161932 201134
rect 162016 200898 162252 201134
rect 162336 200898 162572 201134
rect 162656 200898 162892 201134
rect 162976 200898 163212 201134
rect 163296 200898 163532 201134
rect 163616 200898 163852 201134
rect 163936 200898 164172 201134
rect 164256 200898 164492 201134
rect 164576 200898 164812 201134
rect 164896 200898 165132 201134
rect 165216 200898 165452 201134
rect 132326 169718 132562 169954
rect 132646 169718 132882 169954
rect 132326 169398 132562 169634
rect 132646 169398 132882 169634
rect 168326 169718 168562 169954
rect 168646 169718 168882 169954
rect 168326 169398 168562 169634
rect 168646 169398 168882 169634
rect 172826 210218 173062 210454
rect 173146 210218 173382 210454
rect 172826 209898 173062 210134
rect 173146 209898 173382 210134
rect 172826 174218 173062 174454
rect 173146 174218 173382 174454
rect 172826 173898 173062 174134
rect 173146 173898 173382 174134
rect 177326 214718 177562 214954
rect 177646 214718 177882 214954
rect 177326 214398 177562 214634
rect 177646 214398 177882 214634
rect 177326 178718 177562 178954
rect 177646 178718 177882 178954
rect 177326 178398 177562 178634
rect 177646 178398 177882 178634
rect 177326 142718 177562 142954
rect 177646 142718 177882 142954
rect 177326 142398 177562 142634
rect 177646 142398 177882 142634
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 186326 223718 186562 223954
rect 186646 223718 186882 223954
rect 186326 223398 186562 223634
rect 186646 223398 186882 223634
rect 186326 187718 186562 187954
rect 186646 187718 186882 187954
rect 186326 187398 186562 187634
rect 186646 187398 186882 187634
rect 186326 151718 186562 151954
rect 186646 151718 186882 151954
rect 186326 151398 186562 151634
rect 186646 151398 186882 151634
rect 114326 115718 114562 115954
rect 114646 115718 114882 115954
rect 114326 115398 114562 115634
rect 114646 115398 114882 115634
rect 139610 115718 139846 115954
rect 139610 115398 139846 115634
rect 170330 115718 170566 115954
rect 170330 115398 170566 115634
rect 186326 115718 186562 115954
rect 186646 115718 186882 115954
rect 186326 115398 186562 115634
rect 186646 115398 186882 115634
rect 124250 111218 124486 111454
rect 124250 110898 124486 111134
rect 154970 111218 155206 111454
rect 154970 110898 155206 111134
rect 114326 79718 114562 79954
rect 114646 79718 114882 79954
rect 114326 79398 114562 79634
rect 114646 79398 114882 79634
rect 114326 43718 114562 43954
rect 114646 43718 114882 43954
rect 114326 43398 114562 43634
rect 114646 43398 114882 43634
rect 114326 7718 114562 7954
rect 114646 7718 114882 7954
rect 114326 7398 114562 7634
rect 114646 7398 114882 7634
rect 114326 -1542 114562 -1306
rect 114646 -1542 114882 -1306
rect 114326 -1862 114562 -1626
rect 114646 -1862 114882 -1626
rect 118826 48218 119062 48454
rect 119146 48218 119382 48454
rect 118826 47898 119062 48134
rect 119146 47898 119382 48134
rect 118826 12218 119062 12454
rect 119146 12218 119382 12454
rect 118826 11898 119062 12134
rect 119146 11898 119382 12134
rect 118826 -2502 119062 -2266
rect 119146 -2502 119382 -2266
rect 118826 -2822 119062 -2586
rect 119146 -2822 119382 -2586
rect 123326 52718 123562 52954
rect 123646 52718 123882 52954
rect 123326 52398 123562 52634
rect 123646 52398 123882 52634
rect 123326 16718 123562 16954
rect 123646 16718 123882 16954
rect 123326 16398 123562 16634
rect 123646 16398 123882 16634
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 123326 -3462 123562 -3226
rect 123646 -3462 123882 -3226
rect 123326 -3782 123562 -3546
rect 123646 -3782 123882 -3546
rect 132326 61718 132562 61954
rect 132646 61718 132882 61954
rect 132326 61398 132562 61634
rect 132646 61398 132882 61634
rect 132326 25718 132562 25954
rect 132646 25718 132882 25954
rect 132326 25398 132562 25634
rect 132646 25398 132882 25634
rect 127826 -4422 128062 -4186
rect 128146 -4422 128382 -4186
rect 127826 -4742 128062 -4506
rect 128146 -4742 128382 -4506
rect 136826 66218 137062 66454
rect 137146 66218 137382 66454
rect 136826 65898 137062 66134
rect 137146 65898 137382 66134
rect 136826 30218 137062 30454
rect 137146 30218 137382 30454
rect 136826 29898 137062 30134
rect 137146 29898 137382 30134
rect 132326 -5382 132562 -5146
rect 132646 -5382 132882 -5146
rect 132326 -5702 132562 -5466
rect 132646 -5702 132882 -5466
rect 141326 70718 141562 70954
rect 141646 70718 141882 70954
rect 141326 70398 141562 70634
rect 141646 70398 141882 70634
rect 141326 34718 141562 34954
rect 141646 34718 141882 34954
rect 141326 34398 141562 34634
rect 141646 34398 141882 34634
rect 136826 -6342 137062 -6106
rect 137146 -6342 137382 -6106
rect 136826 -6662 137062 -6426
rect 137146 -6662 137382 -6426
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 141326 -7302 141562 -7066
rect 141646 -7302 141882 -7066
rect 141326 -7622 141562 -7386
rect 141646 -7622 141882 -7386
rect 150326 43718 150562 43954
rect 150646 43718 150882 43954
rect 150326 43398 150562 43634
rect 150646 43398 150882 43634
rect 154826 48218 155062 48454
rect 155146 48218 155382 48454
rect 154826 47898 155062 48134
rect 155146 47898 155382 48134
rect 154826 12218 155062 12454
rect 155146 12218 155382 12454
rect 154826 11898 155062 12134
rect 155146 11898 155382 12134
rect 150326 7718 150562 7954
rect 150646 7718 150882 7954
rect 150326 7398 150562 7634
rect 150646 7398 150882 7634
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 150326 -1542 150562 -1306
rect 150646 -1542 150882 -1306
rect 150326 -1862 150562 -1626
rect 150646 -1862 150882 -1626
rect 159326 52718 159562 52954
rect 159646 52718 159882 52954
rect 159326 52398 159562 52634
rect 159646 52398 159882 52634
rect 159326 16718 159562 16954
rect 159646 16718 159882 16954
rect 159326 16398 159562 16634
rect 159646 16398 159882 16634
rect 154826 -2502 155062 -2266
rect 155146 -2502 155382 -2266
rect 154826 -2822 155062 -2586
rect 155146 -2822 155382 -2586
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 159326 -3462 159562 -3226
rect 159646 -3462 159882 -3226
rect 159326 -3782 159562 -3546
rect 159646 -3782 159882 -3546
rect 168326 61718 168562 61954
rect 168646 61718 168882 61954
rect 168326 61398 168562 61634
rect 168646 61398 168882 61634
rect 168326 25718 168562 25954
rect 168646 25718 168882 25954
rect 168326 25398 168562 25634
rect 168646 25398 168882 25634
rect 163826 -4422 164062 -4186
rect 164146 -4422 164382 -4186
rect 163826 -4742 164062 -4506
rect 164146 -4742 164382 -4506
rect 186326 79718 186562 79954
rect 186646 79718 186882 79954
rect 186326 79398 186562 79634
rect 186646 79398 186882 79634
rect 172826 66218 173062 66454
rect 173146 66218 173382 66454
rect 172826 65898 173062 66134
rect 173146 65898 173382 66134
rect 172826 30218 173062 30454
rect 173146 30218 173382 30454
rect 172826 29898 173062 30134
rect 173146 29898 173382 30134
rect 168326 -5382 168562 -5146
rect 168646 -5382 168882 -5146
rect 168326 -5702 168562 -5466
rect 168646 -5702 168882 -5466
rect 172826 -6342 173062 -6106
rect 173146 -6342 173382 -6106
rect 172826 -6662 173062 -6426
rect 173146 -6662 173382 -6426
rect 177326 70718 177562 70954
rect 177646 70718 177882 70954
rect 177326 70398 177562 70634
rect 177646 70398 177882 70634
rect 177326 34718 177562 34954
rect 177646 34718 177882 34954
rect 177326 34398 177562 34634
rect 177646 34398 177882 34634
rect 177326 -7302 177562 -7066
rect 177646 -7302 177882 -7066
rect 177326 -7622 177562 -7386
rect 177646 -7622 177882 -7386
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 186326 43718 186562 43954
rect 186646 43718 186882 43954
rect 186326 43398 186562 43634
rect 186646 43398 186882 43634
rect 186326 7718 186562 7954
rect 186646 7718 186882 7954
rect 186326 7398 186562 7634
rect 186646 7398 186882 7634
rect 186326 -1542 186562 -1306
rect 186646 -1542 186882 -1306
rect 186326 -1862 186562 -1626
rect 186646 -1862 186882 -1626
rect 190826 228217 191062 228453
rect 191146 228217 191382 228453
rect 190826 227897 191062 228133
rect 191146 227897 191382 228133
rect 190826 192218 191062 192454
rect 191146 192218 191382 192454
rect 190826 191898 191062 192134
rect 191146 191898 191382 192134
rect 190826 156218 191062 156454
rect 191146 156218 191382 156454
rect 190826 155898 191062 156134
rect 191146 155898 191382 156134
rect 190826 120218 191062 120454
rect 191146 120218 191382 120454
rect 190826 119898 191062 120134
rect 191146 119898 191382 120134
rect 190826 84218 191062 84454
rect 191146 84218 191382 84454
rect 190826 83898 191062 84134
rect 191146 83898 191382 84134
rect 190826 48218 191062 48454
rect 191146 48218 191382 48454
rect 190826 47898 191062 48134
rect 191146 47898 191382 48134
rect 190826 12218 191062 12454
rect 191146 12218 191382 12454
rect 190826 11898 191062 12134
rect 191146 11898 191382 12134
rect 190826 -2502 191062 -2266
rect 191146 -2502 191382 -2266
rect 190826 -2822 191062 -2586
rect 191146 -2822 191382 -2586
rect 195326 196718 195562 196954
rect 195646 196718 195882 196954
rect 195326 196398 195562 196634
rect 195646 196398 195882 196634
rect 195326 160718 195562 160954
rect 195646 160718 195882 160954
rect 195326 160398 195562 160634
rect 195646 160398 195882 160634
rect 195326 124718 195562 124954
rect 195646 124718 195882 124954
rect 195326 124398 195562 124634
rect 195646 124398 195882 124634
rect 195326 88718 195562 88954
rect 195646 88718 195882 88954
rect 195326 88398 195562 88634
rect 195646 88398 195882 88634
rect 195326 52718 195562 52954
rect 195646 52718 195882 52954
rect 195326 52398 195562 52634
rect 195646 52398 195882 52634
rect 195326 16718 195562 16954
rect 195646 16718 195882 16954
rect 195326 16398 195562 16634
rect 195646 16398 195882 16634
rect 195326 -3462 195562 -3226
rect 195646 -3462 195882 -3226
rect 195326 -3782 195562 -3546
rect 195646 -3782 195882 -3546
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -4422 200062 -4186
rect 200146 -4422 200382 -4186
rect 199826 -4742 200062 -4506
rect 200146 -4742 200382 -4506
rect 204326 205718 204562 205954
rect 204646 205718 204882 205954
rect 204326 205398 204562 205634
rect 204646 205398 204882 205634
rect 204326 169718 204562 169954
rect 204646 169718 204882 169954
rect 204326 169398 204562 169634
rect 204646 169398 204882 169634
rect 204326 133718 204562 133954
rect 204646 133718 204882 133954
rect 204326 133398 204562 133634
rect 204646 133398 204882 133634
rect 204326 97718 204562 97954
rect 204646 97718 204882 97954
rect 204326 97398 204562 97634
rect 204646 97398 204882 97634
rect 204326 61718 204562 61954
rect 204646 61718 204882 61954
rect 204326 61398 204562 61634
rect 204646 61398 204882 61634
rect 204326 25718 204562 25954
rect 204646 25718 204882 25954
rect 204326 25398 204562 25634
rect 204646 25398 204882 25634
rect 204326 -5382 204562 -5146
rect 204646 -5382 204882 -5146
rect 204326 -5702 204562 -5466
rect 204646 -5702 204882 -5466
rect 208826 210218 209062 210454
rect 209146 210218 209382 210454
rect 208826 209898 209062 210134
rect 209146 209898 209382 210134
rect 208826 174218 209062 174454
rect 209146 174218 209382 174454
rect 208826 173898 209062 174134
rect 209146 173898 209382 174134
rect 208826 138218 209062 138454
rect 209146 138218 209382 138454
rect 208826 137898 209062 138134
rect 209146 137898 209382 138134
rect 208826 102218 209062 102454
rect 209146 102218 209382 102454
rect 208826 101898 209062 102134
rect 209146 101898 209382 102134
rect 208826 66218 209062 66454
rect 209146 66218 209382 66454
rect 208826 65898 209062 66134
rect 209146 65898 209382 66134
rect 208826 30218 209062 30454
rect 209146 30218 209382 30454
rect 208826 29898 209062 30134
rect 209146 29898 209382 30134
rect 208826 -6342 209062 -6106
rect 209146 -6342 209382 -6106
rect 208826 -6662 209062 -6426
rect 209146 -6662 209382 -6426
rect 213326 214718 213562 214954
rect 213646 214718 213882 214954
rect 213326 214398 213562 214634
rect 213646 214398 213882 214634
rect 213326 178718 213562 178954
rect 213646 178718 213882 178954
rect 213326 178398 213562 178634
rect 213646 178398 213882 178634
rect 213326 142718 213562 142954
rect 213646 142718 213882 142954
rect 213326 142398 213562 142634
rect 213646 142398 213882 142634
rect 213326 106718 213562 106954
rect 213646 106718 213882 106954
rect 213326 106398 213562 106634
rect 213646 106398 213882 106634
rect 213326 70718 213562 70954
rect 213646 70718 213882 70954
rect 213326 70398 213562 70634
rect 213646 70398 213882 70634
rect 213326 34718 213562 34954
rect 213646 34718 213882 34954
rect 213326 34398 213562 34634
rect 213646 34398 213882 34634
rect 213326 -7302 213562 -7066
rect 213646 -7302 213882 -7066
rect 213326 -7622 213562 -7386
rect 213646 -7622 213882 -7386
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 222326 223718 222562 223954
rect 222646 223718 222882 223954
rect 222326 223398 222562 223634
rect 222646 223398 222882 223634
rect 222326 187718 222562 187954
rect 222646 187718 222882 187954
rect 222326 187398 222562 187634
rect 222646 187398 222882 187634
rect 222326 151718 222562 151954
rect 222646 151718 222882 151954
rect 222326 151398 222562 151634
rect 222646 151398 222882 151634
rect 222326 115718 222562 115954
rect 222646 115718 222882 115954
rect 222326 115398 222562 115634
rect 222646 115398 222882 115634
rect 222326 79718 222562 79954
rect 222646 79718 222882 79954
rect 222326 79398 222562 79634
rect 222646 79398 222882 79634
rect 222326 43718 222562 43954
rect 222646 43718 222882 43954
rect 222326 43398 222562 43634
rect 222646 43398 222882 43634
rect 222326 7718 222562 7954
rect 222646 7718 222882 7954
rect 222326 7398 222562 7634
rect 222646 7398 222882 7634
rect 222326 -1542 222562 -1306
rect 222646 -1542 222882 -1306
rect 222326 -1862 222562 -1626
rect 222646 -1862 222882 -1626
rect 226826 228217 227062 228453
rect 227146 228217 227382 228453
rect 226826 227897 227062 228133
rect 227146 227897 227382 228133
rect 226826 192218 227062 192454
rect 227146 192218 227382 192454
rect 226826 191898 227062 192134
rect 227146 191898 227382 192134
rect 226826 156218 227062 156454
rect 227146 156218 227382 156454
rect 226826 155898 227062 156134
rect 227146 155898 227382 156134
rect 226826 120218 227062 120454
rect 227146 120218 227382 120454
rect 226826 119898 227062 120134
rect 227146 119898 227382 120134
rect 226826 84218 227062 84454
rect 227146 84218 227382 84454
rect 226826 83898 227062 84134
rect 227146 83898 227382 84134
rect 226826 48218 227062 48454
rect 227146 48218 227382 48454
rect 226826 47898 227062 48134
rect 227146 47898 227382 48134
rect 226826 12218 227062 12454
rect 227146 12218 227382 12454
rect 226826 11898 227062 12134
rect 227146 11898 227382 12134
rect 226826 -2502 227062 -2266
rect 227146 -2502 227382 -2266
rect 226826 -2822 227062 -2586
rect 227146 -2822 227382 -2586
rect 231326 196718 231562 196954
rect 231646 196718 231882 196954
rect 231326 196398 231562 196634
rect 231646 196398 231882 196634
rect 231326 160718 231562 160954
rect 231646 160718 231882 160954
rect 231326 160398 231562 160634
rect 231646 160398 231882 160634
rect 231326 124718 231562 124954
rect 231646 124718 231882 124954
rect 231326 124398 231562 124634
rect 231646 124398 231882 124634
rect 231326 88718 231562 88954
rect 231646 88718 231882 88954
rect 231326 88398 231562 88634
rect 231646 88398 231882 88634
rect 231326 52718 231562 52954
rect 231646 52718 231882 52954
rect 231326 52398 231562 52634
rect 231646 52398 231882 52634
rect 231326 16718 231562 16954
rect 231646 16718 231882 16954
rect 231326 16398 231562 16634
rect 231646 16398 231882 16634
rect 231326 -3462 231562 -3226
rect 231646 -3462 231882 -3226
rect 231326 -3782 231562 -3546
rect 231646 -3782 231882 -3546
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -4422 236062 -4186
rect 236146 -4422 236382 -4186
rect 235826 -4742 236062 -4506
rect 236146 -4742 236382 -4506
rect 240326 205718 240562 205954
rect 240646 205718 240882 205954
rect 240326 205398 240562 205634
rect 240646 205398 240882 205634
rect 240326 169718 240562 169954
rect 240646 169718 240882 169954
rect 240326 169398 240562 169634
rect 240646 169398 240882 169634
rect 240326 133718 240562 133954
rect 240646 133718 240882 133954
rect 240326 133398 240562 133634
rect 240646 133398 240882 133634
rect 240326 97718 240562 97954
rect 240646 97718 240882 97954
rect 240326 97398 240562 97634
rect 240646 97398 240882 97634
rect 240326 61718 240562 61954
rect 240646 61718 240882 61954
rect 240326 61398 240562 61634
rect 240646 61398 240882 61634
rect 240326 25718 240562 25954
rect 240646 25718 240882 25954
rect 240326 25398 240562 25634
rect 240646 25398 240882 25634
rect 240326 -5382 240562 -5146
rect 240646 -5382 240882 -5146
rect 240326 -5702 240562 -5466
rect 240646 -5702 240882 -5466
rect 244826 210218 245062 210454
rect 245146 210218 245382 210454
rect 244826 209898 245062 210134
rect 245146 209898 245382 210134
rect 244826 174218 245062 174454
rect 245146 174218 245382 174454
rect 244826 173898 245062 174134
rect 245146 173898 245382 174134
rect 244826 138218 245062 138454
rect 245146 138218 245382 138454
rect 244826 137898 245062 138134
rect 245146 137898 245382 138134
rect 244826 102218 245062 102454
rect 245146 102218 245382 102454
rect 244826 101898 245062 102134
rect 245146 101898 245382 102134
rect 244826 66218 245062 66454
rect 245146 66218 245382 66454
rect 244826 65898 245062 66134
rect 245146 65898 245382 66134
rect 244826 30218 245062 30454
rect 245146 30218 245382 30454
rect 244826 29898 245062 30134
rect 245146 29898 245382 30134
rect 244826 -6342 245062 -6106
rect 245146 -6342 245382 -6106
rect 244826 -6662 245062 -6426
rect 245146 -6662 245382 -6426
rect 249326 214718 249562 214954
rect 249646 214718 249882 214954
rect 249326 214398 249562 214634
rect 249646 214398 249882 214634
rect 249326 178718 249562 178954
rect 249646 178718 249882 178954
rect 249326 178398 249562 178634
rect 249646 178398 249882 178634
rect 249326 142718 249562 142954
rect 249646 142718 249882 142954
rect 249326 142398 249562 142634
rect 249646 142398 249882 142634
rect 249326 106718 249562 106954
rect 249646 106718 249882 106954
rect 249326 106398 249562 106634
rect 249646 106398 249882 106634
rect 249326 70718 249562 70954
rect 249646 70718 249882 70954
rect 249326 70398 249562 70634
rect 249646 70398 249882 70634
rect 249326 34718 249562 34954
rect 249646 34718 249882 34954
rect 249326 34398 249562 34634
rect 249646 34398 249882 34634
rect 249326 -7302 249562 -7066
rect 249646 -7302 249882 -7066
rect 249326 -7622 249562 -7386
rect 249646 -7622 249882 -7386
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 258326 223718 258562 223954
rect 258646 223718 258882 223954
rect 258326 223398 258562 223634
rect 258646 223398 258882 223634
rect 258326 187718 258562 187954
rect 258646 187718 258882 187954
rect 258326 187398 258562 187634
rect 258646 187398 258882 187634
rect 258326 151718 258562 151954
rect 258646 151718 258882 151954
rect 258326 151398 258562 151634
rect 258646 151398 258882 151634
rect 258326 115718 258562 115954
rect 258646 115718 258882 115954
rect 258326 115398 258562 115634
rect 258646 115398 258882 115634
rect 258326 79718 258562 79954
rect 258646 79718 258882 79954
rect 258326 79398 258562 79634
rect 258646 79398 258882 79634
rect 258326 43718 258562 43954
rect 258646 43718 258882 43954
rect 258326 43398 258562 43634
rect 258646 43398 258882 43634
rect 258326 7718 258562 7954
rect 258646 7718 258882 7954
rect 258326 7398 258562 7634
rect 258646 7398 258882 7634
rect 258326 -1542 258562 -1306
rect 258646 -1542 258882 -1306
rect 258326 -1862 258562 -1626
rect 258646 -1862 258882 -1626
rect 262826 228217 263062 228453
rect 263146 228217 263382 228453
rect 262826 227897 263062 228133
rect 263146 227897 263382 228133
rect 262826 192218 263062 192454
rect 263146 192218 263382 192454
rect 262826 191898 263062 192134
rect 263146 191898 263382 192134
rect 262826 156218 263062 156454
rect 263146 156218 263382 156454
rect 262826 155898 263062 156134
rect 263146 155898 263382 156134
rect 262826 120218 263062 120454
rect 263146 120218 263382 120454
rect 262826 119898 263062 120134
rect 263146 119898 263382 120134
rect 262826 84218 263062 84454
rect 263146 84218 263382 84454
rect 262826 83898 263062 84134
rect 263146 83898 263382 84134
rect 262826 48218 263062 48454
rect 263146 48218 263382 48454
rect 262826 47898 263062 48134
rect 263146 47898 263382 48134
rect 262826 12218 263062 12454
rect 263146 12218 263382 12454
rect 262826 11898 263062 12134
rect 263146 11898 263382 12134
rect 262826 -2502 263062 -2266
rect 263146 -2502 263382 -2266
rect 262826 -2822 263062 -2586
rect 263146 -2822 263382 -2586
rect 267326 196718 267562 196954
rect 267646 196718 267882 196954
rect 267326 196398 267562 196634
rect 267646 196398 267882 196634
rect 267326 160718 267562 160954
rect 267646 160718 267882 160954
rect 267326 160398 267562 160634
rect 267646 160398 267882 160634
rect 267326 124718 267562 124954
rect 267646 124718 267882 124954
rect 267326 124398 267562 124634
rect 267646 124398 267882 124634
rect 267326 88718 267562 88954
rect 267646 88718 267882 88954
rect 267326 88398 267562 88634
rect 267646 88398 267882 88634
rect 267326 52718 267562 52954
rect 267646 52718 267882 52954
rect 267326 52398 267562 52634
rect 267646 52398 267882 52634
rect 267326 16718 267562 16954
rect 267646 16718 267882 16954
rect 267326 16398 267562 16634
rect 267646 16398 267882 16634
rect 267326 -3462 267562 -3226
rect 267646 -3462 267882 -3226
rect 267326 -3782 267562 -3546
rect 267646 -3782 267882 -3546
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -4422 272062 -4186
rect 272146 -4422 272382 -4186
rect 271826 -4742 272062 -4506
rect 272146 -4742 272382 -4506
rect 276326 205718 276562 205954
rect 276646 205718 276882 205954
rect 276326 205398 276562 205634
rect 276646 205398 276882 205634
rect 276326 169718 276562 169954
rect 276646 169718 276882 169954
rect 276326 169398 276562 169634
rect 276646 169398 276882 169634
rect 276326 133718 276562 133954
rect 276646 133718 276882 133954
rect 276326 133398 276562 133634
rect 276646 133398 276882 133634
rect 276326 97718 276562 97954
rect 276646 97718 276882 97954
rect 276326 97398 276562 97634
rect 276646 97398 276882 97634
rect 276326 61718 276562 61954
rect 276646 61718 276882 61954
rect 276326 61398 276562 61634
rect 276646 61398 276882 61634
rect 276326 25718 276562 25954
rect 276646 25718 276882 25954
rect 276326 25398 276562 25634
rect 276646 25398 276882 25634
rect 276326 -5382 276562 -5146
rect 276646 -5382 276882 -5146
rect 276326 -5702 276562 -5466
rect 276646 -5702 276882 -5466
rect 280826 210218 281062 210454
rect 281146 210218 281382 210454
rect 280826 209898 281062 210134
rect 281146 209898 281382 210134
rect 280826 174218 281062 174454
rect 281146 174218 281382 174454
rect 280826 173898 281062 174134
rect 281146 173898 281382 174134
rect 280826 138218 281062 138454
rect 281146 138218 281382 138454
rect 280826 137898 281062 138134
rect 281146 137898 281382 138134
rect 280826 102218 281062 102454
rect 281146 102218 281382 102454
rect 280826 101898 281062 102134
rect 281146 101898 281382 102134
rect 280826 66218 281062 66454
rect 281146 66218 281382 66454
rect 280826 65898 281062 66134
rect 281146 65898 281382 66134
rect 280826 30218 281062 30454
rect 281146 30218 281382 30454
rect 280826 29898 281062 30134
rect 281146 29898 281382 30134
rect 280826 -6342 281062 -6106
rect 281146 -6342 281382 -6106
rect 280826 -6662 281062 -6426
rect 281146 -6662 281382 -6426
rect 285326 214718 285562 214954
rect 285646 214718 285882 214954
rect 285326 214398 285562 214634
rect 285646 214398 285882 214634
rect 285326 178718 285562 178954
rect 285646 178718 285882 178954
rect 285326 178398 285562 178634
rect 285646 178398 285882 178634
rect 285326 142718 285562 142954
rect 285646 142718 285882 142954
rect 285326 142398 285562 142634
rect 285646 142398 285882 142634
rect 285326 106718 285562 106954
rect 285646 106718 285882 106954
rect 285326 106398 285562 106634
rect 285646 106398 285882 106634
rect 285326 70718 285562 70954
rect 285646 70718 285882 70954
rect 285326 70398 285562 70634
rect 285646 70398 285882 70634
rect 285326 34718 285562 34954
rect 285646 34718 285882 34954
rect 285326 34398 285562 34634
rect 285646 34398 285882 34634
rect 285326 -7302 285562 -7066
rect 285646 -7302 285882 -7066
rect 285326 -7622 285562 -7386
rect 285646 -7622 285882 -7386
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 294326 223718 294562 223954
rect 294646 223718 294882 223954
rect 294326 223398 294562 223634
rect 294646 223398 294882 223634
rect 294326 187718 294562 187954
rect 294646 187718 294882 187954
rect 294326 187398 294562 187634
rect 294646 187398 294882 187634
rect 294326 151718 294562 151954
rect 294646 151718 294882 151954
rect 294326 151398 294562 151634
rect 294646 151398 294882 151634
rect 294326 115718 294562 115954
rect 294646 115718 294882 115954
rect 294326 115398 294562 115634
rect 294646 115398 294882 115634
rect 294326 79718 294562 79954
rect 294646 79718 294882 79954
rect 294326 79398 294562 79634
rect 294646 79398 294882 79634
rect 294326 43718 294562 43954
rect 294646 43718 294882 43954
rect 294326 43398 294562 43634
rect 294646 43398 294882 43634
rect 294326 7718 294562 7954
rect 294646 7718 294882 7954
rect 294326 7398 294562 7634
rect 294646 7398 294882 7634
rect 294326 -1542 294562 -1306
rect 294646 -1542 294882 -1306
rect 294326 -1862 294562 -1626
rect 294646 -1862 294882 -1626
rect 298826 228217 299062 228453
rect 299146 228217 299382 228453
rect 298826 227897 299062 228133
rect 299146 227897 299382 228133
rect 298826 192218 299062 192454
rect 299146 192218 299382 192454
rect 298826 191898 299062 192134
rect 299146 191898 299382 192134
rect 298826 156218 299062 156454
rect 299146 156218 299382 156454
rect 298826 155898 299062 156134
rect 299146 155898 299382 156134
rect 298826 120218 299062 120454
rect 299146 120218 299382 120454
rect 298826 119898 299062 120134
rect 299146 119898 299382 120134
rect 298826 84218 299062 84454
rect 299146 84218 299382 84454
rect 298826 83898 299062 84134
rect 299146 83898 299382 84134
rect 298826 48218 299062 48454
rect 299146 48218 299382 48454
rect 298826 47898 299062 48134
rect 299146 47898 299382 48134
rect 298826 12218 299062 12454
rect 299146 12218 299382 12454
rect 298826 11898 299062 12134
rect 299146 11898 299382 12134
rect 298826 -2502 299062 -2266
rect 299146 -2502 299382 -2266
rect 298826 -2822 299062 -2586
rect 299146 -2822 299382 -2586
rect 303326 196718 303562 196954
rect 303646 196718 303882 196954
rect 303326 196398 303562 196634
rect 303646 196398 303882 196634
rect 303326 160718 303562 160954
rect 303646 160718 303882 160954
rect 303326 160398 303562 160634
rect 303646 160398 303882 160634
rect 303326 124718 303562 124954
rect 303646 124718 303882 124954
rect 303326 124398 303562 124634
rect 303646 124398 303882 124634
rect 303326 88718 303562 88954
rect 303646 88718 303882 88954
rect 303326 88398 303562 88634
rect 303646 88398 303882 88634
rect 303326 52718 303562 52954
rect 303646 52718 303882 52954
rect 303326 52398 303562 52634
rect 303646 52398 303882 52634
rect 303326 16718 303562 16954
rect 303646 16718 303882 16954
rect 303326 16398 303562 16634
rect 303646 16398 303882 16634
rect 303326 -3462 303562 -3226
rect 303646 -3462 303882 -3226
rect 303326 -3782 303562 -3546
rect 303646 -3782 303882 -3546
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -4422 308062 -4186
rect 308146 -4422 308382 -4186
rect 307826 -4742 308062 -4506
rect 308146 -4742 308382 -4506
rect 312326 205718 312562 205954
rect 312646 205718 312882 205954
rect 312326 205398 312562 205634
rect 312646 205398 312882 205634
rect 312326 169718 312562 169954
rect 312646 169718 312882 169954
rect 312326 169398 312562 169634
rect 312646 169398 312882 169634
rect 312326 133718 312562 133954
rect 312646 133718 312882 133954
rect 312326 133398 312562 133634
rect 312646 133398 312882 133634
rect 312326 97718 312562 97954
rect 312646 97718 312882 97954
rect 312326 97398 312562 97634
rect 312646 97398 312882 97634
rect 312326 61718 312562 61954
rect 312646 61718 312882 61954
rect 312326 61398 312562 61634
rect 312646 61398 312882 61634
rect 312326 25718 312562 25954
rect 312646 25718 312882 25954
rect 312326 25398 312562 25634
rect 312646 25398 312882 25634
rect 312326 -5382 312562 -5146
rect 312646 -5382 312882 -5146
rect 312326 -5702 312562 -5466
rect 312646 -5702 312882 -5466
rect 316826 210218 317062 210454
rect 317146 210218 317382 210454
rect 316826 209898 317062 210134
rect 317146 209898 317382 210134
rect 316826 174218 317062 174454
rect 317146 174218 317382 174454
rect 316826 173898 317062 174134
rect 317146 173898 317382 174134
rect 316826 138218 317062 138454
rect 317146 138218 317382 138454
rect 316826 137898 317062 138134
rect 317146 137898 317382 138134
rect 316826 102218 317062 102454
rect 317146 102218 317382 102454
rect 316826 101898 317062 102134
rect 317146 101898 317382 102134
rect 316826 66218 317062 66454
rect 317146 66218 317382 66454
rect 316826 65898 317062 66134
rect 317146 65898 317382 66134
rect 316826 30218 317062 30454
rect 317146 30218 317382 30454
rect 316826 29898 317062 30134
rect 317146 29898 317382 30134
rect 316826 -6342 317062 -6106
rect 317146 -6342 317382 -6106
rect 316826 -6662 317062 -6426
rect 317146 -6662 317382 -6426
rect 321326 214718 321562 214954
rect 321646 214718 321882 214954
rect 321326 214398 321562 214634
rect 321646 214398 321882 214634
rect 321326 178718 321562 178954
rect 321646 178718 321882 178954
rect 321326 178398 321562 178634
rect 321646 178398 321882 178634
rect 321326 142718 321562 142954
rect 321646 142718 321882 142954
rect 321326 142398 321562 142634
rect 321646 142398 321882 142634
rect 321326 106718 321562 106954
rect 321646 106718 321882 106954
rect 321326 106398 321562 106634
rect 321646 106398 321882 106634
rect 321326 70718 321562 70954
rect 321646 70718 321882 70954
rect 321326 70398 321562 70634
rect 321646 70398 321882 70634
rect 321326 34718 321562 34954
rect 321646 34718 321882 34954
rect 321326 34398 321562 34634
rect 321646 34398 321882 34634
rect 321326 -7302 321562 -7066
rect 321646 -7302 321882 -7066
rect 321326 -7622 321562 -7386
rect 321646 -7622 321882 -7386
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 330326 223718 330562 223954
rect 330646 223718 330882 223954
rect 330326 223398 330562 223634
rect 330646 223398 330882 223634
rect 330326 187718 330562 187954
rect 330646 187718 330882 187954
rect 330326 187398 330562 187634
rect 330646 187398 330882 187634
rect 330326 151718 330562 151954
rect 330646 151718 330882 151954
rect 330326 151398 330562 151634
rect 330646 151398 330882 151634
rect 330326 115718 330562 115954
rect 330646 115718 330882 115954
rect 330326 115398 330562 115634
rect 330646 115398 330882 115634
rect 330326 79718 330562 79954
rect 330646 79718 330882 79954
rect 330326 79398 330562 79634
rect 330646 79398 330882 79634
rect 330326 43718 330562 43954
rect 330646 43718 330882 43954
rect 330326 43398 330562 43634
rect 330646 43398 330882 43634
rect 330326 7718 330562 7954
rect 330646 7718 330882 7954
rect 330326 7398 330562 7634
rect 330646 7398 330882 7634
rect 330326 -1542 330562 -1306
rect 330646 -1542 330882 -1306
rect 330326 -1862 330562 -1626
rect 330646 -1862 330882 -1626
rect 334826 228217 335062 228453
rect 335146 228217 335382 228453
rect 334826 227897 335062 228133
rect 335146 227897 335382 228133
rect 334826 192218 335062 192454
rect 335146 192218 335382 192454
rect 334826 191898 335062 192134
rect 335146 191898 335382 192134
rect 334826 156218 335062 156454
rect 335146 156218 335382 156454
rect 334826 155898 335062 156134
rect 335146 155898 335382 156134
rect 334826 120218 335062 120454
rect 335146 120218 335382 120454
rect 334826 119898 335062 120134
rect 335146 119898 335382 120134
rect 334826 84218 335062 84454
rect 335146 84218 335382 84454
rect 334826 83898 335062 84134
rect 335146 83898 335382 84134
rect 334826 48218 335062 48454
rect 335146 48218 335382 48454
rect 334826 47898 335062 48134
rect 335146 47898 335382 48134
rect 334826 12218 335062 12454
rect 335146 12218 335382 12454
rect 334826 11898 335062 12134
rect 335146 11898 335382 12134
rect 334826 -2502 335062 -2266
rect 335146 -2502 335382 -2266
rect 334826 -2822 335062 -2586
rect 335146 -2822 335382 -2586
rect 339326 196718 339562 196954
rect 339646 196718 339882 196954
rect 339326 196398 339562 196634
rect 339646 196398 339882 196634
rect 339326 160718 339562 160954
rect 339646 160718 339882 160954
rect 339326 160398 339562 160634
rect 339646 160398 339882 160634
rect 339326 124718 339562 124954
rect 339646 124718 339882 124954
rect 339326 124398 339562 124634
rect 339646 124398 339882 124634
rect 339326 88718 339562 88954
rect 339646 88718 339882 88954
rect 339326 88398 339562 88634
rect 339646 88398 339882 88634
rect 339326 52718 339562 52954
rect 339646 52718 339882 52954
rect 339326 52398 339562 52634
rect 339646 52398 339882 52634
rect 339326 16718 339562 16954
rect 339646 16718 339882 16954
rect 339326 16398 339562 16634
rect 339646 16398 339882 16634
rect 339326 -3462 339562 -3226
rect 339646 -3462 339882 -3226
rect 339326 -3782 339562 -3546
rect 339646 -3782 339882 -3546
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -4422 344062 -4186
rect 344146 -4422 344382 -4186
rect 343826 -4742 344062 -4506
rect 344146 -4742 344382 -4506
rect 348326 205718 348562 205954
rect 348646 205718 348882 205954
rect 348326 205398 348562 205634
rect 348646 205398 348882 205634
rect 348326 169718 348562 169954
rect 348646 169718 348882 169954
rect 348326 169398 348562 169634
rect 348646 169398 348882 169634
rect 348326 133718 348562 133954
rect 348646 133718 348882 133954
rect 348326 133398 348562 133634
rect 348646 133398 348882 133634
rect 348326 97718 348562 97954
rect 348646 97718 348882 97954
rect 348326 97398 348562 97634
rect 348646 97398 348882 97634
rect 348326 61718 348562 61954
rect 348646 61718 348882 61954
rect 348326 61398 348562 61634
rect 348646 61398 348882 61634
rect 348326 25718 348562 25954
rect 348646 25718 348882 25954
rect 348326 25398 348562 25634
rect 348646 25398 348882 25634
rect 348326 -5382 348562 -5146
rect 348646 -5382 348882 -5146
rect 348326 -5702 348562 -5466
rect 348646 -5702 348882 -5466
rect 352826 210218 353062 210454
rect 353146 210218 353382 210454
rect 352826 209898 353062 210134
rect 353146 209898 353382 210134
rect 352826 174218 353062 174454
rect 353146 174218 353382 174454
rect 352826 173898 353062 174134
rect 353146 173898 353382 174134
rect 352826 138218 353062 138454
rect 353146 138218 353382 138454
rect 352826 137898 353062 138134
rect 353146 137898 353382 138134
rect 352826 102218 353062 102454
rect 353146 102218 353382 102454
rect 352826 101898 353062 102134
rect 353146 101898 353382 102134
rect 352826 66218 353062 66454
rect 353146 66218 353382 66454
rect 352826 65898 353062 66134
rect 353146 65898 353382 66134
rect 352826 30218 353062 30454
rect 353146 30218 353382 30454
rect 352826 29898 353062 30134
rect 353146 29898 353382 30134
rect 352826 -6342 353062 -6106
rect 353146 -6342 353382 -6106
rect 352826 -6662 353062 -6426
rect 353146 -6662 353382 -6426
rect 357326 214718 357562 214954
rect 357646 214718 357882 214954
rect 357326 214398 357562 214634
rect 357646 214398 357882 214634
rect 357326 178718 357562 178954
rect 357646 178718 357882 178954
rect 357326 178398 357562 178634
rect 357646 178398 357882 178634
rect 357326 142718 357562 142954
rect 357646 142718 357882 142954
rect 357326 142398 357562 142634
rect 357646 142398 357882 142634
rect 357326 106718 357562 106954
rect 357646 106718 357882 106954
rect 357326 106398 357562 106634
rect 357646 106398 357882 106634
rect 357326 70718 357562 70954
rect 357646 70718 357882 70954
rect 357326 70398 357562 70634
rect 357646 70398 357882 70634
rect 357326 34718 357562 34954
rect 357646 34718 357882 34954
rect 357326 34398 357562 34634
rect 357646 34398 357882 34634
rect 357326 -7302 357562 -7066
rect 357646 -7302 357882 -7066
rect 357326 -7622 357562 -7386
rect 357646 -7622 357882 -7386
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 366326 223718 366562 223954
rect 366646 223718 366882 223954
rect 366326 223398 366562 223634
rect 366646 223398 366882 223634
rect 366326 187718 366562 187954
rect 366646 187718 366882 187954
rect 366326 187398 366562 187634
rect 366646 187398 366882 187634
rect 366326 151718 366562 151954
rect 366646 151718 366882 151954
rect 366326 151398 366562 151634
rect 366646 151398 366882 151634
rect 366326 115718 366562 115954
rect 366646 115718 366882 115954
rect 366326 115398 366562 115634
rect 366646 115398 366882 115634
rect 366326 79718 366562 79954
rect 366646 79718 366882 79954
rect 366326 79398 366562 79634
rect 366646 79398 366882 79634
rect 366326 43718 366562 43954
rect 366646 43718 366882 43954
rect 366326 43398 366562 43634
rect 366646 43398 366882 43634
rect 366326 7718 366562 7954
rect 366646 7718 366882 7954
rect 366326 7398 366562 7634
rect 366646 7398 366882 7634
rect 366326 -1542 366562 -1306
rect 366646 -1542 366882 -1306
rect 366326 -1862 366562 -1626
rect 366646 -1862 366882 -1626
rect 370826 228217 371062 228453
rect 371146 228217 371382 228453
rect 370826 227897 371062 228133
rect 371146 227897 371382 228133
rect 370826 192218 371062 192454
rect 371146 192218 371382 192454
rect 370826 191898 371062 192134
rect 371146 191898 371382 192134
rect 370826 156218 371062 156454
rect 371146 156218 371382 156454
rect 370826 155898 371062 156134
rect 371146 155898 371382 156134
rect 370826 120218 371062 120454
rect 371146 120218 371382 120454
rect 370826 119898 371062 120134
rect 371146 119898 371382 120134
rect 370826 84218 371062 84454
rect 371146 84218 371382 84454
rect 370826 83898 371062 84134
rect 371146 83898 371382 84134
rect 370826 48218 371062 48454
rect 371146 48218 371382 48454
rect 370826 47898 371062 48134
rect 371146 47898 371382 48134
rect 370826 12218 371062 12454
rect 371146 12218 371382 12454
rect 370826 11898 371062 12134
rect 371146 11898 371382 12134
rect 370826 -2502 371062 -2266
rect 371146 -2502 371382 -2266
rect 370826 -2822 371062 -2586
rect 371146 -2822 371382 -2586
rect 375326 196718 375562 196954
rect 375646 196718 375882 196954
rect 375326 196398 375562 196634
rect 375646 196398 375882 196634
rect 375326 160718 375562 160954
rect 375646 160718 375882 160954
rect 375326 160398 375562 160634
rect 375646 160398 375882 160634
rect 375326 124718 375562 124954
rect 375646 124718 375882 124954
rect 375326 124398 375562 124634
rect 375646 124398 375882 124634
rect 375326 88718 375562 88954
rect 375646 88718 375882 88954
rect 375326 88398 375562 88634
rect 375646 88398 375882 88634
rect 375326 52718 375562 52954
rect 375646 52718 375882 52954
rect 375326 52398 375562 52634
rect 375646 52398 375882 52634
rect 375326 16718 375562 16954
rect 375646 16718 375882 16954
rect 375326 16398 375562 16634
rect 375646 16398 375882 16634
rect 375326 -3462 375562 -3226
rect 375646 -3462 375882 -3226
rect 375326 -3782 375562 -3546
rect 375646 -3782 375882 -3546
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -4422 380062 -4186
rect 380146 -4422 380382 -4186
rect 379826 -4742 380062 -4506
rect 380146 -4742 380382 -4506
rect 384326 205718 384562 205954
rect 384646 205718 384882 205954
rect 384326 205398 384562 205634
rect 384646 205398 384882 205634
rect 384326 169718 384562 169954
rect 384646 169718 384882 169954
rect 384326 169398 384562 169634
rect 384646 169398 384882 169634
rect 384326 133718 384562 133954
rect 384646 133718 384882 133954
rect 384326 133398 384562 133634
rect 384646 133398 384882 133634
rect 384326 97718 384562 97954
rect 384646 97718 384882 97954
rect 384326 97398 384562 97634
rect 384646 97398 384882 97634
rect 384326 61718 384562 61954
rect 384646 61718 384882 61954
rect 384326 61398 384562 61634
rect 384646 61398 384882 61634
rect 384326 25718 384562 25954
rect 384646 25718 384882 25954
rect 384326 25398 384562 25634
rect 384646 25398 384882 25634
rect 384326 -5382 384562 -5146
rect 384646 -5382 384882 -5146
rect 384326 -5702 384562 -5466
rect 384646 -5702 384882 -5466
rect 388826 210218 389062 210454
rect 389146 210218 389382 210454
rect 388826 209898 389062 210134
rect 389146 209898 389382 210134
rect 388826 174218 389062 174454
rect 389146 174218 389382 174454
rect 388826 173898 389062 174134
rect 389146 173898 389382 174134
rect 388826 138218 389062 138454
rect 389146 138218 389382 138454
rect 388826 137898 389062 138134
rect 389146 137898 389382 138134
rect 388826 102218 389062 102454
rect 389146 102218 389382 102454
rect 388826 101898 389062 102134
rect 389146 101898 389382 102134
rect 388826 66218 389062 66454
rect 389146 66218 389382 66454
rect 388826 65898 389062 66134
rect 389146 65898 389382 66134
rect 388826 30218 389062 30454
rect 389146 30218 389382 30454
rect 388826 29898 389062 30134
rect 389146 29898 389382 30134
rect 388826 -6342 389062 -6106
rect 389146 -6342 389382 -6106
rect 388826 -6662 389062 -6426
rect 389146 -6662 389382 -6426
rect 393326 214718 393562 214954
rect 393646 214718 393882 214954
rect 393326 214398 393562 214634
rect 393646 214398 393882 214634
rect 393326 178718 393562 178954
rect 393646 178718 393882 178954
rect 393326 178398 393562 178634
rect 393646 178398 393882 178634
rect 393326 142718 393562 142954
rect 393646 142718 393882 142954
rect 393326 142398 393562 142634
rect 393646 142398 393882 142634
rect 393326 106718 393562 106954
rect 393646 106718 393882 106954
rect 393326 106398 393562 106634
rect 393646 106398 393882 106634
rect 393326 70718 393562 70954
rect 393646 70718 393882 70954
rect 393326 70398 393562 70634
rect 393646 70398 393882 70634
rect 393326 34718 393562 34954
rect 393646 34718 393882 34954
rect 393326 34398 393562 34634
rect 393646 34398 393882 34634
rect 393326 -7302 393562 -7066
rect 393646 -7302 393882 -7066
rect 393326 -7622 393562 -7386
rect 393646 -7622 393882 -7386
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 402326 223718 402562 223954
rect 402646 223718 402882 223954
rect 402326 223398 402562 223634
rect 402646 223398 402882 223634
rect 402326 187718 402562 187954
rect 402646 187718 402882 187954
rect 402326 187398 402562 187634
rect 402646 187398 402882 187634
rect 402326 151718 402562 151954
rect 402646 151718 402882 151954
rect 402326 151398 402562 151634
rect 402646 151398 402882 151634
rect 402326 115718 402562 115954
rect 402646 115718 402882 115954
rect 402326 115398 402562 115634
rect 402646 115398 402882 115634
rect 402326 79718 402562 79954
rect 402646 79718 402882 79954
rect 402326 79398 402562 79634
rect 402646 79398 402882 79634
rect 402326 43718 402562 43954
rect 402646 43718 402882 43954
rect 402326 43398 402562 43634
rect 402646 43398 402882 43634
rect 402326 7718 402562 7954
rect 402646 7718 402882 7954
rect 402326 7398 402562 7634
rect 402646 7398 402882 7634
rect 402326 -1542 402562 -1306
rect 402646 -1542 402882 -1306
rect 402326 -1862 402562 -1626
rect 402646 -1862 402882 -1626
rect 406826 228218 407062 228454
rect 407146 228218 407382 228454
rect 406826 227898 407062 228134
rect 407146 227898 407382 228134
rect 406826 192218 407062 192454
rect 407146 192218 407382 192454
rect 406826 191898 407062 192134
rect 407146 191898 407382 192134
rect 406826 156218 407062 156454
rect 407146 156218 407382 156454
rect 406826 155898 407062 156134
rect 407146 155898 407382 156134
rect 406826 120218 407062 120454
rect 407146 120218 407382 120454
rect 406826 119898 407062 120134
rect 407146 119898 407382 120134
rect 406826 84218 407062 84454
rect 407146 84218 407382 84454
rect 406826 83898 407062 84134
rect 407146 83898 407382 84134
rect 406826 48218 407062 48454
rect 407146 48218 407382 48454
rect 406826 47898 407062 48134
rect 407146 47898 407382 48134
rect 406826 12218 407062 12454
rect 407146 12218 407382 12454
rect 406826 11898 407062 12134
rect 407146 11898 407382 12134
rect 406826 -2502 407062 -2266
rect 407146 -2502 407382 -2266
rect 406826 -2822 407062 -2586
rect 407146 -2822 407382 -2586
rect 411326 707482 411562 707718
rect 411646 707482 411882 707718
rect 411326 707162 411562 707398
rect 411646 707162 411882 707398
rect 411326 700718 411562 700954
rect 411646 700718 411882 700954
rect 411326 700398 411562 700634
rect 411646 700398 411882 700634
rect 411326 664718 411562 664954
rect 411646 664718 411882 664954
rect 411326 664398 411562 664634
rect 411646 664398 411882 664634
rect 411326 628718 411562 628954
rect 411646 628718 411882 628954
rect 411326 628398 411562 628634
rect 411646 628398 411882 628634
rect 411326 592718 411562 592954
rect 411646 592718 411882 592954
rect 411326 592398 411562 592634
rect 411646 592398 411882 592634
rect 411326 556718 411562 556954
rect 411646 556718 411882 556954
rect 411326 556398 411562 556634
rect 411646 556398 411882 556634
rect 411326 520718 411562 520954
rect 411646 520718 411882 520954
rect 411326 520398 411562 520634
rect 411646 520398 411882 520634
rect 411326 484718 411562 484954
rect 411646 484718 411882 484954
rect 411326 484398 411562 484634
rect 411646 484398 411882 484634
rect 411326 448718 411562 448954
rect 411646 448718 411882 448954
rect 411326 448398 411562 448634
rect 411646 448398 411882 448634
rect 411326 412718 411562 412954
rect 411646 412718 411882 412954
rect 411326 412398 411562 412634
rect 411646 412398 411882 412634
rect 411326 376718 411562 376954
rect 411646 376718 411882 376954
rect 411326 376398 411562 376634
rect 411646 376398 411882 376634
rect 411326 340718 411562 340954
rect 411646 340718 411882 340954
rect 411326 340398 411562 340634
rect 411646 340398 411882 340634
rect 411326 304718 411562 304954
rect 411646 304718 411882 304954
rect 411326 304398 411562 304634
rect 411646 304398 411882 304634
rect 411326 268718 411562 268954
rect 411646 268718 411882 268954
rect 411326 268398 411562 268634
rect 411646 268398 411882 268634
rect 411326 232718 411562 232954
rect 411646 232718 411882 232954
rect 411326 232398 411562 232634
rect 411646 232398 411882 232634
rect 411326 196718 411562 196954
rect 411646 196718 411882 196954
rect 411326 196398 411562 196634
rect 411646 196398 411882 196634
rect 411326 160718 411562 160954
rect 411646 160718 411882 160954
rect 411326 160398 411562 160634
rect 411646 160398 411882 160634
rect 411326 124718 411562 124954
rect 411646 124718 411882 124954
rect 411326 124398 411562 124634
rect 411646 124398 411882 124634
rect 411326 88718 411562 88954
rect 411646 88718 411882 88954
rect 411326 88398 411562 88634
rect 411646 88398 411882 88634
rect 411326 52718 411562 52954
rect 411646 52718 411882 52954
rect 411326 52398 411562 52634
rect 411646 52398 411882 52634
rect 411326 16718 411562 16954
rect 411646 16718 411882 16954
rect 411326 16398 411562 16634
rect 411646 16398 411882 16634
rect 411326 -3462 411562 -3226
rect 411646 -3462 411882 -3226
rect 411326 -3782 411562 -3546
rect 411646 -3782 411882 -3546
rect 415826 708442 416062 708678
rect 416146 708442 416382 708678
rect 415826 708122 416062 708358
rect 416146 708122 416382 708358
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -4422 416062 -4186
rect 416146 -4422 416382 -4186
rect 415826 -4742 416062 -4506
rect 416146 -4742 416382 -4506
rect 420326 709402 420562 709638
rect 420646 709402 420882 709638
rect 420326 709082 420562 709318
rect 420646 709082 420882 709318
rect 420326 673718 420562 673954
rect 420646 673718 420882 673954
rect 420326 673398 420562 673634
rect 420646 673398 420882 673634
rect 420326 637718 420562 637954
rect 420646 637718 420882 637954
rect 420326 637398 420562 637634
rect 420646 637398 420882 637634
rect 420326 601718 420562 601954
rect 420646 601718 420882 601954
rect 420326 601398 420562 601634
rect 420646 601398 420882 601634
rect 420326 565718 420562 565954
rect 420646 565718 420882 565954
rect 420326 565398 420562 565634
rect 420646 565398 420882 565634
rect 420326 529718 420562 529954
rect 420646 529718 420882 529954
rect 420326 529398 420562 529634
rect 420646 529398 420882 529634
rect 420326 493718 420562 493954
rect 420646 493718 420882 493954
rect 420326 493398 420562 493634
rect 420646 493398 420882 493634
rect 420326 457718 420562 457954
rect 420646 457718 420882 457954
rect 420326 457398 420562 457634
rect 420646 457398 420882 457634
rect 420326 421718 420562 421954
rect 420646 421718 420882 421954
rect 420326 421398 420562 421634
rect 420646 421398 420882 421634
rect 420326 385718 420562 385954
rect 420646 385718 420882 385954
rect 420326 385398 420562 385634
rect 420646 385398 420882 385634
rect 420326 349718 420562 349954
rect 420646 349718 420882 349954
rect 420326 349398 420562 349634
rect 420646 349398 420882 349634
rect 420326 313718 420562 313954
rect 420646 313718 420882 313954
rect 420326 313398 420562 313634
rect 420646 313398 420882 313634
rect 420326 277718 420562 277954
rect 420646 277718 420882 277954
rect 420326 277398 420562 277634
rect 420646 277398 420882 277634
rect 420326 241718 420562 241954
rect 420646 241718 420882 241954
rect 420326 241398 420562 241634
rect 420646 241398 420882 241634
rect 420326 205718 420562 205954
rect 420646 205718 420882 205954
rect 420326 205398 420562 205634
rect 420646 205398 420882 205634
rect 420326 169718 420562 169954
rect 420646 169718 420882 169954
rect 420326 169398 420562 169634
rect 420646 169398 420882 169634
rect 420326 133718 420562 133954
rect 420646 133718 420882 133954
rect 420326 133398 420562 133634
rect 420646 133398 420882 133634
rect 420326 97718 420562 97954
rect 420646 97718 420882 97954
rect 420326 97398 420562 97634
rect 420646 97398 420882 97634
rect 420326 61718 420562 61954
rect 420646 61718 420882 61954
rect 420326 61398 420562 61634
rect 420646 61398 420882 61634
rect 420326 25718 420562 25954
rect 420646 25718 420882 25954
rect 420326 25398 420562 25634
rect 420646 25398 420882 25634
rect 420326 -5382 420562 -5146
rect 420646 -5382 420882 -5146
rect 420326 -5702 420562 -5466
rect 420646 -5702 420882 -5466
rect 424826 710362 425062 710598
rect 425146 710362 425382 710598
rect 424826 710042 425062 710278
rect 425146 710042 425382 710278
rect 424826 678218 425062 678454
rect 425146 678218 425382 678454
rect 424826 677898 425062 678134
rect 425146 677898 425382 678134
rect 424826 642218 425062 642454
rect 425146 642218 425382 642454
rect 424826 641898 425062 642134
rect 425146 641898 425382 642134
rect 424826 606218 425062 606454
rect 425146 606218 425382 606454
rect 424826 605898 425062 606134
rect 425146 605898 425382 606134
rect 424826 570218 425062 570454
rect 425146 570218 425382 570454
rect 424826 569898 425062 570134
rect 425146 569898 425382 570134
rect 424826 534218 425062 534454
rect 425146 534218 425382 534454
rect 424826 533898 425062 534134
rect 425146 533898 425382 534134
rect 424826 498218 425062 498454
rect 425146 498218 425382 498454
rect 424826 497898 425062 498134
rect 425146 497898 425382 498134
rect 424826 462218 425062 462454
rect 425146 462218 425382 462454
rect 424826 461898 425062 462134
rect 425146 461898 425382 462134
rect 424826 426218 425062 426454
rect 425146 426218 425382 426454
rect 424826 425898 425062 426134
rect 425146 425898 425382 426134
rect 424826 390218 425062 390454
rect 425146 390218 425382 390454
rect 424826 389898 425062 390134
rect 425146 389898 425382 390134
rect 424826 354218 425062 354454
rect 425146 354218 425382 354454
rect 424826 353898 425062 354134
rect 425146 353898 425382 354134
rect 424826 318218 425062 318454
rect 425146 318218 425382 318454
rect 424826 317898 425062 318134
rect 425146 317898 425382 318134
rect 424826 282218 425062 282454
rect 425146 282218 425382 282454
rect 424826 281898 425062 282134
rect 425146 281898 425382 282134
rect 424826 246218 425062 246454
rect 425146 246218 425382 246454
rect 424826 245898 425062 246134
rect 425146 245898 425382 246134
rect 424826 210218 425062 210454
rect 425146 210218 425382 210454
rect 424826 209898 425062 210134
rect 425146 209898 425382 210134
rect 424826 174218 425062 174454
rect 425146 174218 425382 174454
rect 424826 173898 425062 174134
rect 425146 173898 425382 174134
rect 424826 138218 425062 138454
rect 425146 138218 425382 138454
rect 424826 137898 425062 138134
rect 425146 137898 425382 138134
rect 424826 102218 425062 102454
rect 425146 102218 425382 102454
rect 424826 101898 425062 102134
rect 425146 101898 425382 102134
rect 424826 66218 425062 66454
rect 425146 66218 425382 66454
rect 424826 65898 425062 66134
rect 425146 65898 425382 66134
rect 424826 30218 425062 30454
rect 425146 30218 425382 30454
rect 424826 29898 425062 30134
rect 425146 29898 425382 30134
rect 424826 -6342 425062 -6106
rect 425146 -6342 425382 -6106
rect 424826 -6662 425062 -6426
rect 425146 -6662 425382 -6426
rect 429326 711322 429562 711558
rect 429646 711322 429882 711558
rect 429326 711002 429562 711238
rect 429646 711002 429882 711238
rect 429326 682718 429562 682954
rect 429646 682718 429882 682954
rect 429326 682398 429562 682634
rect 429646 682398 429882 682634
rect 429326 646718 429562 646954
rect 429646 646718 429882 646954
rect 429326 646398 429562 646634
rect 429646 646398 429882 646634
rect 429326 610718 429562 610954
rect 429646 610718 429882 610954
rect 429326 610398 429562 610634
rect 429646 610398 429882 610634
rect 429326 574718 429562 574954
rect 429646 574718 429882 574954
rect 429326 574398 429562 574634
rect 429646 574398 429882 574634
rect 429326 538718 429562 538954
rect 429646 538718 429882 538954
rect 429326 538398 429562 538634
rect 429646 538398 429882 538634
rect 429326 502718 429562 502954
rect 429646 502718 429882 502954
rect 429326 502398 429562 502634
rect 429646 502398 429882 502634
rect 429326 466718 429562 466954
rect 429646 466718 429882 466954
rect 429326 466398 429562 466634
rect 429646 466398 429882 466634
rect 429326 430718 429562 430954
rect 429646 430718 429882 430954
rect 429326 430398 429562 430634
rect 429646 430398 429882 430634
rect 429326 394718 429562 394954
rect 429646 394718 429882 394954
rect 429326 394398 429562 394634
rect 429646 394398 429882 394634
rect 429326 358718 429562 358954
rect 429646 358718 429882 358954
rect 429326 358398 429562 358634
rect 429646 358398 429882 358634
rect 429326 322718 429562 322954
rect 429646 322718 429882 322954
rect 429326 322398 429562 322634
rect 429646 322398 429882 322634
rect 429326 286718 429562 286954
rect 429646 286718 429882 286954
rect 429326 286398 429562 286634
rect 429646 286398 429882 286634
rect 429326 250718 429562 250954
rect 429646 250718 429882 250954
rect 429326 250398 429562 250634
rect 429646 250398 429882 250634
rect 429326 214718 429562 214954
rect 429646 214718 429882 214954
rect 429326 214398 429562 214634
rect 429646 214398 429882 214634
rect 429326 178718 429562 178954
rect 429646 178718 429882 178954
rect 429326 178398 429562 178634
rect 429646 178398 429882 178634
rect 429326 142718 429562 142954
rect 429646 142718 429882 142954
rect 429326 142398 429562 142634
rect 429646 142398 429882 142634
rect 429326 106718 429562 106954
rect 429646 106718 429882 106954
rect 429326 106398 429562 106634
rect 429646 106398 429882 106634
rect 429326 70718 429562 70954
rect 429646 70718 429882 70954
rect 429326 70398 429562 70634
rect 429646 70398 429882 70634
rect 429326 34718 429562 34954
rect 429646 34718 429882 34954
rect 429326 34398 429562 34634
rect 429646 34398 429882 34634
rect 429326 -7302 429562 -7066
rect 429646 -7302 429882 -7066
rect 429326 -7622 429562 -7386
rect 429646 -7622 429882 -7386
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 438326 705562 438562 705798
rect 438646 705562 438882 705798
rect 438326 705242 438562 705478
rect 438646 705242 438882 705478
rect 438326 691718 438562 691954
rect 438646 691718 438882 691954
rect 438326 691398 438562 691634
rect 438646 691398 438882 691634
rect 438326 655718 438562 655954
rect 438646 655718 438882 655954
rect 438326 655398 438562 655634
rect 438646 655398 438882 655634
rect 438326 619718 438562 619954
rect 438646 619718 438882 619954
rect 438326 619398 438562 619634
rect 438646 619398 438882 619634
rect 438326 583718 438562 583954
rect 438646 583718 438882 583954
rect 438326 583398 438562 583634
rect 438646 583398 438882 583634
rect 438326 547718 438562 547954
rect 438646 547718 438882 547954
rect 438326 547398 438562 547634
rect 438646 547398 438882 547634
rect 438326 511718 438562 511954
rect 438646 511718 438882 511954
rect 438326 511398 438562 511634
rect 438646 511398 438882 511634
rect 438326 475718 438562 475954
rect 438646 475718 438882 475954
rect 438326 475398 438562 475634
rect 438646 475398 438882 475634
rect 438326 439718 438562 439954
rect 438646 439718 438882 439954
rect 438326 439398 438562 439634
rect 438646 439398 438882 439634
rect 438326 403718 438562 403954
rect 438646 403718 438882 403954
rect 438326 403398 438562 403634
rect 438646 403398 438882 403634
rect 438326 367718 438562 367954
rect 438646 367718 438882 367954
rect 438326 367398 438562 367634
rect 438646 367398 438882 367634
rect 438326 331718 438562 331954
rect 438646 331718 438882 331954
rect 438326 331398 438562 331634
rect 438646 331398 438882 331634
rect 438326 295718 438562 295954
rect 438646 295718 438882 295954
rect 438326 295398 438562 295634
rect 438646 295398 438882 295634
rect 438326 259718 438562 259954
rect 438646 259718 438882 259954
rect 438326 259398 438562 259634
rect 438646 259398 438882 259634
rect 438326 223718 438562 223954
rect 438646 223718 438882 223954
rect 438326 223398 438562 223634
rect 438646 223398 438882 223634
rect 438326 187718 438562 187954
rect 438646 187718 438882 187954
rect 438326 187398 438562 187634
rect 438646 187398 438882 187634
rect 438326 151718 438562 151954
rect 438646 151718 438882 151954
rect 438326 151398 438562 151634
rect 438646 151398 438882 151634
rect 438326 115718 438562 115954
rect 438646 115718 438882 115954
rect 438326 115398 438562 115634
rect 438646 115398 438882 115634
rect 438326 79718 438562 79954
rect 438646 79718 438882 79954
rect 438326 79398 438562 79634
rect 438646 79398 438882 79634
rect 438326 43718 438562 43954
rect 438646 43718 438882 43954
rect 438326 43398 438562 43634
rect 438646 43398 438882 43634
rect 438326 7718 438562 7954
rect 438646 7718 438882 7954
rect 438326 7398 438562 7634
rect 438646 7398 438882 7634
rect 438326 -1542 438562 -1306
rect 438646 -1542 438882 -1306
rect 438326 -1862 438562 -1626
rect 438646 -1862 438882 -1626
rect 442826 706522 443062 706758
rect 443146 706522 443382 706758
rect 442826 706202 443062 706438
rect 443146 706202 443382 706438
rect 442826 696218 443062 696454
rect 443146 696218 443382 696454
rect 442826 695898 443062 696134
rect 443146 695898 443382 696134
rect 442826 660218 443062 660454
rect 443146 660218 443382 660454
rect 442826 659898 443062 660134
rect 443146 659898 443382 660134
rect 442826 624218 443062 624454
rect 443146 624218 443382 624454
rect 442826 623898 443062 624134
rect 443146 623898 443382 624134
rect 442826 588218 443062 588454
rect 443146 588218 443382 588454
rect 442826 587898 443062 588134
rect 443146 587898 443382 588134
rect 442826 552218 443062 552454
rect 443146 552218 443382 552454
rect 442826 551898 443062 552134
rect 443146 551898 443382 552134
rect 442826 516218 443062 516454
rect 443146 516218 443382 516454
rect 442826 515898 443062 516134
rect 443146 515898 443382 516134
rect 442826 480218 443062 480454
rect 443146 480218 443382 480454
rect 442826 479898 443062 480134
rect 443146 479898 443382 480134
rect 442826 444218 443062 444454
rect 443146 444218 443382 444454
rect 442826 443898 443062 444134
rect 443146 443898 443382 444134
rect 442826 408218 443062 408454
rect 443146 408218 443382 408454
rect 442826 407898 443062 408134
rect 443146 407898 443382 408134
rect 442826 372218 443062 372454
rect 443146 372218 443382 372454
rect 442826 371898 443062 372134
rect 443146 371898 443382 372134
rect 442826 336218 443062 336454
rect 443146 336218 443382 336454
rect 442826 335898 443062 336134
rect 443146 335898 443382 336134
rect 442826 300218 443062 300454
rect 443146 300218 443382 300454
rect 442826 299898 443062 300134
rect 443146 299898 443382 300134
rect 442826 264218 443062 264454
rect 443146 264218 443382 264454
rect 442826 263898 443062 264134
rect 443146 263898 443382 264134
rect 442826 228218 443062 228454
rect 443146 228218 443382 228454
rect 442826 227898 443062 228134
rect 443146 227898 443382 228134
rect 442826 192218 443062 192454
rect 443146 192218 443382 192454
rect 442826 191898 443062 192134
rect 443146 191898 443382 192134
rect 442826 156218 443062 156454
rect 443146 156218 443382 156454
rect 442826 155898 443062 156134
rect 443146 155898 443382 156134
rect 442826 120218 443062 120454
rect 443146 120218 443382 120454
rect 442826 119898 443062 120134
rect 443146 119898 443382 120134
rect 442826 84218 443062 84454
rect 443146 84218 443382 84454
rect 442826 83898 443062 84134
rect 443146 83898 443382 84134
rect 442826 48218 443062 48454
rect 443146 48218 443382 48454
rect 442826 47898 443062 48134
rect 443146 47898 443382 48134
rect 442826 12218 443062 12454
rect 443146 12218 443382 12454
rect 442826 11898 443062 12134
rect 443146 11898 443382 12134
rect 442826 -2502 443062 -2266
rect 443146 -2502 443382 -2266
rect 442826 -2822 443062 -2586
rect 443146 -2822 443382 -2586
rect 447326 707482 447562 707718
rect 447646 707482 447882 707718
rect 447326 707162 447562 707398
rect 447646 707162 447882 707398
rect 447326 700718 447562 700954
rect 447646 700718 447882 700954
rect 447326 700398 447562 700634
rect 447646 700398 447882 700634
rect 447326 664718 447562 664954
rect 447646 664718 447882 664954
rect 447326 664398 447562 664634
rect 447646 664398 447882 664634
rect 447326 628718 447562 628954
rect 447646 628718 447882 628954
rect 447326 628398 447562 628634
rect 447646 628398 447882 628634
rect 447326 592718 447562 592954
rect 447646 592718 447882 592954
rect 447326 592398 447562 592634
rect 447646 592398 447882 592634
rect 447326 556718 447562 556954
rect 447646 556718 447882 556954
rect 447326 556398 447562 556634
rect 447646 556398 447882 556634
rect 447326 520718 447562 520954
rect 447646 520718 447882 520954
rect 447326 520398 447562 520634
rect 447646 520398 447882 520634
rect 447326 484718 447562 484954
rect 447646 484718 447882 484954
rect 447326 484398 447562 484634
rect 447646 484398 447882 484634
rect 447326 448718 447562 448954
rect 447646 448718 447882 448954
rect 447326 448398 447562 448634
rect 447646 448398 447882 448634
rect 447326 412718 447562 412954
rect 447646 412718 447882 412954
rect 447326 412398 447562 412634
rect 447646 412398 447882 412634
rect 447326 376718 447562 376954
rect 447646 376718 447882 376954
rect 447326 376398 447562 376634
rect 447646 376398 447882 376634
rect 447326 340718 447562 340954
rect 447646 340718 447882 340954
rect 447326 340398 447562 340634
rect 447646 340398 447882 340634
rect 447326 304718 447562 304954
rect 447646 304718 447882 304954
rect 447326 304398 447562 304634
rect 447646 304398 447882 304634
rect 447326 268718 447562 268954
rect 447646 268718 447882 268954
rect 447326 268398 447562 268634
rect 447646 268398 447882 268634
rect 447326 232718 447562 232954
rect 447646 232718 447882 232954
rect 447326 232398 447562 232634
rect 447646 232398 447882 232634
rect 447326 196718 447562 196954
rect 447646 196718 447882 196954
rect 447326 196398 447562 196634
rect 447646 196398 447882 196634
rect 447326 160718 447562 160954
rect 447646 160718 447882 160954
rect 447326 160398 447562 160634
rect 447646 160398 447882 160634
rect 447326 124718 447562 124954
rect 447646 124718 447882 124954
rect 447326 124398 447562 124634
rect 447646 124398 447882 124634
rect 447326 88718 447562 88954
rect 447646 88718 447882 88954
rect 447326 88398 447562 88634
rect 447646 88398 447882 88634
rect 447326 52718 447562 52954
rect 447646 52718 447882 52954
rect 447326 52398 447562 52634
rect 447646 52398 447882 52634
rect 447326 16718 447562 16954
rect 447646 16718 447882 16954
rect 447326 16398 447562 16634
rect 447646 16398 447882 16634
rect 447326 -3462 447562 -3226
rect 447646 -3462 447882 -3226
rect 447326 -3782 447562 -3546
rect 447646 -3782 447882 -3546
rect 451826 708442 452062 708678
rect 452146 708442 452382 708678
rect 451826 708122 452062 708358
rect 452146 708122 452382 708358
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -4422 452062 -4186
rect 452146 -4422 452382 -4186
rect 451826 -4742 452062 -4506
rect 452146 -4742 452382 -4506
rect 456326 709402 456562 709638
rect 456646 709402 456882 709638
rect 456326 709082 456562 709318
rect 456646 709082 456882 709318
rect 456326 673718 456562 673954
rect 456646 673718 456882 673954
rect 456326 673398 456562 673634
rect 456646 673398 456882 673634
rect 456326 637718 456562 637954
rect 456646 637718 456882 637954
rect 456326 637398 456562 637634
rect 456646 637398 456882 637634
rect 456326 601718 456562 601954
rect 456646 601718 456882 601954
rect 456326 601398 456562 601634
rect 456646 601398 456882 601634
rect 456326 565718 456562 565954
rect 456646 565718 456882 565954
rect 456326 565398 456562 565634
rect 456646 565398 456882 565634
rect 456326 529718 456562 529954
rect 456646 529718 456882 529954
rect 456326 529398 456562 529634
rect 456646 529398 456882 529634
rect 456326 493718 456562 493954
rect 456646 493718 456882 493954
rect 456326 493398 456562 493634
rect 456646 493398 456882 493634
rect 456326 457718 456562 457954
rect 456646 457718 456882 457954
rect 456326 457398 456562 457634
rect 456646 457398 456882 457634
rect 456326 421718 456562 421954
rect 456646 421718 456882 421954
rect 456326 421398 456562 421634
rect 456646 421398 456882 421634
rect 456326 385718 456562 385954
rect 456646 385718 456882 385954
rect 456326 385398 456562 385634
rect 456646 385398 456882 385634
rect 456326 349718 456562 349954
rect 456646 349718 456882 349954
rect 456326 349398 456562 349634
rect 456646 349398 456882 349634
rect 456326 313718 456562 313954
rect 456646 313718 456882 313954
rect 456326 313398 456562 313634
rect 456646 313398 456882 313634
rect 456326 277718 456562 277954
rect 456646 277718 456882 277954
rect 456326 277398 456562 277634
rect 456646 277398 456882 277634
rect 456326 241718 456562 241954
rect 456646 241718 456882 241954
rect 456326 241398 456562 241634
rect 456646 241398 456882 241634
rect 456326 205718 456562 205954
rect 456646 205718 456882 205954
rect 456326 205398 456562 205634
rect 456646 205398 456882 205634
rect 456326 169718 456562 169954
rect 456646 169718 456882 169954
rect 456326 169398 456562 169634
rect 456646 169398 456882 169634
rect 456326 133718 456562 133954
rect 456646 133718 456882 133954
rect 456326 133398 456562 133634
rect 456646 133398 456882 133634
rect 456326 97718 456562 97954
rect 456646 97718 456882 97954
rect 456326 97398 456562 97634
rect 456646 97398 456882 97634
rect 456326 61718 456562 61954
rect 456646 61718 456882 61954
rect 456326 61398 456562 61634
rect 456646 61398 456882 61634
rect 456326 25718 456562 25954
rect 456646 25718 456882 25954
rect 456326 25398 456562 25634
rect 456646 25398 456882 25634
rect 456326 -5382 456562 -5146
rect 456646 -5382 456882 -5146
rect 456326 -5702 456562 -5466
rect 456646 -5702 456882 -5466
rect 460826 710362 461062 710598
rect 461146 710362 461382 710598
rect 460826 710042 461062 710278
rect 461146 710042 461382 710278
rect 460826 678218 461062 678454
rect 461146 678218 461382 678454
rect 460826 677898 461062 678134
rect 461146 677898 461382 678134
rect 460826 642218 461062 642454
rect 461146 642218 461382 642454
rect 460826 641898 461062 642134
rect 461146 641898 461382 642134
rect 460826 606218 461062 606454
rect 461146 606218 461382 606454
rect 460826 605898 461062 606134
rect 461146 605898 461382 606134
rect 460826 570218 461062 570454
rect 461146 570218 461382 570454
rect 460826 569898 461062 570134
rect 461146 569898 461382 570134
rect 460826 534218 461062 534454
rect 461146 534218 461382 534454
rect 460826 533898 461062 534134
rect 461146 533898 461382 534134
rect 460826 498218 461062 498454
rect 461146 498218 461382 498454
rect 460826 497898 461062 498134
rect 461146 497898 461382 498134
rect 460826 462218 461062 462454
rect 461146 462218 461382 462454
rect 460826 461898 461062 462134
rect 461146 461898 461382 462134
rect 460826 426218 461062 426454
rect 461146 426218 461382 426454
rect 460826 425898 461062 426134
rect 461146 425898 461382 426134
rect 460826 390218 461062 390454
rect 461146 390218 461382 390454
rect 460826 389898 461062 390134
rect 461146 389898 461382 390134
rect 460826 354218 461062 354454
rect 461146 354218 461382 354454
rect 460826 353898 461062 354134
rect 461146 353898 461382 354134
rect 460826 318218 461062 318454
rect 461146 318218 461382 318454
rect 460826 317898 461062 318134
rect 461146 317898 461382 318134
rect 460826 282218 461062 282454
rect 461146 282218 461382 282454
rect 460826 281898 461062 282134
rect 461146 281898 461382 282134
rect 460826 246218 461062 246454
rect 461146 246218 461382 246454
rect 460826 245898 461062 246134
rect 461146 245898 461382 246134
rect 460826 210218 461062 210454
rect 461146 210218 461382 210454
rect 460826 209898 461062 210134
rect 461146 209898 461382 210134
rect 460826 174218 461062 174454
rect 461146 174218 461382 174454
rect 460826 173898 461062 174134
rect 461146 173898 461382 174134
rect 460826 138218 461062 138454
rect 461146 138218 461382 138454
rect 460826 137898 461062 138134
rect 461146 137898 461382 138134
rect 460826 102218 461062 102454
rect 461146 102218 461382 102454
rect 460826 101898 461062 102134
rect 461146 101898 461382 102134
rect 460826 66218 461062 66454
rect 461146 66218 461382 66454
rect 460826 65898 461062 66134
rect 461146 65898 461382 66134
rect 460826 30218 461062 30454
rect 461146 30218 461382 30454
rect 460826 29898 461062 30134
rect 461146 29898 461382 30134
rect 460826 -6342 461062 -6106
rect 461146 -6342 461382 -6106
rect 460826 -6662 461062 -6426
rect 461146 -6662 461382 -6426
rect 465326 711322 465562 711558
rect 465646 711322 465882 711558
rect 465326 711002 465562 711238
rect 465646 711002 465882 711238
rect 465326 682718 465562 682954
rect 465646 682718 465882 682954
rect 465326 682398 465562 682634
rect 465646 682398 465882 682634
rect 465326 646718 465562 646954
rect 465646 646718 465882 646954
rect 465326 646398 465562 646634
rect 465646 646398 465882 646634
rect 465326 610718 465562 610954
rect 465646 610718 465882 610954
rect 465326 610398 465562 610634
rect 465646 610398 465882 610634
rect 465326 574718 465562 574954
rect 465646 574718 465882 574954
rect 465326 574398 465562 574634
rect 465646 574398 465882 574634
rect 465326 538718 465562 538954
rect 465646 538718 465882 538954
rect 465326 538398 465562 538634
rect 465646 538398 465882 538634
rect 465326 502718 465562 502954
rect 465646 502718 465882 502954
rect 465326 502398 465562 502634
rect 465646 502398 465882 502634
rect 465326 466718 465562 466954
rect 465646 466718 465882 466954
rect 465326 466398 465562 466634
rect 465646 466398 465882 466634
rect 465326 430718 465562 430954
rect 465646 430718 465882 430954
rect 465326 430398 465562 430634
rect 465646 430398 465882 430634
rect 465326 394718 465562 394954
rect 465646 394718 465882 394954
rect 465326 394398 465562 394634
rect 465646 394398 465882 394634
rect 465326 358718 465562 358954
rect 465646 358718 465882 358954
rect 465326 358398 465562 358634
rect 465646 358398 465882 358634
rect 465326 322718 465562 322954
rect 465646 322718 465882 322954
rect 465326 322398 465562 322634
rect 465646 322398 465882 322634
rect 465326 286718 465562 286954
rect 465646 286718 465882 286954
rect 465326 286398 465562 286634
rect 465646 286398 465882 286634
rect 465326 250718 465562 250954
rect 465646 250718 465882 250954
rect 465326 250398 465562 250634
rect 465646 250398 465882 250634
rect 465326 214718 465562 214954
rect 465646 214718 465882 214954
rect 465326 214398 465562 214634
rect 465646 214398 465882 214634
rect 465326 178718 465562 178954
rect 465646 178718 465882 178954
rect 465326 178398 465562 178634
rect 465646 178398 465882 178634
rect 465326 142718 465562 142954
rect 465646 142718 465882 142954
rect 465326 142398 465562 142634
rect 465646 142398 465882 142634
rect 465326 106718 465562 106954
rect 465646 106718 465882 106954
rect 465326 106398 465562 106634
rect 465646 106398 465882 106634
rect 465326 70718 465562 70954
rect 465646 70718 465882 70954
rect 465326 70398 465562 70634
rect 465646 70398 465882 70634
rect 465326 34718 465562 34954
rect 465646 34718 465882 34954
rect 465326 34398 465562 34634
rect 465646 34398 465882 34634
rect 465326 -7302 465562 -7066
rect 465646 -7302 465882 -7066
rect 465326 -7622 465562 -7386
rect 465646 -7622 465882 -7386
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 474326 705562 474562 705798
rect 474646 705562 474882 705798
rect 474326 705242 474562 705478
rect 474646 705242 474882 705478
rect 474326 691718 474562 691954
rect 474646 691718 474882 691954
rect 474326 691398 474562 691634
rect 474646 691398 474882 691634
rect 474326 655718 474562 655954
rect 474646 655718 474882 655954
rect 474326 655398 474562 655634
rect 474646 655398 474882 655634
rect 474326 619718 474562 619954
rect 474646 619718 474882 619954
rect 474326 619398 474562 619634
rect 474646 619398 474882 619634
rect 474326 583718 474562 583954
rect 474646 583718 474882 583954
rect 474326 583398 474562 583634
rect 474646 583398 474882 583634
rect 474326 547718 474562 547954
rect 474646 547718 474882 547954
rect 474326 547398 474562 547634
rect 474646 547398 474882 547634
rect 474326 511718 474562 511954
rect 474646 511718 474882 511954
rect 474326 511398 474562 511634
rect 474646 511398 474882 511634
rect 474326 475718 474562 475954
rect 474646 475718 474882 475954
rect 474326 475398 474562 475634
rect 474646 475398 474882 475634
rect 474326 439718 474562 439954
rect 474646 439718 474882 439954
rect 474326 439398 474562 439634
rect 474646 439398 474882 439634
rect 474326 403718 474562 403954
rect 474646 403718 474882 403954
rect 474326 403398 474562 403634
rect 474646 403398 474882 403634
rect 474326 367718 474562 367954
rect 474646 367718 474882 367954
rect 474326 367398 474562 367634
rect 474646 367398 474882 367634
rect 474326 331718 474562 331954
rect 474646 331718 474882 331954
rect 474326 331398 474562 331634
rect 474646 331398 474882 331634
rect 474326 295718 474562 295954
rect 474646 295718 474882 295954
rect 474326 295398 474562 295634
rect 474646 295398 474882 295634
rect 474326 259718 474562 259954
rect 474646 259718 474882 259954
rect 474326 259398 474562 259634
rect 474646 259398 474882 259634
rect 474326 223718 474562 223954
rect 474646 223718 474882 223954
rect 474326 223398 474562 223634
rect 474646 223398 474882 223634
rect 474326 187718 474562 187954
rect 474646 187718 474882 187954
rect 474326 187398 474562 187634
rect 474646 187398 474882 187634
rect 474326 151718 474562 151954
rect 474646 151718 474882 151954
rect 474326 151398 474562 151634
rect 474646 151398 474882 151634
rect 474326 115718 474562 115954
rect 474646 115718 474882 115954
rect 474326 115398 474562 115634
rect 474646 115398 474882 115634
rect 474326 79718 474562 79954
rect 474646 79718 474882 79954
rect 474326 79398 474562 79634
rect 474646 79398 474882 79634
rect 474326 43718 474562 43954
rect 474646 43718 474882 43954
rect 474326 43398 474562 43634
rect 474646 43398 474882 43634
rect 474326 7718 474562 7954
rect 474646 7718 474882 7954
rect 474326 7398 474562 7634
rect 474646 7398 474882 7634
rect 474326 -1542 474562 -1306
rect 474646 -1542 474882 -1306
rect 474326 -1862 474562 -1626
rect 474646 -1862 474882 -1626
rect 478826 706522 479062 706758
rect 479146 706522 479382 706758
rect 478826 706202 479062 706438
rect 479146 706202 479382 706438
rect 478826 696218 479062 696454
rect 479146 696218 479382 696454
rect 478826 695898 479062 696134
rect 479146 695898 479382 696134
rect 478826 660218 479062 660454
rect 479146 660218 479382 660454
rect 478826 659898 479062 660134
rect 479146 659898 479382 660134
rect 478826 624218 479062 624454
rect 479146 624218 479382 624454
rect 478826 623898 479062 624134
rect 479146 623898 479382 624134
rect 478826 588218 479062 588454
rect 479146 588218 479382 588454
rect 478826 587898 479062 588134
rect 479146 587898 479382 588134
rect 478826 552218 479062 552454
rect 479146 552218 479382 552454
rect 478826 551898 479062 552134
rect 479146 551898 479382 552134
rect 478826 516218 479062 516454
rect 479146 516218 479382 516454
rect 478826 515898 479062 516134
rect 479146 515898 479382 516134
rect 478826 480218 479062 480454
rect 479146 480218 479382 480454
rect 478826 479898 479062 480134
rect 479146 479898 479382 480134
rect 478826 444218 479062 444454
rect 479146 444218 479382 444454
rect 478826 443898 479062 444134
rect 479146 443898 479382 444134
rect 478826 408218 479062 408454
rect 479146 408218 479382 408454
rect 478826 407898 479062 408134
rect 479146 407898 479382 408134
rect 478826 372218 479062 372454
rect 479146 372218 479382 372454
rect 478826 371898 479062 372134
rect 479146 371898 479382 372134
rect 478826 336218 479062 336454
rect 479146 336218 479382 336454
rect 478826 335898 479062 336134
rect 479146 335898 479382 336134
rect 478826 300218 479062 300454
rect 479146 300218 479382 300454
rect 478826 299898 479062 300134
rect 479146 299898 479382 300134
rect 478826 264218 479062 264454
rect 479146 264218 479382 264454
rect 478826 263898 479062 264134
rect 479146 263898 479382 264134
rect 478826 228218 479062 228454
rect 479146 228218 479382 228454
rect 478826 227898 479062 228134
rect 479146 227898 479382 228134
rect 478826 192218 479062 192454
rect 479146 192218 479382 192454
rect 478826 191898 479062 192134
rect 479146 191898 479382 192134
rect 478826 156218 479062 156454
rect 479146 156218 479382 156454
rect 478826 155898 479062 156134
rect 479146 155898 479382 156134
rect 478826 120218 479062 120454
rect 479146 120218 479382 120454
rect 478826 119898 479062 120134
rect 479146 119898 479382 120134
rect 478826 84218 479062 84454
rect 479146 84218 479382 84454
rect 478826 83898 479062 84134
rect 479146 83898 479382 84134
rect 478826 48218 479062 48454
rect 479146 48218 479382 48454
rect 478826 47898 479062 48134
rect 479146 47898 479382 48134
rect 478826 12218 479062 12454
rect 479146 12218 479382 12454
rect 478826 11898 479062 12134
rect 479146 11898 479382 12134
rect 478826 -2502 479062 -2266
rect 479146 -2502 479382 -2266
rect 478826 -2822 479062 -2586
rect 479146 -2822 479382 -2586
rect 483326 707482 483562 707718
rect 483646 707482 483882 707718
rect 483326 707162 483562 707398
rect 483646 707162 483882 707398
rect 483326 700718 483562 700954
rect 483646 700718 483882 700954
rect 483326 700398 483562 700634
rect 483646 700398 483882 700634
rect 483326 664718 483562 664954
rect 483646 664718 483882 664954
rect 483326 664398 483562 664634
rect 483646 664398 483882 664634
rect 483326 628718 483562 628954
rect 483646 628718 483882 628954
rect 483326 628398 483562 628634
rect 483646 628398 483882 628634
rect 483326 592718 483562 592954
rect 483646 592718 483882 592954
rect 483326 592398 483562 592634
rect 483646 592398 483882 592634
rect 483326 556718 483562 556954
rect 483646 556718 483882 556954
rect 483326 556398 483562 556634
rect 483646 556398 483882 556634
rect 483326 520718 483562 520954
rect 483646 520718 483882 520954
rect 483326 520398 483562 520634
rect 483646 520398 483882 520634
rect 483326 484718 483562 484954
rect 483646 484718 483882 484954
rect 483326 484398 483562 484634
rect 483646 484398 483882 484634
rect 483326 448718 483562 448954
rect 483646 448718 483882 448954
rect 483326 448398 483562 448634
rect 483646 448398 483882 448634
rect 483326 412718 483562 412954
rect 483646 412718 483882 412954
rect 483326 412398 483562 412634
rect 483646 412398 483882 412634
rect 483326 376718 483562 376954
rect 483646 376718 483882 376954
rect 483326 376398 483562 376634
rect 483646 376398 483882 376634
rect 483326 340718 483562 340954
rect 483646 340718 483882 340954
rect 483326 340398 483562 340634
rect 483646 340398 483882 340634
rect 483326 304718 483562 304954
rect 483646 304718 483882 304954
rect 483326 304398 483562 304634
rect 483646 304398 483882 304634
rect 483326 268718 483562 268954
rect 483646 268718 483882 268954
rect 483326 268398 483562 268634
rect 483646 268398 483882 268634
rect 483326 232718 483562 232954
rect 483646 232718 483882 232954
rect 483326 232398 483562 232634
rect 483646 232398 483882 232634
rect 483326 196718 483562 196954
rect 483646 196718 483882 196954
rect 483326 196398 483562 196634
rect 483646 196398 483882 196634
rect 483326 160718 483562 160954
rect 483646 160718 483882 160954
rect 483326 160398 483562 160634
rect 483646 160398 483882 160634
rect 483326 124718 483562 124954
rect 483646 124718 483882 124954
rect 483326 124398 483562 124634
rect 483646 124398 483882 124634
rect 483326 88718 483562 88954
rect 483646 88718 483882 88954
rect 483326 88398 483562 88634
rect 483646 88398 483882 88634
rect 483326 52718 483562 52954
rect 483646 52718 483882 52954
rect 483326 52398 483562 52634
rect 483646 52398 483882 52634
rect 483326 16718 483562 16954
rect 483646 16718 483882 16954
rect 483326 16398 483562 16634
rect 483646 16398 483882 16634
rect 483326 -3462 483562 -3226
rect 483646 -3462 483882 -3226
rect 483326 -3782 483562 -3546
rect 483646 -3782 483882 -3546
rect 487826 708442 488062 708678
rect 488146 708442 488382 708678
rect 487826 708122 488062 708358
rect 488146 708122 488382 708358
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -4422 488062 -4186
rect 488146 -4422 488382 -4186
rect 487826 -4742 488062 -4506
rect 488146 -4742 488382 -4506
rect 492326 709402 492562 709638
rect 492646 709402 492882 709638
rect 492326 709082 492562 709318
rect 492646 709082 492882 709318
rect 492326 673718 492562 673954
rect 492646 673718 492882 673954
rect 492326 673398 492562 673634
rect 492646 673398 492882 673634
rect 492326 637718 492562 637954
rect 492646 637718 492882 637954
rect 492326 637398 492562 637634
rect 492646 637398 492882 637634
rect 492326 601718 492562 601954
rect 492646 601718 492882 601954
rect 492326 601398 492562 601634
rect 492646 601398 492882 601634
rect 492326 565718 492562 565954
rect 492646 565718 492882 565954
rect 492326 565398 492562 565634
rect 492646 565398 492882 565634
rect 492326 529718 492562 529954
rect 492646 529718 492882 529954
rect 492326 529398 492562 529634
rect 492646 529398 492882 529634
rect 492326 493718 492562 493954
rect 492646 493718 492882 493954
rect 492326 493398 492562 493634
rect 492646 493398 492882 493634
rect 492326 457718 492562 457954
rect 492646 457718 492882 457954
rect 492326 457398 492562 457634
rect 492646 457398 492882 457634
rect 492326 421718 492562 421954
rect 492646 421718 492882 421954
rect 492326 421398 492562 421634
rect 492646 421398 492882 421634
rect 492326 385718 492562 385954
rect 492646 385718 492882 385954
rect 492326 385398 492562 385634
rect 492646 385398 492882 385634
rect 492326 349718 492562 349954
rect 492646 349718 492882 349954
rect 492326 349398 492562 349634
rect 492646 349398 492882 349634
rect 492326 313718 492562 313954
rect 492646 313718 492882 313954
rect 492326 313398 492562 313634
rect 492646 313398 492882 313634
rect 492326 277718 492562 277954
rect 492646 277718 492882 277954
rect 492326 277398 492562 277634
rect 492646 277398 492882 277634
rect 492326 241718 492562 241954
rect 492646 241718 492882 241954
rect 492326 241398 492562 241634
rect 492646 241398 492882 241634
rect 492326 205718 492562 205954
rect 492646 205718 492882 205954
rect 492326 205398 492562 205634
rect 492646 205398 492882 205634
rect 492326 169718 492562 169954
rect 492646 169718 492882 169954
rect 492326 169398 492562 169634
rect 492646 169398 492882 169634
rect 492326 133718 492562 133954
rect 492646 133718 492882 133954
rect 492326 133398 492562 133634
rect 492646 133398 492882 133634
rect 492326 97718 492562 97954
rect 492646 97718 492882 97954
rect 492326 97398 492562 97634
rect 492646 97398 492882 97634
rect 492326 61718 492562 61954
rect 492646 61718 492882 61954
rect 492326 61398 492562 61634
rect 492646 61398 492882 61634
rect 492326 25718 492562 25954
rect 492646 25718 492882 25954
rect 492326 25398 492562 25634
rect 492646 25398 492882 25634
rect 492326 -5382 492562 -5146
rect 492646 -5382 492882 -5146
rect 492326 -5702 492562 -5466
rect 492646 -5702 492882 -5466
rect 496826 710362 497062 710598
rect 497146 710362 497382 710598
rect 496826 710042 497062 710278
rect 497146 710042 497382 710278
rect 496826 678218 497062 678454
rect 497146 678218 497382 678454
rect 496826 677898 497062 678134
rect 497146 677898 497382 678134
rect 496826 642218 497062 642454
rect 497146 642218 497382 642454
rect 496826 641898 497062 642134
rect 497146 641898 497382 642134
rect 496826 606218 497062 606454
rect 497146 606218 497382 606454
rect 496826 605898 497062 606134
rect 497146 605898 497382 606134
rect 496826 570218 497062 570454
rect 497146 570218 497382 570454
rect 496826 569898 497062 570134
rect 497146 569898 497382 570134
rect 496826 534218 497062 534454
rect 497146 534218 497382 534454
rect 496826 533898 497062 534134
rect 497146 533898 497382 534134
rect 496826 498218 497062 498454
rect 497146 498218 497382 498454
rect 496826 497898 497062 498134
rect 497146 497898 497382 498134
rect 496826 462218 497062 462454
rect 497146 462218 497382 462454
rect 496826 461898 497062 462134
rect 497146 461898 497382 462134
rect 496826 426218 497062 426454
rect 497146 426218 497382 426454
rect 496826 425898 497062 426134
rect 497146 425898 497382 426134
rect 496826 390218 497062 390454
rect 497146 390218 497382 390454
rect 496826 389898 497062 390134
rect 497146 389898 497382 390134
rect 496826 354218 497062 354454
rect 497146 354218 497382 354454
rect 496826 353898 497062 354134
rect 497146 353898 497382 354134
rect 496826 318218 497062 318454
rect 497146 318218 497382 318454
rect 496826 317898 497062 318134
rect 497146 317898 497382 318134
rect 496826 282218 497062 282454
rect 497146 282218 497382 282454
rect 496826 281898 497062 282134
rect 497146 281898 497382 282134
rect 496826 246218 497062 246454
rect 497146 246218 497382 246454
rect 496826 245898 497062 246134
rect 497146 245898 497382 246134
rect 496826 210218 497062 210454
rect 497146 210218 497382 210454
rect 496826 209898 497062 210134
rect 497146 209898 497382 210134
rect 496826 174218 497062 174454
rect 497146 174218 497382 174454
rect 496826 173898 497062 174134
rect 497146 173898 497382 174134
rect 496826 138218 497062 138454
rect 497146 138218 497382 138454
rect 496826 137898 497062 138134
rect 497146 137898 497382 138134
rect 496826 102218 497062 102454
rect 497146 102218 497382 102454
rect 496826 101898 497062 102134
rect 497146 101898 497382 102134
rect 496826 66218 497062 66454
rect 497146 66218 497382 66454
rect 496826 65898 497062 66134
rect 497146 65898 497382 66134
rect 496826 30218 497062 30454
rect 497146 30218 497382 30454
rect 496826 29898 497062 30134
rect 497146 29898 497382 30134
rect 496826 -6342 497062 -6106
rect 497146 -6342 497382 -6106
rect 496826 -6662 497062 -6426
rect 497146 -6662 497382 -6426
rect 501326 711322 501562 711558
rect 501646 711322 501882 711558
rect 501326 711002 501562 711238
rect 501646 711002 501882 711238
rect 501326 682718 501562 682954
rect 501646 682718 501882 682954
rect 501326 682398 501562 682634
rect 501646 682398 501882 682634
rect 501326 646718 501562 646954
rect 501646 646718 501882 646954
rect 501326 646398 501562 646634
rect 501646 646398 501882 646634
rect 501326 610718 501562 610954
rect 501646 610718 501882 610954
rect 501326 610398 501562 610634
rect 501646 610398 501882 610634
rect 501326 574718 501562 574954
rect 501646 574718 501882 574954
rect 501326 574398 501562 574634
rect 501646 574398 501882 574634
rect 501326 538718 501562 538954
rect 501646 538718 501882 538954
rect 501326 538398 501562 538634
rect 501646 538398 501882 538634
rect 501326 502718 501562 502954
rect 501646 502718 501882 502954
rect 501326 502398 501562 502634
rect 501646 502398 501882 502634
rect 501326 466718 501562 466954
rect 501646 466718 501882 466954
rect 501326 466398 501562 466634
rect 501646 466398 501882 466634
rect 501326 430718 501562 430954
rect 501646 430718 501882 430954
rect 501326 430398 501562 430634
rect 501646 430398 501882 430634
rect 501326 394718 501562 394954
rect 501646 394718 501882 394954
rect 501326 394398 501562 394634
rect 501646 394398 501882 394634
rect 501326 358718 501562 358954
rect 501646 358718 501882 358954
rect 501326 358398 501562 358634
rect 501646 358398 501882 358634
rect 501326 322718 501562 322954
rect 501646 322718 501882 322954
rect 501326 322398 501562 322634
rect 501646 322398 501882 322634
rect 501326 286718 501562 286954
rect 501646 286718 501882 286954
rect 501326 286398 501562 286634
rect 501646 286398 501882 286634
rect 501326 250718 501562 250954
rect 501646 250718 501882 250954
rect 501326 250398 501562 250634
rect 501646 250398 501882 250634
rect 501326 214718 501562 214954
rect 501646 214718 501882 214954
rect 501326 214398 501562 214634
rect 501646 214398 501882 214634
rect 501326 178718 501562 178954
rect 501646 178718 501882 178954
rect 501326 178398 501562 178634
rect 501646 178398 501882 178634
rect 501326 142718 501562 142954
rect 501646 142718 501882 142954
rect 501326 142398 501562 142634
rect 501646 142398 501882 142634
rect 501326 106718 501562 106954
rect 501646 106718 501882 106954
rect 501326 106398 501562 106634
rect 501646 106398 501882 106634
rect 501326 70718 501562 70954
rect 501646 70718 501882 70954
rect 501326 70398 501562 70634
rect 501646 70398 501882 70634
rect 501326 34718 501562 34954
rect 501646 34718 501882 34954
rect 501326 34398 501562 34634
rect 501646 34398 501882 34634
rect 501326 -7302 501562 -7066
rect 501646 -7302 501882 -7066
rect 501326 -7622 501562 -7386
rect 501646 -7622 501882 -7386
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 510326 705562 510562 705798
rect 510646 705562 510882 705798
rect 510326 705242 510562 705478
rect 510646 705242 510882 705478
rect 510326 691718 510562 691954
rect 510646 691718 510882 691954
rect 510326 691398 510562 691634
rect 510646 691398 510882 691634
rect 510326 655718 510562 655954
rect 510646 655718 510882 655954
rect 510326 655398 510562 655634
rect 510646 655398 510882 655634
rect 510326 619718 510562 619954
rect 510646 619718 510882 619954
rect 510326 619398 510562 619634
rect 510646 619398 510882 619634
rect 510326 583718 510562 583954
rect 510646 583718 510882 583954
rect 510326 583398 510562 583634
rect 510646 583398 510882 583634
rect 510326 547718 510562 547954
rect 510646 547718 510882 547954
rect 510326 547398 510562 547634
rect 510646 547398 510882 547634
rect 510326 511718 510562 511954
rect 510646 511718 510882 511954
rect 510326 511398 510562 511634
rect 510646 511398 510882 511634
rect 510326 475718 510562 475954
rect 510646 475718 510882 475954
rect 510326 475398 510562 475634
rect 510646 475398 510882 475634
rect 510326 439718 510562 439954
rect 510646 439718 510882 439954
rect 510326 439398 510562 439634
rect 510646 439398 510882 439634
rect 510326 403718 510562 403954
rect 510646 403718 510882 403954
rect 510326 403398 510562 403634
rect 510646 403398 510882 403634
rect 510326 367718 510562 367954
rect 510646 367718 510882 367954
rect 510326 367398 510562 367634
rect 510646 367398 510882 367634
rect 510326 331718 510562 331954
rect 510646 331718 510882 331954
rect 510326 331398 510562 331634
rect 510646 331398 510882 331634
rect 510326 295718 510562 295954
rect 510646 295718 510882 295954
rect 510326 295398 510562 295634
rect 510646 295398 510882 295634
rect 510326 259718 510562 259954
rect 510646 259718 510882 259954
rect 510326 259398 510562 259634
rect 510646 259398 510882 259634
rect 510326 223718 510562 223954
rect 510646 223718 510882 223954
rect 510326 223398 510562 223634
rect 510646 223398 510882 223634
rect 510326 187718 510562 187954
rect 510646 187718 510882 187954
rect 510326 187398 510562 187634
rect 510646 187398 510882 187634
rect 510326 151718 510562 151954
rect 510646 151718 510882 151954
rect 510326 151398 510562 151634
rect 510646 151398 510882 151634
rect 510326 115718 510562 115954
rect 510646 115718 510882 115954
rect 510326 115398 510562 115634
rect 510646 115398 510882 115634
rect 510326 79718 510562 79954
rect 510646 79718 510882 79954
rect 510326 79398 510562 79634
rect 510646 79398 510882 79634
rect 510326 43718 510562 43954
rect 510646 43718 510882 43954
rect 510326 43398 510562 43634
rect 510646 43398 510882 43634
rect 510326 7718 510562 7954
rect 510646 7718 510882 7954
rect 510326 7398 510562 7634
rect 510646 7398 510882 7634
rect 510326 -1542 510562 -1306
rect 510646 -1542 510882 -1306
rect 510326 -1862 510562 -1626
rect 510646 -1862 510882 -1626
rect 514826 706522 515062 706758
rect 515146 706522 515382 706758
rect 514826 706202 515062 706438
rect 515146 706202 515382 706438
rect 514826 696218 515062 696454
rect 515146 696218 515382 696454
rect 514826 695898 515062 696134
rect 515146 695898 515382 696134
rect 514826 660218 515062 660454
rect 515146 660218 515382 660454
rect 514826 659898 515062 660134
rect 515146 659898 515382 660134
rect 514826 624218 515062 624454
rect 515146 624218 515382 624454
rect 514826 623898 515062 624134
rect 515146 623898 515382 624134
rect 514826 588218 515062 588454
rect 515146 588218 515382 588454
rect 514826 587898 515062 588134
rect 515146 587898 515382 588134
rect 514826 552218 515062 552454
rect 515146 552218 515382 552454
rect 514826 551898 515062 552134
rect 515146 551898 515382 552134
rect 514826 516218 515062 516454
rect 515146 516218 515382 516454
rect 514826 515898 515062 516134
rect 515146 515898 515382 516134
rect 514826 480218 515062 480454
rect 515146 480218 515382 480454
rect 514826 479898 515062 480134
rect 515146 479898 515382 480134
rect 514826 444218 515062 444454
rect 515146 444218 515382 444454
rect 514826 443898 515062 444134
rect 515146 443898 515382 444134
rect 514826 408218 515062 408454
rect 515146 408218 515382 408454
rect 514826 407898 515062 408134
rect 515146 407898 515382 408134
rect 514826 372218 515062 372454
rect 515146 372218 515382 372454
rect 514826 371898 515062 372134
rect 515146 371898 515382 372134
rect 514826 336218 515062 336454
rect 515146 336218 515382 336454
rect 514826 335898 515062 336134
rect 515146 335898 515382 336134
rect 514826 300218 515062 300454
rect 515146 300218 515382 300454
rect 514826 299898 515062 300134
rect 515146 299898 515382 300134
rect 514826 264218 515062 264454
rect 515146 264218 515382 264454
rect 514826 263898 515062 264134
rect 515146 263898 515382 264134
rect 514826 228218 515062 228454
rect 515146 228218 515382 228454
rect 514826 227898 515062 228134
rect 515146 227898 515382 228134
rect 514826 192218 515062 192454
rect 515146 192218 515382 192454
rect 514826 191898 515062 192134
rect 515146 191898 515382 192134
rect 514826 156218 515062 156454
rect 515146 156218 515382 156454
rect 514826 155898 515062 156134
rect 515146 155898 515382 156134
rect 514826 120218 515062 120454
rect 515146 120218 515382 120454
rect 514826 119898 515062 120134
rect 515146 119898 515382 120134
rect 514826 84218 515062 84454
rect 515146 84218 515382 84454
rect 514826 83898 515062 84134
rect 515146 83898 515382 84134
rect 514826 48218 515062 48454
rect 515146 48218 515382 48454
rect 514826 47898 515062 48134
rect 515146 47898 515382 48134
rect 514826 12218 515062 12454
rect 515146 12218 515382 12454
rect 514826 11898 515062 12134
rect 515146 11898 515382 12134
rect 514826 -2502 515062 -2266
rect 515146 -2502 515382 -2266
rect 514826 -2822 515062 -2586
rect 515146 -2822 515382 -2586
rect 519326 707482 519562 707718
rect 519646 707482 519882 707718
rect 519326 707162 519562 707398
rect 519646 707162 519882 707398
rect 519326 700718 519562 700954
rect 519646 700718 519882 700954
rect 519326 700398 519562 700634
rect 519646 700398 519882 700634
rect 519326 664718 519562 664954
rect 519646 664718 519882 664954
rect 519326 664398 519562 664634
rect 519646 664398 519882 664634
rect 519326 628718 519562 628954
rect 519646 628718 519882 628954
rect 519326 628398 519562 628634
rect 519646 628398 519882 628634
rect 519326 592718 519562 592954
rect 519646 592718 519882 592954
rect 519326 592398 519562 592634
rect 519646 592398 519882 592634
rect 519326 556718 519562 556954
rect 519646 556718 519882 556954
rect 519326 556398 519562 556634
rect 519646 556398 519882 556634
rect 519326 520718 519562 520954
rect 519646 520718 519882 520954
rect 519326 520398 519562 520634
rect 519646 520398 519882 520634
rect 519326 484718 519562 484954
rect 519646 484718 519882 484954
rect 519326 484398 519562 484634
rect 519646 484398 519882 484634
rect 519326 448718 519562 448954
rect 519646 448718 519882 448954
rect 519326 448398 519562 448634
rect 519646 448398 519882 448634
rect 519326 412718 519562 412954
rect 519646 412718 519882 412954
rect 519326 412398 519562 412634
rect 519646 412398 519882 412634
rect 519326 376718 519562 376954
rect 519646 376718 519882 376954
rect 519326 376398 519562 376634
rect 519646 376398 519882 376634
rect 519326 340718 519562 340954
rect 519646 340718 519882 340954
rect 519326 340398 519562 340634
rect 519646 340398 519882 340634
rect 519326 304718 519562 304954
rect 519646 304718 519882 304954
rect 519326 304398 519562 304634
rect 519646 304398 519882 304634
rect 519326 268718 519562 268954
rect 519646 268718 519882 268954
rect 519326 268398 519562 268634
rect 519646 268398 519882 268634
rect 519326 232718 519562 232954
rect 519646 232718 519882 232954
rect 519326 232398 519562 232634
rect 519646 232398 519882 232634
rect 519326 196718 519562 196954
rect 519646 196718 519882 196954
rect 519326 196398 519562 196634
rect 519646 196398 519882 196634
rect 519326 160718 519562 160954
rect 519646 160718 519882 160954
rect 519326 160398 519562 160634
rect 519646 160398 519882 160634
rect 519326 124718 519562 124954
rect 519646 124718 519882 124954
rect 519326 124398 519562 124634
rect 519646 124398 519882 124634
rect 519326 88718 519562 88954
rect 519646 88718 519882 88954
rect 519326 88398 519562 88634
rect 519646 88398 519882 88634
rect 519326 52718 519562 52954
rect 519646 52718 519882 52954
rect 519326 52398 519562 52634
rect 519646 52398 519882 52634
rect 519326 16718 519562 16954
rect 519646 16718 519882 16954
rect 519326 16398 519562 16634
rect 519646 16398 519882 16634
rect 519326 -3462 519562 -3226
rect 519646 -3462 519882 -3226
rect 519326 -3782 519562 -3546
rect 519646 -3782 519882 -3546
rect 523826 708442 524062 708678
rect 524146 708442 524382 708678
rect 523826 708122 524062 708358
rect 524146 708122 524382 708358
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -4422 524062 -4186
rect 524146 -4422 524382 -4186
rect 523826 -4742 524062 -4506
rect 524146 -4742 524382 -4506
rect 528326 709402 528562 709638
rect 528646 709402 528882 709638
rect 528326 709082 528562 709318
rect 528646 709082 528882 709318
rect 528326 673718 528562 673954
rect 528646 673718 528882 673954
rect 528326 673398 528562 673634
rect 528646 673398 528882 673634
rect 528326 637718 528562 637954
rect 528646 637718 528882 637954
rect 528326 637398 528562 637634
rect 528646 637398 528882 637634
rect 528326 601718 528562 601954
rect 528646 601718 528882 601954
rect 528326 601398 528562 601634
rect 528646 601398 528882 601634
rect 528326 565718 528562 565954
rect 528646 565718 528882 565954
rect 528326 565398 528562 565634
rect 528646 565398 528882 565634
rect 528326 529718 528562 529954
rect 528646 529718 528882 529954
rect 528326 529398 528562 529634
rect 528646 529398 528882 529634
rect 528326 493718 528562 493954
rect 528646 493718 528882 493954
rect 528326 493398 528562 493634
rect 528646 493398 528882 493634
rect 528326 457718 528562 457954
rect 528646 457718 528882 457954
rect 528326 457398 528562 457634
rect 528646 457398 528882 457634
rect 528326 421718 528562 421954
rect 528646 421718 528882 421954
rect 528326 421398 528562 421634
rect 528646 421398 528882 421634
rect 528326 385718 528562 385954
rect 528646 385718 528882 385954
rect 528326 385398 528562 385634
rect 528646 385398 528882 385634
rect 528326 349718 528562 349954
rect 528646 349718 528882 349954
rect 528326 349398 528562 349634
rect 528646 349398 528882 349634
rect 528326 313718 528562 313954
rect 528646 313718 528882 313954
rect 528326 313398 528562 313634
rect 528646 313398 528882 313634
rect 528326 277718 528562 277954
rect 528646 277718 528882 277954
rect 528326 277398 528562 277634
rect 528646 277398 528882 277634
rect 528326 241718 528562 241954
rect 528646 241718 528882 241954
rect 528326 241398 528562 241634
rect 528646 241398 528882 241634
rect 528326 205718 528562 205954
rect 528646 205718 528882 205954
rect 528326 205398 528562 205634
rect 528646 205398 528882 205634
rect 528326 169718 528562 169954
rect 528646 169718 528882 169954
rect 528326 169398 528562 169634
rect 528646 169398 528882 169634
rect 528326 133718 528562 133954
rect 528646 133718 528882 133954
rect 528326 133398 528562 133634
rect 528646 133398 528882 133634
rect 528326 97718 528562 97954
rect 528646 97718 528882 97954
rect 528326 97398 528562 97634
rect 528646 97398 528882 97634
rect 528326 61718 528562 61954
rect 528646 61718 528882 61954
rect 528326 61398 528562 61634
rect 528646 61398 528882 61634
rect 528326 25718 528562 25954
rect 528646 25718 528882 25954
rect 528326 25398 528562 25634
rect 528646 25398 528882 25634
rect 528326 -5382 528562 -5146
rect 528646 -5382 528882 -5146
rect 528326 -5702 528562 -5466
rect 528646 -5702 528882 -5466
rect 532826 710362 533062 710598
rect 533146 710362 533382 710598
rect 532826 710042 533062 710278
rect 533146 710042 533382 710278
rect 532826 678218 533062 678454
rect 533146 678218 533382 678454
rect 532826 677898 533062 678134
rect 533146 677898 533382 678134
rect 532826 642218 533062 642454
rect 533146 642218 533382 642454
rect 532826 641898 533062 642134
rect 533146 641898 533382 642134
rect 532826 606218 533062 606454
rect 533146 606218 533382 606454
rect 532826 605898 533062 606134
rect 533146 605898 533382 606134
rect 532826 570218 533062 570454
rect 533146 570218 533382 570454
rect 532826 569898 533062 570134
rect 533146 569898 533382 570134
rect 532826 534218 533062 534454
rect 533146 534218 533382 534454
rect 532826 533898 533062 534134
rect 533146 533898 533382 534134
rect 532826 498218 533062 498454
rect 533146 498218 533382 498454
rect 532826 497898 533062 498134
rect 533146 497898 533382 498134
rect 532826 462218 533062 462454
rect 533146 462218 533382 462454
rect 532826 461898 533062 462134
rect 533146 461898 533382 462134
rect 532826 426218 533062 426454
rect 533146 426218 533382 426454
rect 532826 425898 533062 426134
rect 533146 425898 533382 426134
rect 532826 390218 533062 390454
rect 533146 390218 533382 390454
rect 532826 389898 533062 390134
rect 533146 389898 533382 390134
rect 532826 354218 533062 354454
rect 533146 354218 533382 354454
rect 532826 353898 533062 354134
rect 533146 353898 533382 354134
rect 532826 318218 533062 318454
rect 533146 318218 533382 318454
rect 532826 317898 533062 318134
rect 533146 317898 533382 318134
rect 532826 282218 533062 282454
rect 533146 282218 533382 282454
rect 532826 281898 533062 282134
rect 533146 281898 533382 282134
rect 532826 246218 533062 246454
rect 533146 246218 533382 246454
rect 532826 245898 533062 246134
rect 533146 245898 533382 246134
rect 532826 210218 533062 210454
rect 533146 210218 533382 210454
rect 532826 209898 533062 210134
rect 533146 209898 533382 210134
rect 532826 174218 533062 174454
rect 533146 174218 533382 174454
rect 532826 173898 533062 174134
rect 533146 173898 533382 174134
rect 532826 138218 533062 138454
rect 533146 138218 533382 138454
rect 532826 137898 533062 138134
rect 533146 137898 533382 138134
rect 532826 102218 533062 102454
rect 533146 102218 533382 102454
rect 532826 101898 533062 102134
rect 533146 101898 533382 102134
rect 532826 66218 533062 66454
rect 533146 66218 533382 66454
rect 532826 65898 533062 66134
rect 533146 65898 533382 66134
rect 532826 30218 533062 30454
rect 533146 30218 533382 30454
rect 532826 29898 533062 30134
rect 533146 29898 533382 30134
rect 532826 -6342 533062 -6106
rect 533146 -6342 533382 -6106
rect 532826 -6662 533062 -6426
rect 533146 -6662 533382 -6426
rect 537326 711322 537562 711558
rect 537646 711322 537882 711558
rect 537326 711002 537562 711238
rect 537646 711002 537882 711238
rect 537326 682718 537562 682954
rect 537646 682718 537882 682954
rect 537326 682398 537562 682634
rect 537646 682398 537882 682634
rect 537326 646718 537562 646954
rect 537646 646718 537882 646954
rect 537326 646398 537562 646634
rect 537646 646398 537882 646634
rect 537326 610718 537562 610954
rect 537646 610718 537882 610954
rect 537326 610398 537562 610634
rect 537646 610398 537882 610634
rect 537326 574718 537562 574954
rect 537646 574718 537882 574954
rect 537326 574398 537562 574634
rect 537646 574398 537882 574634
rect 537326 538718 537562 538954
rect 537646 538718 537882 538954
rect 537326 538398 537562 538634
rect 537646 538398 537882 538634
rect 537326 502718 537562 502954
rect 537646 502718 537882 502954
rect 537326 502398 537562 502634
rect 537646 502398 537882 502634
rect 537326 466718 537562 466954
rect 537646 466718 537882 466954
rect 537326 466398 537562 466634
rect 537646 466398 537882 466634
rect 537326 430718 537562 430954
rect 537646 430718 537882 430954
rect 537326 430398 537562 430634
rect 537646 430398 537882 430634
rect 537326 394718 537562 394954
rect 537646 394718 537882 394954
rect 537326 394398 537562 394634
rect 537646 394398 537882 394634
rect 537326 358718 537562 358954
rect 537646 358718 537882 358954
rect 537326 358398 537562 358634
rect 537646 358398 537882 358634
rect 537326 322718 537562 322954
rect 537646 322718 537882 322954
rect 537326 322398 537562 322634
rect 537646 322398 537882 322634
rect 537326 286718 537562 286954
rect 537646 286718 537882 286954
rect 537326 286398 537562 286634
rect 537646 286398 537882 286634
rect 537326 250718 537562 250954
rect 537646 250718 537882 250954
rect 537326 250398 537562 250634
rect 537646 250398 537882 250634
rect 537326 214718 537562 214954
rect 537646 214718 537882 214954
rect 537326 214398 537562 214634
rect 537646 214398 537882 214634
rect 537326 178718 537562 178954
rect 537646 178718 537882 178954
rect 537326 178398 537562 178634
rect 537646 178398 537882 178634
rect 537326 142718 537562 142954
rect 537646 142718 537882 142954
rect 537326 142398 537562 142634
rect 537646 142398 537882 142634
rect 537326 106718 537562 106954
rect 537646 106718 537882 106954
rect 537326 106398 537562 106634
rect 537646 106398 537882 106634
rect 537326 70718 537562 70954
rect 537646 70718 537882 70954
rect 537326 70398 537562 70634
rect 537646 70398 537882 70634
rect 537326 34718 537562 34954
rect 537646 34718 537882 34954
rect 537326 34398 537562 34634
rect 537646 34398 537882 34634
rect 537326 -7302 537562 -7066
rect 537646 -7302 537882 -7066
rect 537326 -7622 537562 -7386
rect 537646 -7622 537882 -7386
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 546326 705562 546562 705798
rect 546646 705562 546882 705798
rect 546326 705242 546562 705478
rect 546646 705242 546882 705478
rect 546326 691718 546562 691954
rect 546646 691718 546882 691954
rect 546326 691398 546562 691634
rect 546646 691398 546882 691634
rect 546326 655718 546562 655954
rect 546646 655718 546882 655954
rect 546326 655398 546562 655634
rect 546646 655398 546882 655634
rect 546326 619718 546562 619954
rect 546646 619718 546882 619954
rect 546326 619398 546562 619634
rect 546646 619398 546882 619634
rect 546326 583718 546562 583954
rect 546646 583718 546882 583954
rect 546326 583398 546562 583634
rect 546646 583398 546882 583634
rect 546326 547718 546562 547954
rect 546646 547718 546882 547954
rect 546326 547398 546562 547634
rect 546646 547398 546882 547634
rect 546326 511718 546562 511954
rect 546646 511718 546882 511954
rect 546326 511398 546562 511634
rect 546646 511398 546882 511634
rect 546326 475718 546562 475954
rect 546646 475718 546882 475954
rect 546326 475398 546562 475634
rect 546646 475398 546882 475634
rect 546326 439718 546562 439954
rect 546646 439718 546882 439954
rect 546326 439398 546562 439634
rect 546646 439398 546882 439634
rect 546326 403718 546562 403954
rect 546646 403718 546882 403954
rect 546326 403398 546562 403634
rect 546646 403398 546882 403634
rect 546326 367718 546562 367954
rect 546646 367718 546882 367954
rect 546326 367398 546562 367634
rect 546646 367398 546882 367634
rect 546326 331718 546562 331954
rect 546646 331718 546882 331954
rect 546326 331398 546562 331634
rect 546646 331398 546882 331634
rect 546326 295718 546562 295954
rect 546646 295718 546882 295954
rect 546326 295398 546562 295634
rect 546646 295398 546882 295634
rect 546326 259718 546562 259954
rect 546646 259718 546882 259954
rect 546326 259398 546562 259634
rect 546646 259398 546882 259634
rect 546326 223718 546562 223954
rect 546646 223718 546882 223954
rect 546326 223398 546562 223634
rect 546646 223398 546882 223634
rect 546326 187718 546562 187954
rect 546646 187718 546882 187954
rect 546326 187398 546562 187634
rect 546646 187398 546882 187634
rect 546326 151718 546562 151954
rect 546646 151718 546882 151954
rect 546326 151398 546562 151634
rect 546646 151398 546882 151634
rect 546326 115718 546562 115954
rect 546646 115718 546882 115954
rect 546326 115398 546562 115634
rect 546646 115398 546882 115634
rect 546326 79718 546562 79954
rect 546646 79718 546882 79954
rect 546326 79398 546562 79634
rect 546646 79398 546882 79634
rect 546326 43718 546562 43954
rect 546646 43718 546882 43954
rect 546326 43398 546562 43634
rect 546646 43398 546882 43634
rect 546326 7718 546562 7954
rect 546646 7718 546882 7954
rect 546326 7398 546562 7634
rect 546646 7398 546882 7634
rect 546326 -1542 546562 -1306
rect 546646 -1542 546882 -1306
rect 546326 -1862 546562 -1626
rect 546646 -1862 546882 -1626
rect 550826 706522 551062 706758
rect 551146 706522 551382 706758
rect 550826 706202 551062 706438
rect 551146 706202 551382 706438
rect 550826 696218 551062 696454
rect 551146 696218 551382 696454
rect 550826 695898 551062 696134
rect 551146 695898 551382 696134
rect 550826 660218 551062 660454
rect 551146 660218 551382 660454
rect 550826 659898 551062 660134
rect 551146 659898 551382 660134
rect 550826 624218 551062 624454
rect 551146 624218 551382 624454
rect 550826 623898 551062 624134
rect 551146 623898 551382 624134
rect 550826 588218 551062 588454
rect 551146 588218 551382 588454
rect 550826 587898 551062 588134
rect 551146 587898 551382 588134
rect 550826 552218 551062 552454
rect 551146 552218 551382 552454
rect 550826 551898 551062 552134
rect 551146 551898 551382 552134
rect 550826 516218 551062 516454
rect 551146 516218 551382 516454
rect 550826 515898 551062 516134
rect 551146 515898 551382 516134
rect 550826 480218 551062 480454
rect 551146 480218 551382 480454
rect 550826 479898 551062 480134
rect 551146 479898 551382 480134
rect 550826 444218 551062 444454
rect 551146 444218 551382 444454
rect 550826 443898 551062 444134
rect 551146 443898 551382 444134
rect 550826 408218 551062 408454
rect 551146 408218 551382 408454
rect 550826 407898 551062 408134
rect 551146 407898 551382 408134
rect 550826 372218 551062 372454
rect 551146 372218 551382 372454
rect 550826 371898 551062 372134
rect 551146 371898 551382 372134
rect 550826 336218 551062 336454
rect 551146 336218 551382 336454
rect 550826 335898 551062 336134
rect 551146 335898 551382 336134
rect 550826 300218 551062 300454
rect 551146 300218 551382 300454
rect 550826 299898 551062 300134
rect 551146 299898 551382 300134
rect 550826 264218 551062 264454
rect 551146 264218 551382 264454
rect 550826 263898 551062 264134
rect 551146 263898 551382 264134
rect 550826 228218 551062 228454
rect 551146 228218 551382 228454
rect 550826 227898 551062 228134
rect 551146 227898 551382 228134
rect 550826 192218 551062 192454
rect 551146 192218 551382 192454
rect 550826 191898 551062 192134
rect 551146 191898 551382 192134
rect 550826 156218 551062 156454
rect 551146 156218 551382 156454
rect 550826 155898 551062 156134
rect 551146 155898 551382 156134
rect 550826 120218 551062 120454
rect 551146 120218 551382 120454
rect 550826 119898 551062 120134
rect 551146 119898 551382 120134
rect 550826 84218 551062 84454
rect 551146 84218 551382 84454
rect 550826 83898 551062 84134
rect 551146 83898 551382 84134
rect 550826 48218 551062 48454
rect 551146 48218 551382 48454
rect 550826 47898 551062 48134
rect 551146 47898 551382 48134
rect 550826 12218 551062 12454
rect 551146 12218 551382 12454
rect 550826 11898 551062 12134
rect 551146 11898 551382 12134
rect 550826 -2502 551062 -2266
rect 551146 -2502 551382 -2266
rect 550826 -2822 551062 -2586
rect 551146 -2822 551382 -2586
rect 555326 707482 555562 707718
rect 555646 707482 555882 707718
rect 555326 707162 555562 707398
rect 555646 707162 555882 707398
rect 555326 700718 555562 700954
rect 555646 700718 555882 700954
rect 555326 700398 555562 700634
rect 555646 700398 555882 700634
rect 555326 664718 555562 664954
rect 555646 664718 555882 664954
rect 555326 664398 555562 664634
rect 555646 664398 555882 664634
rect 555326 628718 555562 628954
rect 555646 628718 555882 628954
rect 555326 628398 555562 628634
rect 555646 628398 555882 628634
rect 555326 592718 555562 592954
rect 555646 592718 555882 592954
rect 555326 592398 555562 592634
rect 555646 592398 555882 592634
rect 555326 556718 555562 556954
rect 555646 556718 555882 556954
rect 555326 556398 555562 556634
rect 555646 556398 555882 556634
rect 555326 520718 555562 520954
rect 555646 520718 555882 520954
rect 555326 520398 555562 520634
rect 555646 520398 555882 520634
rect 555326 484718 555562 484954
rect 555646 484718 555882 484954
rect 555326 484398 555562 484634
rect 555646 484398 555882 484634
rect 555326 448718 555562 448954
rect 555646 448718 555882 448954
rect 555326 448398 555562 448634
rect 555646 448398 555882 448634
rect 555326 412718 555562 412954
rect 555646 412718 555882 412954
rect 555326 412398 555562 412634
rect 555646 412398 555882 412634
rect 555326 376718 555562 376954
rect 555646 376718 555882 376954
rect 555326 376398 555562 376634
rect 555646 376398 555882 376634
rect 555326 340718 555562 340954
rect 555646 340718 555882 340954
rect 555326 340398 555562 340634
rect 555646 340398 555882 340634
rect 555326 304718 555562 304954
rect 555646 304718 555882 304954
rect 555326 304398 555562 304634
rect 555646 304398 555882 304634
rect 555326 268718 555562 268954
rect 555646 268718 555882 268954
rect 555326 268398 555562 268634
rect 555646 268398 555882 268634
rect 555326 232718 555562 232954
rect 555646 232718 555882 232954
rect 555326 232398 555562 232634
rect 555646 232398 555882 232634
rect 555326 196718 555562 196954
rect 555646 196718 555882 196954
rect 555326 196398 555562 196634
rect 555646 196398 555882 196634
rect 555326 160718 555562 160954
rect 555646 160718 555882 160954
rect 555326 160398 555562 160634
rect 555646 160398 555882 160634
rect 555326 124718 555562 124954
rect 555646 124718 555882 124954
rect 555326 124398 555562 124634
rect 555646 124398 555882 124634
rect 555326 88718 555562 88954
rect 555646 88718 555882 88954
rect 555326 88398 555562 88634
rect 555646 88398 555882 88634
rect 555326 52718 555562 52954
rect 555646 52718 555882 52954
rect 555326 52398 555562 52634
rect 555646 52398 555882 52634
rect 555326 16718 555562 16954
rect 555646 16718 555882 16954
rect 555326 16398 555562 16634
rect 555646 16398 555882 16634
rect 555326 -3462 555562 -3226
rect 555646 -3462 555882 -3226
rect 555326 -3782 555562 -3546
rect 555646 -3782 555882 -3546
rect 559826 708442 560062 708678
rect 560146 708442 560382 708678
rect 559826 708122 560062 708358
rect 560146 708122 560382 708358
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -4422 560062 -4186
rect 560146 -4422 560382 -4186
rect 559826 -4742 560062 -4506
rect 560146 -4742 560382 -4506
rect 564326 709402 564562 709638
rect 564646 709402 564882 709638
rect 564326 709082 564562 709318
rect 564646 709082 564882 709318
rect 564326 673718 564562 673954
rect 564646 673718 564882 673954
rect 564326 673398 564562 673634
rect 564646 673398 564882 673634
rect 564326 637718 564562 637954
rect 564646 637718 564882 637954
rect 564326 637398 564562 637634
rect 564646 637398 564882 637634
rect 564326 601718 564562 601954
rect 564646 601718 564882 601954
rect 564326 601398 564562 601634
rect 564646 601398 564882 601634
rect 564326 565718 564562 565954
rect 564646 565718 564882 565954
rect 564326 565398 564562 565634
rect 564646 565398 564882 565634
rect 564326 529718 564562 529954
rect 564646 529718 564882 529954
rect 564326 529398 564562 529634
rect 564646 529398 564882 529634
rect 564326 493718 564562 493954
rect 564646 493718 564882 493954
rect 564326 493398 564562 493634
rect 564646 493398 564882 493634
rect 564326 457718 564562 457954
rect 564646 457718 564882 457954
rect 564326 457398 564562 457634
rect 564646 457398 564882 457634
rect 564326 421718 564562 421954
rect 564646 421718 564882 421954
rect 564326 421398 564562 421634
rect 564646 421398 564882 421634
rect 564326 385718 564562 385954
rect 564646 385718 564882 385954
rect 564326 385398 564562 385634
rect 564646 385398 564882 385634
rect 564326 349718 564562 349954
rect 564646 349718 564882 349954
rect 564326 349398 564562 349634
rect 564646 349398 564882 349634
rect 564326 313718 564562 313954
rect 564646 313718 564882 313954
rect 564326 313398 564562 313634
rect 564646 313398 564882 313634
rect 564326 277718 564562 277954
rect 564646 277718 564882 277954
rect 564326 277398 564562 277634
rect 564646 277398 564882 277634
rect 564326 241718 564562 241954
rect 564646 241718 564882 241954
rect 564326 241398 564562 241634
rect 564646 241398 564882 241634
rect 564326 205718 564562 205954
rect 564646 205718 564882 205954
rect 564326 205398 564562 205634
rect 564646 205398 564882 205634
rect 564326 169718 564562 169954
rect 564646 169718 564882 169954
rect 564326 169398 564562 169634
rect 564646 169398 564882 169634
rect 564326 133718 564562 133954
rect 564646 133718 564882 133954
rect 564326 133398 564562 133634
rect 564646 133398 564882 133634
rect 564326 97718 564562 97954
rect 564646 97718 564882 97954
rect 564326 97398 564562 97634
rect 564646 97398 564882 97634
rect 564326 61718 564562 61954
rect 564646 61718 564882 61954
rect 564326 61398 564562 61634
rect 564646 61398 564882 61634
rect 564326 25718 564562 25954
rect 564646 25718 564882 25954
rect 564326 25398 564562 25634
rect 564646 25398 564882 25634
rect 564326 -5382 564562 -5146
rect 564646 -5382 564882 -5146
rect 564326 -5702 564562 -5466
rect 564646 -5702 564882 -5466
rect 568826 710362 569062 710598
rect 569146 710362 569382 710598
rect 568826 710042 569062 710278
rect 569146 710042 569382 710278
rect 568826 678218 569062 678454
rect 569146 678218 569382 678454
rect 568826 677898 569062 678134
rect 569146 677898 569382 678134
rect 568826 642218 569062 642454
rect 569146 642218 569382 642454
rect 568826 641898 569062 642134
rect 569146 641898 569382 642134
rect 568826 606218 569062 606454
rect 569146 606218 569382 606454
rect 568826 605898 569062 606134
rect 569146 605898 569382 606134
rect 568826 570218 569062 570454
rect 569146 570218 569382 570454
rect 568826 569898 569062 570134
rect 569146 569898 569382 570134
rect 568826 534218 569062 534454
rect 569146 534218 569382 534454
rect 568826 533898 569062 534134
rect 569146 533898 569382 534134
rect 568826 498218 569062 498454
rect 569146 498218 569382 498454
rect 568826 497898 569062 498134
rect 569146 497898 569382 498134
rect 568826 462218 569062 462454
rect 569146 462218 569382 462454
rect 568826 461898 569062 462134
rect 569146 461898 569382 462134
rect 568826 426218 569062 426454
rect 569146 426218 569382 426454
rect 568826 425898 569062 426134
rect 569146 425898 569382 426134
rect 568826 390218 569062 390454
rect 569146 390218 569382 390454
rect 568826 389898 569062 390134
rect 569146 389898 569382 390134
rect 568826 354218 569062 354454
rect 569146 354218 569382 354454
rect 568826 353898 569062 354134
rect 569146 353898 569382 354134
rect 568826 318218 569062 318454
rect 569146 318218 569382 318454
rect 568826 317898 569062 318134
rect 569146 317898 569382 318134
rect 568826 282218 569062 282454
rect 569146 282218 569382 282454
rect 568826 281898 569062 282134
rect 569146 281898 569382 282134
rect 568826 246218 569062 246454
rect 569146 246218 569382 246454
rect 568826 245898 569062 246134
rect 569146 245898 569382 246134
rect 568826 210218 569062 210454
rect 569146 210218 569382 210454
rect 568826 209898 569062 210134
rect 569146 209898 569382 210134
rect 568826 174218 569062 174454
rect 569146 174218 569382 174454
rect 568826 173898 569062 174134
rect 569146 173898 569382 174134
rect 568826 138218 569062 138454
rect 569146 138218 569382 138454
rect 568826 137898 569062 138134
rect 569146 137898 569382 138134
rect 568826 102218 569062 102454
rect 569146 102218 569382 102454
rect 568826 101898 569062 102134
rect 569146 101898 569382 102134
rect 568826 66218 569062 66454
rect 569146 66218 569382 66454
rect 568826 65898 569062 66134
rect 569146 65898 569382 66134
rect 568826 30218 569062 30454
rect 569146 30218 569382 30454
rect 568826 29898 569062 30134
rect 569146 29898 569382 30134
rect 568826 -6342 569062 -6106
rect 569146 -6342 569382 -6106
rect 568826 -6662 569062 -6426
rect 569146 -6662 569382 -6426
rect 573326 711322 573562 711558
rect 573646 711322 573882 711558
rect 573326 711002 573562 711238
rect 573646 711002 573882 711238
rect 573326 682718 573562 682954
rect 573646 682718 573882 682954
rect 573326 682398 573562 682634
rect 573646 682398 573882 682634
rect 573326 646718 573562 646954
rect 573646 646718 573882 646954
rect 573326 646398 573562 646634
rect 573646 646398 573882 646634
rect 573326 610718 573562 610954
rect 573646 610718 573882 610954
rect 573326 610398 573562 610634
rect 573646 610398 573882 610634
rect 573326 574718 573562 574954
rect 573646 574718 573882 574954
rect 573326 574398 573562 574634
rect 573646 574398 573882 574634
rect 573326 538718 573562 538954
rect 573646 538718 573882 538954
rect 573326 538398 573562 538634
rect 573646 538398 573882 538634
rect 573326 502718 573562 502954
rect 573646 502718 573882 502954
rect 573326 502398 573562 502634
rect 573646 502398 573882 502634
rect 573326 466718 573562 466954
rect 573646 466718 573882 466954
rect 573326 466398 573562 466634
rect 573646 466398 573882 466634
rect 573326 430718 573562 430954
rect 573646 430718 573882 430954
rect 573326 430398 573562 430634
rect 573646 430398 573882 430634
rect 573326 394718 573562 394954
rect 573646 394718 573882 394954
rect 573326 394398 573562 394634
rect 573646 394398 573882 394634
rect 573326 358718 573562 358954
rect 573646 358718 573882 358954
rect 573326 358398 573562 358634
rect 573646 358398 573882 358634
rect 573326 322718 573562 322954
rect 573646 322718 573882 322954
rect 573326 322398 573562 322634
rect 573646 322398 573882 322634
rect 573326 286718 573562 286954
rect 573646 286718 573882 286954
rect 573326 286398 573562 286634
rect 573646 286398 573882 286634
rect 573326 250718 573562 250954
rect 573646 250718 573882 250954
rect 573326 250398 573562 250634
rect 573646 250398 573882 250634
rect 573326 214718 573562 214954
rect 573646 214718 573882 214954
rect 573326 214398 573562 214634
rect 573646 214398 573882 214634
rect 573326 178718 573562 178954
rect 573646 178718 573882 178954
rect 573326 178398 573562 178634
rect 573646 178398 573882 178634
rect 573326 142718 573562 142954
rect 573646 142718 573882 142954
rect 573326 142398 573562 142634
rect 573646 142398 573882 142634
rect 573326 106718 573562 106954
rect 573646 106718 573882 106954
rect 573326 106398 573562 106634
rect 573646 106398 573882 106634
rect 573326 70718 573562 70954
rect 573646 70718 573882 70954
rect 573326 70398 573562 70634
rect 573646 70398 573882 70634
rect 573326 34718 573562 34954
rect 573646 34718 573882 34954
rect 573326 34398 573562 34634
rect 573646 34398 573882 34634
rect 573326 -7302 573562 -7066
rect 573646 -7302 573882 -7066
rect 573326 -7622 573562 -7386
rect 573646 -7622 573882 -7386
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 582326 705562 582562 705798
rect 582646 705562 582882 705798
rect 582326 705242 582562 705478
rect 582646 705242 582882 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 582326 691718 582562 691954
rect 582646 691718 582882 691954
rect 582326 691398 582562 691634
rect 582646 691398 582882 691634
rect 582326 655718 582562 655954
rect 582646 655718 582882 655954
rect 582326 655398 582562 655634
rect 582646 655398 582882 655634
rect 582326 619718 582562 619954
rect 582646 619718 582882 619954
rect 582326 619398 582562 619634
rect 582646 619398 582882 619634
rect 582326 583718 582562 583954
rect 582646 583718 582882 583954
rect 582326 583398 582562 583634
rect 582646 583398 582882 583634
rect 582326 547718 582562 547954
rect 582646 547718 582882 547954
rect 582326 547398 582562 547634
rect 582646 547398 582882 547634
rect 582326 511718 582562 511954
rect 582646 511718 582882 511954
rect 582326 511398 582562 511634
rect 582646 511398 582882 511634
rect 582326 475718 582562 475954
rect 582646 475718 582882 475954
rect 582326 475398 582562 475634
rect 582646 475398 582882 475634
rect 582326 439718 582562 439954
rect 582646 439718 582882 439954
rect 582326 439398 582562 439634
rect 582646 439398 582882 439634
rect 582326 403718 582562 403954
rect 582646 403718 582882 403954
rect 582326 403398 582562 403634
rect 582646 403398 582882 403634
rect 582326 367718 582562 367954
rect 582646 367718 582882 367954
rect 582326 367398 582562 367634
rect 582646 367398 582882 367634
rect 582326 331718 582562 331954
rect 582646 331718 582882 331954
rect 582326 331398 582562 331634
rect 582646 331398 582882 331634
rect 582326 295718 582562 295954
rect 582646 295718 582882 295954
rect 582326 295398 582562 295634
rect 582646 295398 582882 295634
rect 582326 259718 582562 259954
rect 582646 259718 582882 259954
rect 582326 259398 582562 259634
rect 582646 259398 582882 259634
rect 582326 223718 582562 223954
rect 582646 223718 582882 223954
rect 582326 223398 582562 223634
rect 582646 223398 582882 223634
rect 582326 187718 582562 187954
rect 582646 187718 582882 187954
rect 582326 187398 582562 187634
rect 582646 187398 582882 187634
rect 582326 151718 582562 151954
rect 582646 151718 582882 151954
rect 582326 151398 582562 151634
rect 582646 151398 582882 151634
rect 582326 115718 582562 115954
rect 582646 115718 582882 115954
rect 582326 115398 582562 115634
rect 582646 115398 582882 115634
rect 582326 79718 582562 79954
rect 582646 79718 582882 79954
rect 582326 79398 582562 79634
rect 582646 79398 582882 79634
rect 582326 43718 582562 43954
rect 582646 43718 582882 43954
rect 582326 43398 582562 43634
rect 582646 43398 582882 43634
rect 582326 7718 582562 7954
rect 582646 7718 582882 7954
rect 582326 7398 582562 7634
rect 582646 7398 582882 7634
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 691718 586538 691954
rect 586622 691718 586858 691954
rect 586302 691398 586538 691634
rect 586622 691398 586858 691634
rect 586302 655718 586538 655954
rect 586622 655718 586858 655954
rect 586302 655398 586538 655634
rect 586622 655398 586858 655634
rect 586302 619718 586538 619954
rect 586622 619718 586858 619954
rect 586302 619398 586538 619634
rect 586622 619398 586858 619634
rect 586302 583718 586538 583954
rect 586622 583718 586858 583954
rect 586302 583398 586538 583634
rect 586622 583398 586858 583634
rect 586302 547718 586538 547954
rect 586622 547718 586858 547954
rect 586302 547398 586538 547634
rect 586622 547398 586858 547634
rect 586302 511718 586538 511954
rect 586622 511718 586858 511954
rect 586302 511398 586538 511634
rect 586622 511398 586858 511634
rect 586302 475718 586538 475954
rect 586622 475718 586858 475954
rect 586302 475398 586538 475634
rect 586622 475398 586858 475634
rect 586302 439718 586538 439954
rect 586622 439718 586858 439954
rect 586302 439398 586538 439634
rect 586622 439398 586858 439634
rect 586302 403718 586538 403954
rect 586622 403718 586858 403954
rect 586302 403398 586538 403634
rect 586622 403398 586858 403634
rect 586302 367718 586538 367954
rect 586622 367718 586858 367954
rect 586302 367398 586538 367634
rect 586622 367398 586858 367634
rect 586302 331718 586538 331954
rect 586622 331718 586858 331954
rect 586302 331398 586538 331634
rect 586622 331398 586858 331634
rect 586302 295718 586538 295954
rect 586622 295718 586858 295954
rect 586302 295398 586538 295634
rect 586622 295398 586858 295634
rect 586302 259718 586538 259954
rect 586622 259718 586858 259954
rect 586302 259398 586538 259634
rect 586622 259398 586858 259634
rect 586302 223718 586538 223954
rect 586622 223718 586858 223954
rect 586302 223398 586538 223634
rect 586622 223398 586858 223634
rect 586302 187718 586538 187954
rect 586622 187718 586858 187954
rect 586302 187398 586538 187634
rect 586622 187398 586858 187634
rect 586302 151718 586538 151954
rect 586622 151718 586858 151954
rect 586302 151398 586538 151634
rect 586622 151398 586858 151634
rect 586302 115718 586538 115954
rect 586622 115718 586858 115954
rect 586302 115398 586538 115634
rect 586622 115398 586858 115634
rect 586302 79718 586538 79954
rect 586622 79718 586858 79954
rect 586302 79398 586538 79634
rect 586622 79398 586858 79634
rect 586302 43718 586538 43954
rect 586622 43718 586858 43954
rect 586302 43398 586538 43634
rect 586622 43398 586858 43634
rect 586302 7718 586538 7954
rect 586622 7718 586858 7954
rect 586302 7398 586538 7634
rect 586622 7398 586858 7634
rect 582326 -1542 582562 -1306
rect 582646 -1542 582882 -1306
rect 582326 -1862 582562 -1626
rect 582646 -1862 582882 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 696218 587498 696454
rect 587582 696218 587818 696454
rect 587262 695898 587498 696134
rect 587582 695898 587818 696134
rect 587262 660218 587498 660454
rect 587582 660218 587818 660454
rect 587262 659898 587498 660134
rect 587582 659898 587818 660134
rect 587262 624218 587498 624454
rect 587582 624218 587818 624454
rect 587262 623898 587498 624134
rect 587582 623898 587818 624134
rect 587262 588218 587498 588454
rect 587582 588218 587818 588454
rect 587262 587898 587498 588134
rect 587582 587898 587818 588134
rect 587262 552218 587498 552454
rect 587582 552218 587818 552454
rect 587262 551898 587498 552134
rect 587582 551898 587818 552134
rect 587262 516218 587498 516454
rect 587582 516218 587818 516454
rect 587262 515898 587498 516134
rect 587582 515898 587818 516134
rect 587262 480218 587498 480454
rect 587582 480218 587818 480454
rect 587262 479898 587498 480134
rect 587582 479898 587818 480134
rect 587262 444218 587498 444454
rect 587582 444218 587818 444454
rect 587262 443898 587498 444134
rect 587582 443898 587818 444134
rect 587262 408218 587498 408454
rect 587582 408218 587818 408454
rect 587262 407898 587498 408134
rect 587582 407898 587818 408134
rect 587262 372218 587498 372454
rect 587582 372218 587818 372454
rect 587262 371898 587498 372134
rect 587582 371898 587818 372134
rect 587262 336218 587498 336454
rect 587582 336218 587818 336454
rect 587262 335898 587498 336134
rect 587582 335898 587818 336134
rect 587262 300218 587498 300454
rect 587582 300218 587818 300454
rect 587262 299898 587498 300134
rect 587582 299898 587818 300134
rect 587262 264218 587498 264454
rect 587582 264218 587818 264454
rect 587262 263898 587498 264134
rect 587582 263898 587818 264134
rect 587262 228218 587498 228454
rect 587582 228218 587818 228454
rect 587262 227898 587498 228134
rect 587582 227898 587818 228134
rect 587262 192218 587498 192454
rect 587582 192218 587818 192454
rect 587262 191898 587498 192134
rect 587582 191898 587818 192134
rect 587262 156218 587498 156454
rect 587582 156218 587818 156454
rect 587262 155898 587498 156134
rect 587582 155898 587818 156134
rect 587262 120218 587498 120454
rect 587582 120218 587818 120454
rect 587262 119898 587498 120134
rect 587582 119898 587818 120134
rect 587262 84218 587498 84454
rect 587582 84218 587818 84454
rect 587262 83898 587498 84134
rect 587582 83898 587818 84134
rect 587262 48218 587498 48454
rect 587582 48218 587818 48454
rect 587262 47898 587498 48134
rect 587582 47898 587818 48134
rect 587262 12218 587498 12454
rect 587582 12218 587818 12454
rect 587262 11898 587498 12134
rect 587582 11898 587818 12134
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 700718 588458 700954
rect 588542 700718 588778 700954
rect 588222 700398 588458 700634
rect 588542 700398 588778 700634
rect 588222 664718 588458 664954
rect 588542 664718 588778 664954
rect 588222 664398 588458 664634
rect 588542 664398 588778 664634
rect 588222 628718 588458 628954
rect 588542 628718 588778 628954
rect 588222 628398 588458 628634
rect 588542 628398 588778 628634
rect 588222 592718 588458 592954
rect 588542 592718 588778 592954
rect 588222 592398 588458 592634
rect 588542 592398 588778 592634
rect 588222 556718 588458 556954
rect 588542 556718 588778 556954
rect 588222 556398 588458 556634
rect 588542 556398 588778 556634
rect 588222 520718 588458 520954
rect 588542 520718 588778 520954
rect 588222 520398 588458 520634
rect 588542 520398 588778 520634
rect 588222 484718 588458 484954
rect 588542 484718 588778 484954
rect 588222 484398 588458 484634
rect 588542 484398 588778 484634
rect 588222 448718 588458 448954
rect 588542 448718 588778 448954
rect 588222 448398 588458 448634
rect 588542 448398 588778 448634
rect 588222 412718 588458 412954
rect 588542 412718 588778 412954
rect 588222 412398 588458 412634
rect 588542 412398 588778 412634
rect 588222 376718 588458 376954
rect 588542 376718 588778 376954
rect 588222 376398 588458 376634
rect 588542 376398 588778 376634
rect 588222 340718 588458 340954
rect 588542 340718 588778 340954
rect 588222 340398 588458 340634
rect 588542 340398 588778 340634
rect 588222 304718 588458 304954
rect 588542 304718 588778 304954
rect 588222 304398 588458 304634
rect 588542 304398 588778 304634
rect 588222 268718 588458 268954
rect 588542 268718 588778 268954
rect 588222 268398 588458 268634
rect 588542 268398 588778 268634
rect 588222 232718 588458 232954
rect 588542 232718 588778 232954
rect 588222 232398 588458 232634
rect 588542 232398 588778 232634
rect 588222 196718 588458 196954
rect 588542 196718 588778 196954
rect 588222 196398 588458 196634
rect 588542 196398 588778 196634
rect 588222 160718 588458 160954
rect 588542 160718 588778 160954
rect 588222 160398 588458 160634
rect 588542 160398 588778 160634
rect 588222 124718 588458 124954
rect 588542 124718 588778 124954
rect 588222 124398 588458 124634
rect 588542 124398 588778 124634
rect 588222 88718 588458 88954
rect 588542 88718 588778 88954
rect 588222 88398 588458 88634
rect 588542 88398 588778 88634
rect 588222 52718 588458 52954
rect 588542 52718 588778 52954
rect 588222 52398 588458 52634
rect 588542 52398 588778 52634
rect 588222 16718 588458 16954
rect 588542 16718 588778 16954
rect 588222 16398 588458 16634
rect 588542 16398 588778 16634
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 669218 589418 669454
rect 589502 669218 589738 669454
rect 589182 668898 589418 669134
rect 589502 668898 589738 669134
rect 589182 633218 589418 633454
rect 589502 633218 589738 633454
rect 589182 632898 589418 633134
rect 589502 632898 589738 633134
rect 589182 597218 589418 597454
rect 589502 597218 589738 597454
rect 589182 596898 589418 597134
rect 589502 596898 589738 597134
rect 589182 561218 589418 561454
rect 589502 561218 589738 561454
rect 589182 560898 589418 561134
rect 589502 560898 589738 561134
rect 589182 525218 589418 525454
rect 589502 525218 589738 525454
rect 589182 524898 589418 525134
rect 589502 524898 589738 525134
rect 589182 489218 589418 489454
rect 589502 489218 589738 489454
rect 589182 488898 589418 489134
rect 589502 488898 589738 489134
rect 589182 453218 589418 453454
rect 589502 453218 589738 453454
rect 589182 452898 589418 453134
rect 589502 452898 589738 453134
rect 589182 417218 589418 417454
rect 589502 417218 589738 417454
rect 589182 416898 589418 417134
rect 589502 416898 589738 417134
rect 589182 381218 589418 381454
rect 589502 381218 589738 381454
rect 589182 380898 589418 381134
rect 589502 380898 589738 381134
rect 589182 345218 589418 345454
rect 589502 345218 589738 345454
rect 589182 344898 589418 345134
rect 589502 344898 589738 345134
rect 589182 309218 589418 309454
rect 589502 309218 589738 309454
rect 589182 308898 589418 309134
rect 589502 308898 589738 309134
rect 589182 273218 589418 273454
rect 589502 273218 589738 273454
rect 589182 272898 589418 273134
rect 589502 272898 589738 273134
rect 589182 237218 589418 237454
rect 589502 237218 589738 237454
rect 589182 236898 589418 237134
rect 589502 236898 589738 237134
rect 589182 201218 589418 201454
rect 589502 201218 589738 201454
rect 589182 200898 589418 201134
rect 589502 200898 589738 201134
rect 589182 165218 589418 165454
rect 589502 165218 589738 165454
rect 589182 164898 589418 165134
rect 589502 164898 589738 165134
rect 589182 129218 589418 129454
rect 589502 129218 589738 129454
rect 589182 128898 589418 129134
rect 589502 128898 589738 129134
rect 589182 93218 589418 93454
rect 589502 93218 589738 93454
rect 589182 92898 589418 93134
rect 589502 92898 589738 93134
rect 589182 57218 589418 57454
rect 589502 57218 589738 57454
rect 589182 56898 589418 57134
rect 589502 56898 589738 57134
rect 589182 21218 589418 21454
rect 589502 21218 589738 21454
rect 589182 20898 589418 21134
rect 589502 20898 589738 21134
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 673718 590378 673954
rect 590462 673718 590698 673954
rect 590142 673398 590378 673634
rect 590462 673398 590698 673634
rect 590142 637718 590378 637954
rect 590462 637718 590698 637954
rect 590142 637398 590378 637634
rect 590462 637398 590698 637634
rect 590142 601718 590378 601954
rect 590462 601718 590698 601954
rect 590142 601398 590378 601634
rect 590462 601398 590698 601634
rect 590142 565718 590378 565954
rect 590462 565718 590698 565954
rect 590142 565398 590378 565634
rect 590462 565398 590698 565634
rect 590142 529718 590378 529954
rect 590462 529718 590698 529954
rect 590142 529398 590378 529634
rect 590462 529398 590698 529634
rect 590142 493718 590378 493954
rect 590462 493718 590698 493954
rect 590142 493398 590378 493634
rect 590462 493398 590698 493634
rect 590142 457718 590378 457954
rect 590462 457718 590698 457954
rect 590142 457398 590378 457634
rect 590462 457398 590698 457634
rect 590142 421718 590378 421954
rect 590462 421718 590698 421954
rect 590142 421398 590378 421634
rect 590462 421398 590698 421634
rect 590142 385718 590378 385954
rect 590462 385718 590698 385954
rect 590142 385398 590378 385634
rect 590462 385398 590698 385634
rect 590142 349718 590378 349954
rect 590462 349718 590698 349954
rect 590142 349398 590378 349634
rect 590462 349398 590698 349634
rect 590142 313718 590378 313954
rect 590462 313718 590698 313954
rect 590142 313398 590378 313634
rect 590462 313398 590698 313634
rect 590142 277718 590378 277954
rect 590462 277718 590698 277954
rect 590142 277398 590378 277634
rect 590462 277398 590698 277634
rect 590142 241718 590378 241954
rect 590462 241718 590698 241954
rect 590142 241398 590378 241634
rect 590462 241398 590698 241634
rect 590142 205718 590378 205954
rect 590462 205718 590698 205954
rect 590142 205398 590378 205634
rect 590462 205398 590698 205634
rect 590142 169718 590378 169954
rect 590462 169718 590698 169954
rect 590142 169398 590378 169634
rect 590462 169398 590698 169634
rect 590142 133718 590378 133954
rect 590462 133718 590698 133954
rect 590142 133398 590378 133634
rect 590462 133398 590698 133634
rect 590142 97718 590378 97954
rect 590462 97718 590698 97954
rect 590142 97398 590378 97634
rect 590462 97398 590698 97634
rect 590142 61718 590378 61954
rect 590462 61718 590698 61954
rect 590142 61398 590378 61634
rect 590462 61398 590698 61634
rect 590142 25718 590378 25954
rect 590462 25718 590698 25954
rect 590142 25398 590378 25634
rect 590462 25398 590698 25634
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 678218 591338 678454
rect 591422 678218 591658 678454
rect 591102 677898 591338 678134
rect 591422 677898 591658 678134
rect 591102 642218 591338 642454
rect 591422 642218 591658 642454
rect 591102 641898 591338 642134
rect 591422 641898 591658 642134
rect 591102 606218 591338 606454
rect 591422 606218 591658 606454
rect 591102 605898 591338 606134
rect 591422 605898 591658 606134
rect 591102 570218 591338 570454
rect 591422 570218 591658 570454
rect 591102 569898 591338 570134
rect 591422 569898 591658 570134
rect 591102 534218 591338 534454
rect 591422 534218 591658 534454
rect 591102 533898 591338 534134
rect 591422 533898 591658 534134
rect 591102 498218 591338 498454
rect 591422 498218 591658 498454
rect 591102 497898 591338 498134
rect 591422 497898 591658 498134
rect 591102 462218 591338 462454
rect 591422 462218 591658 462454
rect 591102 461898 591338 462134
rect 591422 461898 591658 462134
rect 591102 426218 591338 426454
rect 591422 426218 591658 426454
rect 591102 425898 591338 426134
rect 591422 425898 591658 426134
rect 591102 390218 591338 390454
rect 591422 390218 591658 390454
rect 591102 389898 591338 390134
rect 591422 389898 591658 390134
rect 591102 354218 591338 354454
rect 591422 354218 591658 354454
rect 591102 353898 591338 354134
rect 591422 353898 591658 354134
rect 591102 318218 591338 318454
rect 591422 318218 591658 318454
rect 591102 317898 591338 318134
rect 591422 317898 591658 318134
rect 591102 282218 591338 282454
rect 591422 282218 591658 282454
rect 591102 281898 591338 282134
rect 591422 281898 591658 282134
rect 591102 246218 591338 246454
rect 591422 246218 591658 246454
rect 591102 245898 591338 246134
rect 591422 245898 591658 246134
rect 591102 210218 591338 210454
rect 591422 210218 591658 210454
rect 591102 209898 591338 210134
rect 591422 209898 591658 210134
rect 591102 174218 591338 174454
rect 591422 174218 591658 174454
rect 591102 173898 591338 174134
rect 591422 173898 591658 174134
rect 591102 138218 591338 138454
rect 591422 138218 591658 138454
rect 591102 137898 591338 138134
rect 591422 137898 591658 138134
rect 591102 102218 591338 102454
rect 591422 102218 591658 102454
rect 591102 101898 591338 102134
rect 591422 101898 591658 102134
rect 591102 66218 591338 66454
rect 591422 66218 591658 66454
rect 591102 65898 591338 66134
rect 591422 65898 591658 66134
rect 591102 30218 591338 30454
rect 591422 30218 591658 30454
rect 591102 29898 591338 30134
rect 591422 29898 591658 30134
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 682718 592298 682954
rect 592382 682718 592618 682954
rect 592062 682398 592298 682634
rect 592382 682398 592618 682634
rect 592062 646718 592298 646954
rect 592382 646718 592618 646954
rect 592062 646398 592298 646634
rect 592382 646398 592618 646634
rect 592062 610718 592298 610954
rect 592382 610718 592618 610954
rect 592062 610398 592298 610634
rect 592382 610398 592618 610634
rect 592062 574718 592298 574954
rect 592382 574718 592618 574954
rect 592062 574398 592298 574634
rect 592382 574398 592618 574634
rect 592062 538718 592298 538954
rect 592382 538718 592618 538954
rect 592062 538398 592298 538634
rect 592382 538398 592618 538634
rect 592062 502718 592298 502954
rect 592382 502718 592618 502954
rect 592062 502398 592298 502634
rect 592382 502398 592618 502634
rect 592062 466718 592298 466954
rect 592382 466718 592618 466954
rect 592062 466398 592298 466634
rect 592382 466398 592618 466634
rect 592062 430718 592298 430954
rect 592382 430718 592618 430954
rect 592062 430398 592298 430634
rect 592382 430398 592618 430634
rect 592062 394718 592298 394954
rect 592382 394718 592618 394954
rect 592062 394398 592298 394634
rect 592382 394398 592618 394634
rect 592062 358718 592298 358954
rect 592382 358718 592618 358954
rect 592062 358398 592298 358634
rect 592382 358398 592618 358634
rect 592062 322718 592298 322954
rect 592382 322718 592618 322954
rect 592062 322398 592298 322634
rect 592382 322398 592618 322634
rect 592062 286718 592298 286954
rect 592382 286718 592618 286954
rect 592062 286398 592298 286634
rect 592382 286398 592618 286634
rect 592062 250718 592298 250954
rect 592382 250718 592618 250954
rect 592062 250398 592298 250634
rect 592382 250398 592618 250634
rect 592062 214718 592298 214954
rect 592382 214718 592618 214954
rect 592062 214398 592298 214634
rect 592382 214398 592618 214634
rect 592062 178718 592298 178954
rect 592382 178718 592618 178954
rect 592062 178398 592298 178634
rect 592382 178398 592618 178634
rect 592062 142718 592298 142954
rect 592382 142718 592618 142954
rect 592062 142398 592298 142634
rect 592382 142398 592618 142634
rect 592062 106718 592298 106954
rect 592382 106718 592618 106954
rect 592062 106398 592298 106634
rect 592382 106398 592618 106634
rect 592062 70718 592298 70954
rect 592382 70718 592618 70954
rect 592062 70398 592298 70634
rect 592382 70398 592618 70634
rect 592062 34718 592298 34954
rect 592382 34718 592618 34954
rect 592062 34398 592298 34634
rect 592382 34398 592618 34634
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 700954 592650 700986
rect -8726 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 592650 700954
rect -8726 700634 592650 700718
rect -8726 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 592650 700634
rect -8726 700366 592650 700398
rect -8726 696454 592650 696486
rect -8726 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 592650 696454
rect -8726 696134 592650 696218
rect -8726 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 592650 696134
rect -8726 695866 592650 695898
rect -8726 691954 592650 691986
rect -8726 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 592650 691954
rect -8726 691634 592650 691718
rect -8726 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 592650 691634
rect -8726 691366 592650 691398
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 682954 592650 682986
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect -8726 682634 592650 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect -8726 682366 592650 682398
rect -8726 678454 592650 678486
rect -8726 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 592650 678454
rect -8726 678134 592650 678218
rect -8726 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 592650 678134
rect -8726 677866 592650 677898
rect -8726 673954 592650 673986
rect -8726 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 592650 673954
rect -8726 673634 592650 673718
rect -8726 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 592650 673634
rect -8726 673366 592650 673398
rect -8726 669454 592650 669486
rect -8726 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 592650 669454
rect -8726 669134 592650 669218
rect -8726 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 592650 669134
rect -8726 668866 592650 668898
rect -8726 664954 592650 664986
rect -8726 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 592650 664954
rect -8726 664634 592650 664718
rect -8726 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 592650 664634
rect -8726 664366 592650 664398
rect -8726 660454 592650 660486
rect -8726 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 592650 660454
rect -8726 660134 592650 660218
rect -8726 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 592650 660134
rect -8726 659866 592650 659898
rect -8726 655954 592650 655986
rect -8726 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 592650 655954
rect -8726 655634 592650 655718
rect -8726 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 592650 655634
rect -8726 655366 592650 655398
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 646954 592650 646986
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect -8726 646634 592650 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect -8726 646366 592650 646398
rect -8726 642454 592650 642486
rect -8726 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 592650 642454
rect -8726 642134 592650 642218
rect -8726 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 592650 642134
rect -8726 641866 592650 641898
rect -8726 637954 592650 637986
rect -8726 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 592650 637954
rect -8726 637634 592650 637718
rect -8726 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 592650 637634
rect -8726 637366 592650 637398
rect -8726 633454 592650 633486
rect -8726 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 592650 633454
rect -8726 633134 592650 633218
rect -8726 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 592650 633134
rect -8726 632866 592650 632898
rect -8726 628954 592650 628986
rect -8726 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 592650 628954
rect -8726 628634 592650 628718
rect -8726 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 592650 628634
rect -8726 628366 592650 628398
rect -8726 624454 592650 624486
rect -8726 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 592650 624454
rect -8726 624134 592650 624218
rect -8726 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 592650 624134
rect -8726 623866 592650 623898
rect -8726 619954 592650 619986
rect -8726 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 592650 619954
rect -8726 619634 592650 619718
rect -8726 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 592650 619634
rect -8726 619366 592650 619398
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 610954 592650 610986
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect -8726 610634 592650 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect -8726 610366 592650 610398
rect -8726 606454 592650 606486
rect -8726 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 592650 606454
rect -8726 606134 592650 606218
rect -8726 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 592650 606134
rect -8726 605866 592650 605898
rect -8726 601954 592650 601986
rect -8726 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 592650 601954
rect -8726 601634 592650 601718
rect -8726 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 592650 601634
rect -8726 601366 592650 601398
rect -8726 597454 592650 597486
rect -8726 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 592650 597454
rect -8726 597134 592650 597218
rect -8726 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 592650 597134
rect -8726 596866 592650 596898
rect -8726 592954 592650 592986
rect -8726 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 592650 592954
rect -8726 592634 592650 592718
rect -8726 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 592650 592634
rect -8726 592366 592650 592398
rect -8726 588454 592650 588486
rect -8726 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 592650 588454
rect -8726 588134 592650 588218
rect -8726 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 592650 588134
rect -8726 587866 592650 587898
rect -8726 583954 592650 583986
rect -8726 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 592650 583954
rect -8726 583634 592650 583718
rect -8726 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 592650 583634
rect -8726 583366 592650 583398
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 574954 592650 574986
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect -8726 574634 592650 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect -8726 574366 592650 574398
rect -8726 570454 592650 570486
rect -8726 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 592650 570454
rect -8726 570134 592650 570218
rect -8726 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 592650 570134
rect -8726 569866 592650 569898
rect -8726 565954 592650 565986
rect -8726 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 592650 565954
rect -8726 565634 592650 565718
rect -8726 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 592650 565634
rect -8726 565366 592650 565398
rect -8726 561454 592650 561486
rect -8726 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 592650 561454
rect -8726 561134 592650 561218
rect -8726 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 592650 561134
rect -8726 560866 592650 560898
rect -8726 556954 592650 556986
rect -8726 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 592650 556954
rect -8726 556634 592650 556718
rect -8726 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 592650 556634
rect -8726 556366 592650 556398
rect -8726 552454 592650 552486
rect -8726 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 592650 552454
rect -8726 552134 592650 552218
rect -8726 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 592650 552134
rect -8726 551866 592650 551898
rect -8726 547954 592650 547986
rect -8726 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 592650 547954
rect -8726 547634 592650 547718
rect -8726 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 592650 547634
rect -8726 547366 592650 547398
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 538954 592650 538986
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect -8726 538634 592650 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect -8726 538366 592650 538398
rect -8726 534454 592650 534486
rect -8726 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 592650 534454
rect -8726 534134 592650 534218
rect -8726 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 592650 534134
rect -8726 533866 592650 533898
rect -8726 529954 592650 529986
rect -8726 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 592650 529954
rect -8726 529634 592650 529718
rect -8726 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 592650 529634
rect -8726 529366 592650 529398
rect -8726 525454 592650 525486
rect -8726 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 592650 525454
rect -8726 525134 592650 525218
rect -8726 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 592650 525134
rect -8726 524866 592650 524898
rect -8726 520954 592650 520986
rect -8726 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 592650 520954
rect -8726 520634 592650 520718
rect -8726 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 592650 520634
rect -8726 520366 592650 520398
rect -8726 516454 592650 516486
rect -8726 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 592650 516454
rect -8726 516134 592650 516218
rect -8726 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 592650 516134
rect -8726 515866 592650 515898
rect -8726 511954 592650 511986
rect -8726 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 592650 511954
rect -8726 511634 592650 511718
rect -8726 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 592650 511634
rect -8726 511366 592650 511398
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 502954 592650 502986
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect -8726 502634 592650 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect -8726 502366 592650 502398
rect -8726 498454 592650 498486
rect -8726 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 592650 498454
rect -8726 498134 592650 498218
rect -8726 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 592650 498134
rect -8726 497866 592650 497898
rect -8726 493954 592650 493986
rect -8726 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 592650 493954
rect -8726 493634 592650 493718
rect -8726 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 592650 493634
rect -8726 493366 592650 493398
rect -8726 489454 592650 489486
rect -8726 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 592650 489454
rect -8726 489134 592650 489218
rect -8726 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 592650 489134
rect -8726 488866 592650 488898
rect -8726 484954 592650 484986
rect -8726 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 592650 484954
rect -8726 484634 592650 484718
rect -8726 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 592650 484634
rect -8726 484366 592650 484398
rect -8726 480454 592650 480486
rect -8726 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 592650 480454
rect -8726 480134 592650 480218
rect -8726 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 592650 480134
rect -8726 479866 592650 479898
rect -8726 475954 592650 475986
rect -8726 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 592650 475954
rect -8726 475634 592650 475718
rect -8726 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 592650 475634
rect -8726 475366 592650 475398
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 466954 592650 466986
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect -8726 466634 592650 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect -8726 466366 592650 466398
rect -8726 462454 592650 462486
rect -8726 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 592650 462454
rect -8726 462134 592650 462218
rect -8726 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 592650 462134
rect -8726 461866 592650 461898
rect -8726 457954 592650 457986
rect -8726 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 592650 457954
rect -8726 457634 592650 457718
rect -8726 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 592650 457634
rect -8726 457366 592650 457398
rect -8726 453454 592650 453486
rect -8726 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 592650 453454
rect -8726 453134 592650 453218
rect -8726 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 592650 453134
rect -8726 452866 592650 452898
rect -8726 448954 592650 448986
rect -8726 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 592650 448954
rect -8726 448634 592650 448718
rect -8726 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 592650 448634
rect -8726 448366 592650 448398
rect -8726 444454 592650 444486
rect -8726 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 592650 444454
rect -8726 444134 592650 444218
rect -8726 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 592650 444134
rect -8726 443866 592650 443898
rect -8726 439954 592650 439986
rect -8726 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 592650 439954
rect -8726 439634 592650 439718
rect -8726 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 592650 439634
rect -8726 439366 592650 439398
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 430954 592650 430986
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect -8726 430634 592650 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect -8726 430366 592650 430398
rect -8726 426454 592650 426486
rect -8726 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 592650 426454
rect -8726 426134 592650 426218
rect -8726 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 592650 426134
rect -8726 425866 592650 425898
rect -8726 421954 592650 421986
rect -8726 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 592650 421954
rect -8726 421634 592650 421718
rect -8726 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 592650 421634
rect -8726 421366 592650 421398
rect -8726 417454 592650 417486
rect -8726 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 592650 417454
rect -8726 417134 592650 417218
rect -8726 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 592650 417134
rect -8726 416866 592650 416898
rect -8726 412954 592650 412986
rect -8726 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 592650 412954
rect -8726 412634 592650 412718
rect -8726 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 592650 412634
rect -8726 412366 592650 412398
rect -8726 408454 592650 408486
rect -8726 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 592650 408454
rect -8726 408134 592650 408218
rect -8726 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 592650 408134
rect -8726 407866 592650 407898
rect -8726 403954 592650 403986
rect -8726 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 592650 403954
rect -8726 403634 592650 403718
rect -8726 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 592650 403634
rect -8726 403366 592650 403398
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 394954 592650 394986
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect -8726 394634 592650 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect -8726 394366 592650 394398
rect -8726 390454 592650 390486
rect -8726 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 592650 390454
rect -8726 390134 592650 390218
rect -8726 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 592650 390134
rect -8726 389866 592650 389898
rect -8726 385954 592650 385986
rect -8726 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 592650 385954
rect -8726 385634 592650 385718
rect -8726 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 592650 385634
rect -8726 385366 592650 385398
rect -8726 381454 592650 381486
rect -8726 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 592650 381454
rect -8726 381134 592650 381218
rect -8726 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 592650 381134
rect -8726 380866 592650 380898
rect -8726 376954 592650 376986
rect -8726 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 592650 376954
rect -8726 376634 592650 376718
rect -8726 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 592650 376634
rect -8726 376366 592650 376398
rect -8726 372454 592650 372486
rect -8726 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 592650 372454
rect -8726 372134 592650 372218
rect -8726 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 592650 372134
rect -8726 371866 592650 371898
rect -8726 367954 592650 367986
rect -8726 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 592650 367954
rect -8726 367634 592650 367718
rect -8726 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 592650 367634
rect -8726 367366 592650 367398
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 358954 592650 358986
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect -8726 358634 592650 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect -8726 358366 592650 358398
rect -8726 354454 592650 354486
rect -8726 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 244826 354454
rect 245062 354218 245146 354454
rect 245382 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 592650 354454
rect -8726 354134 592650 354218
rect -8726 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 244826 354134
rect 245062 353898 245146 354134
rect 245382 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 592650 354134
rect -8726 353866 592650 353898
rect -8726 349954 592650 349986
rect -8726 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 240326 349954
rect 240562 349718 240646 349954
rect 240882 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 592650 349954
rect -8726 349634 592650 349718
rect -8726 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 240326 349634
rect 240562 349398 240646 349634
rect 240882 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 592650 349634
rect -8726 349366 592650 349398
rect -8726 345454 592650 345486
rect -8726 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 592650 345454
rect -8726 345134 592650 345218
rect -8726 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 592650 345134
rect -8726 344866 592650 344898
rect -8726 340954 592650 340986
rect -8726 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 592650 340954
rect -8726 340634 592650 340718
rect -8726 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 592650 340634
rect -8726 340366 592650 340398
rect -8726 336454 592650 336486
rect -8726 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 592650 336454
rect -8726 336134 592650 336218
rect -8726 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 592650 336134
rect -8726 335866 592650 335898
rect -8726 331954 592650 331986
rect -8726 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 592650 331954
rect -8726 331634 592650 331718
rect -8726 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 592650 331634
rect -8726 331366 592650 331398
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 322954 592650 322986
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect -8726 322634 592650 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect -8726 322366 592650 322398
rect -8726 318454 592650 318486
rect -8726 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 592650 318454
rect -8726 318134 592650 318218
rect -8726 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 592650 318134
rect -8726 317866 592650 317898
rect -8726 313954 592650 313986
rect -8726 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 592650 313954
rect -8726 313634 592650 313718
rect -8726 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 592650 313634
rect -8726 313366 592650 313398
rect -8726 309454 592650 309486
rect -8726 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 592650 309454
rect -8726 309134 592650 309218
rect -8726 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 592650 309134
rect -8726 308866 592650 308898
rect -8726 304954 592650 304986
rect -8726 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 592650 304954
rect -8726 304634 592650 304718
rect -8726 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 592650 304634
rect -8726 304366 592650 304398
rect -8726 300454 592650 300486
rect -8726 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 592650 300454
rect -8726 300134 592650 300218
rect -8726 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 592650 300134
rect -8726 299866 592650 299898
rect -8726 295954 592650 295986
rect -8726 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 592650 295954
rect -8726 295634 592650 295718
rect -8726 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 592650 295634
rect -8726 295366 592650 295398
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 286954 592650 286986
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect -8726 286634 592650 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect -8726 286366 592650 286398
rect -8726 282454 592650 282486
rect -8726 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 592650 282454
rect -8726 282134 592650 282218
rect -8726 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 592650 282134
rect -8726 281866 592650 281898
rect -8726 277954 592650 277986
rect -8726 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 592650 277954
rect -8726 277634 592650 277718
rect -8726 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 592650 277634
rect -8726 277366 592650 277398
rect -8726 273454 592650 273486
rect -8726 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 592650 273454
rect -8726 273134 592650 273218
rect -8726 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 592650 273134
rect -8726 272866 592650 272898
rect -8726 268954 592650 268986
rect -8726 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 592650 268954
rect -8726 268634 592650 268718
rect -8726 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 592650 268634
rect -8726 268366 592650 268398
rect -8726 264454 592650 264486
rect -8726 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 592650 264454
rect -8726 264134 592650 264218
rect -8726 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 592650 264134
rect -8726 263866 592650 263898
rect -8726 259954 592650 259986
rect -8726 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 592650 259954
rect -8726 259634 592650 259718
rect -8726 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 592650 259634
rect -8726 259366 592650 259398
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 250954 592650 250986
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect -8726 250634 592650 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect -8726 250366 592650 250398
rect -8726 246454 592650 246486
rect -8726 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 136826 246454
rect 137062 246218 137146 246454
rect 137382 246218 172826 246454
rect 173062 246218 173146 246454
rect 173382 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 592650 246454
rect -8726 246134 592650 246218
rect -8726 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 136826 246134
rect 137062 245898 137146 246134
rect 137382 245898 172826 246134
rect 173062 245898 173146 246134
rect 173382 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 592650 246134
rect -8726 245866 592650 245898
rect -8726 241954 592650 241986
rect -8726 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241953 420326 241954
rect 24882 241718 71462 241953
rect -8726 241717 71462 241718
rect 71698 241717 71782 241953
rect 72018 241717 72102 241953
rect 72338 241717 72422 241953
rect 72658 241717 72742 241953
rect 72978 241717 73062 241953
rect 73298 241717 73382 241953
rect 73618 241717 73702 241953
rect 73938 241717 74022 241953
rect 74258 241717 74342 241953
rect 74578 241717 74662 241953
rect 74898 241717 74982 241953
rect 75218 241717 75302 241953
rect 75538 241717 75622 241953
rect 75858 241717 75942 241953
rect 76178 241717 76262 241953
rect 76498 241717 76582 241953
rect 76818 241717 76902 241953
rect 77138 241718 420326 241953
rect 420562 241718 420646 241954
rect 420882 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 592650 241954
rect 77138 241717 592650 241718
rect -8726 241634 592650 241717
rect -8726 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241633 420326 241634
rect 24882 241398 71462 241633
rect -8726 241397 71462 241398
rect 71698 241397 71782 241633
rect 72018 241397 72102 241633
rect 72338 241397 72422 241633
rect 72658 241397 72742 241633
rect 72978 241397 73062 241633
rect 73298 241397 73382 241633
rect 73618 241397 73702 241633
rect 73938 241397 74022 241633
rect 74258 241397 74342 241633
rect 74578 241397 74662 241633
rect 74898 241397 74982 241633
rect 75218 241397 75302 241633
rect 75538 241397 75622 241633
rect 75858 241397 75942 241633
rect 76178 241397 76262 241633
rect 76498 241397 76582 241633
rect 76818 241397 76902 241633
rect 77138 241398 420326 241633
rect 420562 241398 420646 241634
rect 420882 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 592650 241634
rect 77138 241397 592650 241398
rect -8726 241366 592650 241397
rect -8726 237454 592650 237486
rect -8726 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237453 415826 237454
rect 20382 237218 46039 237453
rect -8726 237217 46039 237218
rect 46275 237217 46359 237453
rect 46595 237217 46679 237453
rect 46915 237217 46999 237453
rect 47235 237217 47319 237453
rect 47555 237217 47639 237453
rect 47875 237217 47959 237453
rect 48195 237217 48279 237453
rect 48515 237217 48599 237453
rect 48835 237217 48919 237453
rect 49155 237217 49239 237453
rect 49475 237217 49559 237453
rect 49795 237217 49879 237453
rect 50115 237217 50199 237453
rect 50435 237217 50519 237453
rect 50755 237218 415826 237453
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 592650 237454
rect 50755 237217 592650 237218
rect -8726 237134 592650 237217
rect -8726 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 237133 415826 237134
rect 20382 236898 46039 237133
rect -8726 236897 46039 236898
rect 46275 236897 46359 237133
rect 46595 236897 46679 237133
rect 46915 236897 46999 237133
rect 47235 236897 47319 237133
rect 47555 236897 47639 237133
rect 47875 236897 47959 237133
rect 48195 236897 48279 237133
rect 48515 236897 48599 237133
rect 48835 236897 48919 237133
rect 49155 236897 49239 237133
rect 49475 236897 49559 237133
rect 49795 236897 49879 237133
rect 50115 236897 50199 237133
rect 50435 236897 50519 237133
rect 50755 236898 415826 237133
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 592650 237134
rect 50755 236897 592650 236898
rect -8726 236866 592650 236897
rect -8726 232954 592650 232986
rect -8726 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 592650 232954
rect -8726 232634 592650 232718
rect -8726 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 592650 232634
rect -8726 232366 592650 232398
rect -8726 228454 592650 228486
rect -8726 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228453 406826 228454
rect 11382 228218 46826 228453
rect -8726 228217 46826 228218
rect 47062 228217 47146 228453
rect 47382 228217 82826 228453
rect 83062 228217 83146 228453
rect 83382 228217 118826 228453
rect 119062 228217 119146 228453
rect 119382 228217 190826 228453
rect 191062 228217 191146 228453
rect 191382 228217 226826 228453
rect 227062 228217 227146 228453
rect 227382 228217 262826 228453
rect 263062 228217 263146 228453
rect 263382 228217 298826 228453
rect 299062 228217 299146 228453
rect 299382 228217 334826 228453
rect 335062 228217 335146 228453
rect 335382 228217 370826 228453
rect 371062 228217 371146 228453
rect 371382 228218 406826 228453
rect 407062 228218 407146 228454
rect 407382 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 592650 228454
rect 371382 228217 592650 228218
rect -8726 228134 592650 228217
rect -8726 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 228133 406826 228134
rect 11382 227898 46826 228133
rect -8726 227897 46826 227898
rect 47062 227897 47146 228133
rect 47382 227897 82826 228133
rect 83062 227897 83146 228133
rect 83382 227897 118826 228133
rect 119062 227897 119146 228133
rect 119382 227897 190826 228133
rect 191062 227897 191146 228133
rect 191382 227897 226826 228133
rect 227062 227897 227146 228133
rect 227382 227897 262826 228133
rect 263062 227897 263146 228133
rect 263382 227897 298826 228133
rect 299062 227897 299146 228133
rect 299382 227897 334826 228133
rect 335062 227897 335146 228133
rect 335382 227897 370826 228133
rect 371062 227897 371146 228133
rect 371382 227898 406826 228133
rect 407062 227898 407146 228134
rect 407382 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 592650 228134
rect 371382 227897 592650 227898
rect -8726 227866 592650 227897
rect -8726 223954 592650 223986
rect -8726 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 592650 223954
rect -8726 223634 592650 223718
rect -8726 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 592650 223634
rect -8726 223366 592650 223398
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 214954 592650 214986
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect -8726 214634 592650 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect -8726 214366 592650 214398
rect -8726 210454 592650 210486
rect -8726 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 592650 210454
rect -8726 210134 592650 210218
rect -8726 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 592650 210134
rect -8726 209866 592650 209898
rect -8726 205954 592650 205986
rect -8726 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205718 136036 205954
rect 136272 205718 136356 205954
rect 136592 205718 136676 205954
rect 136912 205718 136996 205954
rect 137232 205718 137316 205954
rect 137552 205718 137636 205954
rect 137872 205718 137956 205954
rect 138192 205718 138276 205954
rect 138512 205718 138596 205954
rect 138832 205718 138916 205954
rect 139152 205718 139236 205954
rect 139472 205718 139556 205954
rect 139792 205718 139876 205954
rect 140112 205718 140196 205954
rect 140432 205718 140516 205954
rect 140752 205718 140836 205954
rect 141072 205718 141156 205954
rect 141392 205718 141476 205954
rect 141712 205718 141796 205954
rect 142032 205718 142116 205954
rect 142352 205718 142436 205954
rect 142672 205718 142756 205954
rect 142992 205718 143076 205954
rect 143312 205718 143396 205954
rect 143632 205718 143716 205954
rect 143952 205718 144036 205954
rect 144272 205718 144356 205954
rect 144592 205718 144676 205954
rect 144912 205718 144996 205954
rect 145232 205718 145316 205954
rect 145552 205718 145636 205954
rect 145872 205718 145956 205954
rect 146192 205718 146276 205954
rect 146512 205718 146596 205954
rect 146832 205718 146916 205954
rect 147152 205718 147236 205954
rect 147472 205718 147556 205954
rect 147792 205718 147876 205954
rect 148112 205718 148196 205954
rect 148432 205718 148516 205954
rect 148752 205718 148836 205954
rect 149072 205718 149156 205954
rect 149392 205718 149476 205954
rect 149712 205718 149796 205954
rect 150032 205718 150116 205954
rect 150352 205718 150436 205954
rect 150672 205718 150756 205954
rect 150992 205718 151076 205954
rect 151312 205718 151396 205954
rect 151632 205718 151716 205954
rect 151952 205718 152036 205954
rect 152272 205718 152356 205954
rect 152592 205718 152676 205954
rect 152912 205718 152996 205954
rect 153232 205718 153316 205954
rect 153552 205718 153636 205954
rect 153872 205718 153956 205954
rect 154192 205718 154276 205954
rect 154512 205718 154596 205954
rect 154832 205718 154916 205954
rect 155152 205718 155236 205954
rect 155472 205718 155556 205954
rect 155792 205718 155876 205954
rect 156112 205718 156196 205954
rect 156432 205718 156516 205954
rect 156752 205718 156836 205954
rect 157072 205718 157156 205954
rect 157392 205718 157476 205954
rect 157712 205718 157796 205954
rect 158032 205718 158116 205954
rect 158352 205718 158436 205954
rect 158672 205718 158756 205954
rect 158992 205718 159076 205954
rect 159312 205718 159396 205954
rect 159632 205718 159716 205954
rect 159952 205718 160036 205954
rect 160272 205718 160356 205954
rect 160592 205718 160676 205954
rect 160912 205718 160996 205954
rect 161232 205718 161316 205954
rect 161552 205718 161636 205954
rect 161872 205718 161956 205954
rect 162192 205718 162276 205954
rect 162512 205718 162596 205954
rect 162832 205718 162916 205954
rect 163152 205718 163236 205954
rect 163472 205718 163556 205954
rect 163792 205718 163876 205954
rect 164112 205718 164196 205954
rect 164432 205718 164516 205954
rect 164752 205718 164836 205954
rect 165072 205718 165156 205954
rect 165392 205718 168326 205954
rect 168562 205718 168646 205954
rect 168882 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 592650 205954
rect -8726 205634 592650 205718
rect -8726 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205398 136036 205634
rect 136272 205398 136356 205634
rect 136592 205398 136676 205634
rect 136912 205398 136996 205634
rect 137232 205398 137316 205634
rect 137552 205398 137636 205634
rect 137872 205398 137956 205634
rect 138192 205398 138276 205634
rect 138512 205398 138596 205634
rect 138832 205398 138916 205634
rect 139152 205398 139236 205634
rect 139472 205398 139556 205634
rect 139792 205398 139876 205634
rect 140112 205398 140196 205634
rect 140432 205398 140516 205634
rect 140752 205398 140836 205634
rect 141072 205398 141156 205634
rect 141392 205398 141476 205634
rect 141712 205398 141796 205634
rect 142032 205398 142116 205634
rect 142352 205398 142436 205634
rect 142672 205398 142756 205634
rect 142992 205398 143076 205634
rect 143312 205398 143396 205634
rect 143632 205398 143716 205634
rect 143952 205398 144036 205634
rect 144272 205398 144356 205634
rect 144592 205398 144676 205634
rect 144912 205398 144996 205634
rect 145232 205398 145316 205634
rect 145552 205398 145636 205634
rect 145872 205398 145956 205634
rect 146192 205398 146276 205634
rect 146512 205398 146596 205634
rect 146832 205398 146916 205634
rect 147152 205398 147236 205634
rect 147472 205398 147556 205634
rect 147792 205398 147876 205634
rect 148112 205398 148196 205634
rect 148432 205398 148516 205634
rect 148752 205398 148836 205634
rect 149072 205398 149156 205634
rect 149392 205398 149476 205634
rect 149712 205398 149796 205634
rect 150032 205398 150116 205634
rect 150352 205398 150436 205634
rect 150672 205398 150756 205634
rect 150992 205398 151076 205634
rect 151312 205398 151396 205634
rect 151632 205398 151716 205634
rect 151952 205398 152036 205634
rect 152272 205398 152356 205634
rect 152592 205398 152676 205634
rect 152912 205398 152996 205634
rect 153232 205398 153316 205634
rect 153552 205398 153636 205634
rect 153872 205398 153956 205634
rect 154192 205398 154276 205634
rect 154512 205398 154596 205634
rect 154832 205398 154916 205634
rect 155152 205398 155236 205634
rect 155472 205398 155556 205634
rect 155792 205398 155876 205634
rect 156112 205398 156196 205634
rect 156432 205398 156516 205634
rect 156752 205398 156836 205634
rect 157072 205398 157156 205634
rect 157392 205398 157476 205634
rect 157712 205398 157796 205634
rect 158032 205398 158116 205634
rect 158352 205398 158436 205634
rect 158672 205398 158756 205634
rect 158992 205398 159076 205634
rect 159312 205398 159396 205634
rect 159632 205398 159716 205634
rect 159952 205398 160036 205634
rect 160272 205398 160356 205634
rect 160592 205398 160676 205634
rect 160912 205398 160996 205634
rect 161232 205398 161316 205634
rect 161552 205398 161636 205634
rect 161872 205398 161956 205634
rect 162192 205398 162276 205634
rect 162512 205398 162596 205634
rect 162832 205398 162916 205634
rect 163152 205398 163236 205634
rect 163472 205398 163556 205634
rect 163792 205398 163876 205634
rect 164112 205398 164196 205634
rect 164432 205398 164516 205634
rect 164752 205398 164836 205634
rect 165072 205398 165156 205634
rect 165392 205398 168326 205634
rect 168562 205398 168646 205634
rect 168882 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 592650 205634
rect -8726 205366 592650 205398
rect -8726 201454 592650 201486
rect -8726 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 137376 201454
rect 137612 201218 137696 201454
rect 137932 201218 138016 201454
rect 138252 201218 138336 201454
rect 138572 201218 138656 201454
rect 138892 201218 138976 201454
rect 139212 201218 139296 201454
rect 139532 201218 139616 201454
rect 139852 201218 139936 201454
rect 140172 201218 140256 201454
rect 140492 201218 140576 201454
rect 140812 201218 140896 201454
rect 141132 201218 141216 201454
rect 141452 201218 141536 201454
rect 141772 201218 141856 201454
rect 142092 201218 142176 201454
rect 142412 201218 142496 201454
rect 142732 201218 142816 201454
rect 143052 201218 143136 201454
rect 143372 201218 143456 201454
rect 143692 201218 143776 201454
rect 144012 201218 144096 201454
rect 144332 201218 144416 201454
rect 144652 201218 144736 201454
rect 144972 201218 145056 201454
rect 145292 201218 145376 201454
rect 145612 201218 145696 201454
rect 145932 201218 146016 201454
rect 146252 201218 146336 201454
rect 146572 201218 146656 201454
rect 146892 201218 146976 201454
rect 147212 201218 147296 201454
rect 147532 201218 147616 201454
rect 147852 201218 147936 201454
rect 148172 201218 148256 201454
rect 148492 201218 148576 201454
rect 148812 201218 148896 201454
rect 149132 201218 149216 201454
rect 149452 201218 149536 201454
rect 149772 201218 149856 201454
rect 150092 201218 150176 201454
rect 150412 201218 150496 201454
rect 150732 201218 150816 201454
rect 151052 201218 151136 201454
rect 151372 201218 151456 201454
rect 151692 201218 151776 201454
rect 152012 201218 152096 201454
rect 152332 201218 152416 201454
rect 152652 201218 152736 201454
rect 152972 201218 153056 201454
rect 153292 201218 153376 201454
rect 153612 201218 153696 201454
rect 153932 201218 154016 201454
rect 154252 201218 154336 201454
rect 154572 201218 154656 201454
rect 154892 201218 154976 201454
rect 155212 201218 155296 201454
rect 155532 201218 155616 201454
rect 155852 201218 155936 201454
rect 156172 201218 156256 201454
rect 156492 201218 156576 201454
rect 156812 201218 156896 201454
rect 157132 201218 157216 201454
rect 157452 201218 157536 201454
rect 157772 201218 157856 201454
rect 158092 201218 158176 201454
rect 158412 201218 158496 201454
rect 158732 201218 158816 201454
rect 159052 201218 159136 201454
rect 159372 201218 159456 201454
rect 159692 201218 159776 201454
rect 160012 201218 160096 201454
rect 160332 201218 160416 201454
rect 160652 201218 160736 201454
rect 160972 201218 161056 201454
rect 161292 201218 161376 201454
rect 161612 201218 161696 201454
rect 161932 201218 162016 201454
rect 162252 201218 162336 201454
rect 162572 201218 162656 201454
rect 162892 201218 162976 201454
rect 163212 201218 163296 201454
rect 163532 201218 163616 201454
rect 163852 201218 163936 201454
rect 164172 201218 164256 201454
rect 164492 201218 164576 201454
rect 164812 201218 164896 201454
rect 165132 201218 165216 201454
rect 165452 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 592650 201454
rect -8726 201134 592650 201218
rect -8726 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 137376 201134
rect 137612 200898 137696 201134
rect 137932 200898 138016 201134
rect 138252 200898 138336 201134
rect 138572 200898 138656 201134
rect 138892 200898 138976 201134
rect 139212 200898 139296 201134
rect 139532 200898 139616 201134
rect 139852 200898 139936 201134
rect 140172 200898 140256 201134
rect 140492 200898 140576 201134
rect 140812 200898 140896 201134
rect 141132 200898 141216 201134
rect 141452 200898 141536 201134
rect 141772 200898 141856 201134
rect 142092 200898 142176 201134
rect 142412 200898 142496 201134
rect 142732 200898 142816 201134
rect 143052 200898 143136 201134
rect 143372 200898 143456 201134
rect 143692 200898 143776 201134
rect 144012 200898 144096 201134
rect 144332 200898 144416 201134
rect 144652 200898 144736 201134
rect 144972 200898 145056 201134
rect 145292 200898 145376 201134
rect 145612 200898 145696 201134
rect 145932 200898 146016 201134
rect 146252 200898 146336 201134
rect 146572 200898 146656 201134
rect 146892 200898 146976 201134
rect 147212 200898 147296 201134
rect 147532 200898 147616 201134
rect 147852 200898 147936 201134
rect 148172 200898 148256 201134
rect 148492 200898 148576 201134
rect 148812 200898 148896 201134
rect 149132 200898 149216 201134
rect 149452 200898 149536 201134
rect 149772 200898 149856 201134
rect 150092 200898 150176 201134
rect 150412 200898 150496 201134
rect 150732 200898 150816 201134
rect 151052 200898 151136 201134
rect 151372 200898 151456 201134
rect 151692 200898 151776 201134
rect 152012 200898 152096 201134
rect 152332 200898 152416 201134
rect 152652 200898 152736 201134
rect 152972 200898 153056 201134
rect 153292 200898 153376 201134
rect 153612 200898 153696 201134
rect 153932 200898 154016 201134
rect 154252 200898 154336 201134
rect 154572 200898 154656 201134
rect 154892 200898 154976 201134
rect 155212 200898 155296 201134
rect 155532 200898 155616 201134
rect 155852 200898 155936 201134
rect 156172 200898 156256 201134
rect 156492 200898 156576 201134
rect 156812 200898 156896 201134
rect 157132 200898 157216 201134
rect 157452 200898 157536 201134
rect 157772 200898 157856 201134
rect 158092 200898 158176 201134
rect 158412 200898 158496 201134
rect 158732 200898 158816 201134
rect 159052 200898 159136 201134
rect 159372 200898 159456 201134
rect 159692 200898 159776 201134
rect 160012 200898 160096 201134
rect 160332 200898 160416 201134
rect 160652 200898 160736 201134
rect 160972 200898 161056 201134
rect 161292 200898 161376 201134
rect 161612 200898 161696 201134
rect 161932 200898 162016 201134
rect 162252 200898 162336 201134
rect 162572 200898 162656 201134
rect 162892 200898 162976 201134
rect 163212 200898 163296 201134
rect 163532 200898 163616 201134
rect 163852 200898 163936 201134
rect 164172 200898 164256 201134
rect 164492 200898 164576 201134
rect 164812 200898 164896 201134
rect 165132 200898 165216 201134
rect 165452 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 592650 201134
rect -8726 200866 592650 200898
rect -8726 196954 592650 196986
rect -8726 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 592650 196954
rect -8726 196634 592650 196718
rect -8726 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 592650 196634
rect -8726 196366 592650 196398
rect -8726 192454 592650 192486
rect -8726 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 592650 192454
rect -8726 192134 592650 192218
rect -8726 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 592650 192134
rect -8726 191866 592650 191898
rect -8726 187954 592650 187986
rect -8726 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 592650 187954
rect -8726 187634 592650 187718
rect -8726 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 592650 187634
rect -8726 187366 592650 187398
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 178954 592650 178986
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect -8726 178634 592650 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect -8726 178366 592650 178398
rect -8726 174454 592650 174486
rect -8726 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 316826 174454
rect 317062 174218 317146 174454
rect 317382 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 592650 174454
rect -8726 174134 592650 174218
rect -8726 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 316826 174134
rect 317062 173898 317146 174134
rect 317382 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 592650 174134
rect -8726 173866 592650 173898
rect -8726 169954 592650 169986
rect -8726 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 132326 169954
rect 132562 169718 132646 169954
rect 132882 169718 168326 169954
rect 168562 169718 168646 169954
rect 168882 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 312326 169954
rect 312562 169718 312646 169954
rect 312882 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 592650 169954
rect -8726 169634 592650 169718
rect -8726 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 132326 169634
rect 132562 169398 132646 169634
rect 132882 169398 168326 169634
rect 168562 169398 168646 169634
rect 168882 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 312326 169634
rect 312562 169398 312646 169634
rect 312882 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 592650 169634
rect -8726 169366 592650 169398
rect -8726 165454 592650 165486
rect -8726 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 592650 165454
rect -8726 165134 592650 165218
rect -8726 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 592650 165134
rect -8726 164866 592650 164898
rect -8726 160954 592650 160986
rect -8726 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 592650 160954
rect -8726 160634 592650 160718
rect -8726 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 592650 160634
rect -8726 160366 592650 160398
rect -8726 156454 592650 156486
rect -8726 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 592650 156454
rect -8726 156134 592650 156218
rect -8726 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 592650 156134
rect -8726 155866 592650 155898
rect -8726 151954 592650 151986
rect -8726 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 592650 151954
rect -8726 151634 592650 151718
rect -8726 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 592650 151634
rect -8726 151366 592650 151398
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 142954 592650 142986
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect -8726 142634 592650 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect -8726 142366 592650 142398
rect -8726 138454 592650 138486
rect -8726 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 592650 138454
rect -8726 138134 592650 138218
rect -8726 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 592650 138134
rect -8726 137866 592650 137898
rect -8726 133954 592650 133986
rect -8726 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 592650 133954
rect -8726 133634 592650 133718
rect -8726 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 592650 133634
rect -8726 133366 592650 133398
rect -8726 129454 592650 129486
rect -8726 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 592650 129454
rect -8726 129134 592650 129218
rect -8726 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 592650 129134
rect -8726 128866 592650 128898
rect -8726 124954 592650 124986
rect -8726 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 592650 124954
rect -8726 124634 592650 124718
rect -8726 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 592650 124634
rect -8726 124366 592650 124398
rect -8726 120454 592650 120486
rect -8726 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 592650 120454
rect -8726 120134 592650 120218
rect -8726 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 592650 120134
rect -8726 119866 592650 119898
rect -8726 115954 592650 115986
rect -8726 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 139610 115954
rect 139846 115718 170330 115954
rect 170566 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 592650 115954
rect -8726 115634 592650 115718
rect -8726 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 139610 115634
rect 139846 115398 170330 115634
rect 170566 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 592650 115634
rect -8726 115366 592650 115398
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 124250 111454
rect 124486 111218 154970 111454
rect 155206 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 124250 111134
rect 124486 110898 154970 111134
rect 155206 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 106954 592650 106986
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect -8726 106634 592650 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect -8726 106366 592650 106398
rect -8726 102454 592650 102486
rect -8726 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 592650 102454
rect -8726 102134 592650 102218
rect -8726 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 592650 102134
rect -8726 101866 592650 101898
rect -8726 97954 592650 97986
rect -8726 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 592650 97954
rect -8726 97634 592650 97718
rect -8726 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 592650 97634
rect -8726 97366 592650 97398
rect -8726 93454 592650 93486
rect -8726 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 592650 93454
rect -8726 93134 592650 93218
rect -8726 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 592650 93134
rect -8726 92866 592650 92898
rect -8726 88954 592650 88986
rect -8726 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 592650 88954
rect -8726 88634 592650 88718
rect -8726 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 592650 88634
rect -8726 88366 592650 88398
rect -8726 84454 592650 84486
rect -8726 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 592650 84454
rect -8726 84134 592650 84218
rect -8726 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 592650 84134
rect -8726 83866 592650 83898
rect -8726 79954 592650 79986
rect -8726 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 592650 79954
rect -8726 79634 592650 79718
rect -8726 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 592650 79634
rect -8726 79366 592650 79398
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 70954 592650 70986
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect -8726 70634 592650 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect -8726 70366 592650 70398
rect -8726 66454 592650 66486
rect -8726 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 592650 66454
rect -8726 66134 592650 66218
rect -8726 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 592650 66134
rect -8726 65866 592650 65898
rect -8726 61954 592650 61986
rect -8726 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 592650 61954
rect -8726 61634 592650 61718
rect -8726 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 592650 61634
rect -8726 61366 592650 61398
rect -8726 57454 592650 57486
rect -8726 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 592650 57454
rect -8726 57134 592650 57218
rect -8726 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 592650 57134
rect -8726 56866 592650 56898
rect -8726 52954 592650 52986
rect -8726 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 592650 52954
rect -8726 52634 592650 52718
rect -8726 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 592650 52634
rect -8726 52366 592650 52398
rect -8726 48454 592650 48486
rect -8726 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 592650 48454
rect -8726 48134 592650 48218
rect -8726 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 592650 48134
rect -8726 47866 592650 47898
rect -8726 43954 592650 43986
rect -8726 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 592650 43954
rect -8726 43634 592650 43718
rect -8726 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 592650 43634
rect -8726 43366 592650 43398
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 34954 592650 34986
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect -8726 34634 592650 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect -8726 34366 592650 34398
rect -8726 30454 592650 30486
rect -8726 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 592650 30454
rect -8726 30134 592650 30218
rect -8726 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 592650 30134
rect -8726 29866 592650 29898
rect -8726 25954 592650 25986
rect -8726 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 592650 25954
rect -8726 25634 592650 25718
rect -8726 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 592650 25634
rect -8726 25366 592650 25398
rect -8726 21454 592650 21486
rect -8726 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 592650 21454
rect -8726 21134 592650 21218
rect -8726 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 592650 21134
rect -8726 20866 592650 20898
rect -8726 16954 592650 16986
rect -8726 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 592650 16954
rect -8726 16634 592650 16718
rect -8726 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 592650 16634
rect -8726 16366 592650 16398
rect -8726 12454 592650 12486
rect -8726 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 592650 12454
rect -8726 12134 592650 12218
rect -8726 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 592650 12134
rect -8726 11866 592650 11898
rect -8726 7954 592650 7986
rect -8726 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 592650 7954
rect -8726 7634 592650 7718
rect -8726 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 592650 7634
rect -8726 7366 592650 7398
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use PD1  PD1_macro0
timestamp 0
transform 1 0 22000 0 1 232484
box 24000 -2000 380300 9600
use rlbp_macro  rlbp_macro0
timestamp 0
transform 1 0 120000 0 1 80000
box 0 0 60000 60000
use SystemLevel  sl_macro0
timestamp 0
transform 1 0 148914 0 1 188066
box -13000 -14480 17120 18000
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 244084 74414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 244084 110414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 78000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 244084 146414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 78000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 142000 182414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 244084 182414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 244084 218414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 244084 254414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 244084 290414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 244084 326414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 244084 362414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 244084 398414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 10794 -7654 11414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 46794 -7654 47414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 46794 244084 47414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 -7654 83414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 244084 83414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 -7654 119414 78000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 142000 119414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 244084 119414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 -7654 155414 78000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 244084 155414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 -7654 191414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 244084 191414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 -7654 227414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 244084 227414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 -7654 263414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 244084 263414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 -7654 299414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 244084 299414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 -7654 335414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 244084 335414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 -7654 371414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 244084 371414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 406794 -7654 407414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 442794 -7654 443414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 478794 -7654 479414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 514794 -7654 515414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 550794 -7654 551414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 11866 592650 12486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 47866 592650 48486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 83866 592650 84486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 119866 592650 120486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 155866 592650 156486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 191866 592650 192486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 227866 592650 228486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 263866 592650 264486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 299866 592650 300486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 335866 592650 336486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 371866 592650 372486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 407866 592650 408486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 443866 592650 444486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 479866 592650 480486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 515866 592650 516486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 551866 592650 552486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 587866 592650 588486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 623866 592650 624486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 659866 592650 660486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 695866 592650 696486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 19794 -7654 20414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 55794 -7654 56414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 55794 244084 56414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 -7654 92414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 244084 92414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 -7654 128414 78000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 142000 128414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 244084 128414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 -7654 164414 78000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 244084 164414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 -7654 200414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 244084 200414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 -7654 236414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 244084 236414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 271794 -7654 272414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 271794 244084 272414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 -7654 308414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 244084 308414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 343794 -7654 344414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 343794 244084 344414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 -7654 380414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 244084 380414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 415794 -7654 416414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 451794 -7654 452414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 487794 -7654 488414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 523794 -7654 524414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 559794 -7654 560414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 20866 592650 21486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 56866 592650 57486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 92866 592650 93486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 128866 592650 129486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 164866 592650 165486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 200866 592650 201486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 236866 592650 237486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 272866 592650 273486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 308866 592650 309486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 344866 592650 345486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 380866 592650 381486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 416866 592650 417486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 452866 592650 453486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 488866 592650 489486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 524866 592650 525486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 560866 592650 561486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 596866 592650 597486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 632866 592650 633486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 668866 592650 669486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 28794 -7654 29414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 64794 -7654 65414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 64794 244084 65414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 100794 -7654 101414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 100794 244084 101414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 -7654 137414 78000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 244084 137414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 -7654 173414 78000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 142000 173414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 244084 173414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 208794 -7654 209414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 208794 244084 209414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 244794 -7654 245414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 244794 244084 245414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 280794 -7654 281414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 280794 244084 281414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 316794 -7654 317414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 316794 244084 317414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 352794 -7654 353414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 352794 244084 353414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 388794 -7654 389414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 388794 244084 389414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 424794 -7654 425414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 460794 -7654 461414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 496794 -7654 497414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 532794 -7654 533414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 568794 -7654 569414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 29866 592650 30486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 65866 592650 66486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 101866 592650 102486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 137866 592650 138486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 173866 592650 174486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 209866 592650 210486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 245866 592650 246486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 281866 592650 282486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 317866 592650 318486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 353866 592650 354486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 389866 592650 390486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 425866 592650 426486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 461866 592650 462486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 497866 592650 498486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 533866 592650 534486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 569866 592650 570486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 605866 592650 606486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 641866 592650 642486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 677866 592650 678486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 24294 -7654 24914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 60294 -7654 60914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 60294 244084 60914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 96294 -7654 96914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 96294 244084 96914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 -7654 132914 78000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 142000 132914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 244084 132914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 -7654 168914 78000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 142000 168914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 244084 168914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 204294 -7654 204914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 204294 244084 204914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 240294 -7654 240914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 240294 244084 240914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 276294 -7654 276914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 276294 244084 276914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 -7654 312914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 244084 312914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 348294 -7654 348914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 348294 244084 348914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 384294 -7654 384914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 384294 244084 384914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 420294 -7654 420914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 456294 -7654 456914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 492294 -7654 492914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 528294 -7654 528914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 564294 -7654 564914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 25366 592650 25986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 61366 592650 61986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 97366 592650 97986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 133366 592650 133986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 169366 592650 169986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 205366 592650 205986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 241366 592650 241986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 277366 592650 277986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 313366 592650 313986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 349366 592650 349986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 385366 592650 385986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 421366 592650 421986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 457366 592650 457986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 493366 592650 493986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 529366 592650 529986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 565366 592650 565986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 601366 592650 601986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 637366 592650 637986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 673366 592650 673986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 33294 -7654 33914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 69294 -7654 69914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 69294 244084 69914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 -7654 105914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 244084 105914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 -7654 141914 78000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 244084 141914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 -7654 177914 78000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 142000 177914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 244084 177914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 213294 -7654 213914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 213294 244084 213914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 -7654 249914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 244084 249914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 285294 -7654 285914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 285294 244084 285914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 321294 -7654 321914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 321294 244084 321914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 357294 -7654 357914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 357294 244084 357914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 393294 -7654 393914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 393294 244084 393914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 429294 -7654 429914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 465294 -7654 465914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 501294 -7654 501914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 537294 -7654 537914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 573294 -7654 573914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 34366 592650 34986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 70366 592650 70986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 106366 592650 106986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 142366 592650 142986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 178366 592650 178986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 214366 592650 214986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 250366 592650 250986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 286366 592650 286986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 322366 592650 322986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 358366 592650 358986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 394366 592650 394986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 430366 592650 430986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 466366 592650 466986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 502366 592650 502986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 538366 592650 538986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 574366 592650 574986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 610366 592650 610986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 646366 592650 646986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 682366 592650 682986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 6294 -7654 6914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 42294 -7654 42914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 -7654 78914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 244084 78914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 -7654 114914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 244084 114914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 -7654 150914 78000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 244084 150914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 -7654 186914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 244084 186914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 -7654 222914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 244084 222914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 -7654 258914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 244084 258914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 -7654 294914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 244084 294914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 -7654 330914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 244084 330914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 -7654 366914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 244084 366914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 402294 -7654 402914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 402294 244084 402914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 438294 -7654 438914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 474294 -7654 474914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 510294 -7654 510914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 546294 -7654 546914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 582294 -7654 582914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 7366 592650 7986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 43366 592650 43986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 79366 592650 79986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 115366 592650 115986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 151366 592650 151986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 187366 592650 187986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 223366 592650 223986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 259366 592650 259986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 295366 592650 295986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 331366 592650 331986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 367366 592650 367986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 403366 592650 403986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 439366 592650 439986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 475366 592650 475986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 511366 592650 511986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 547366 592650 547986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 583366 592650 583986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 619366 592650 619986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 655366 592650 655986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 691366 592650 691986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 15294 -7654 15914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 51294 -7654 51914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 51294 244084 51914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 -7654 87914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 244084 87914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 -7654 123914 78000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 142000 123914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 244084 123914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 -7654 159914 78000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 244084 159914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 -7654 195914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 244084 195914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 -7654 231914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 244084 231914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 -7654 267914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 244084 267914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 -7654 303914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 244084 303914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 -7654 339914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 244084 339914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 -7654 375914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 244084 375914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 411294 -7654 411914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 447294 -7654 447914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 483294 -7654 483914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 519294 -7654 519914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 555294 -7654 555914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 16366 592650 16986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 52366 592650 52986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 88366 592650 88986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 124366 592650 124986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 160366 592650 160986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 196366 592650 196986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 232366 592650 232986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 268366 592650 268986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 304366 592650 304986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 340366 592650 340986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 376366 592650 376986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 412366 592650 412986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 448366 592650 448986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 484366 592650 484986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 520366 592650 520986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 556366 592650 556986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 592366 592650 592986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 628366 592650 628986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 664366 592650 664986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 700366 592650 700986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
