magic
tech sky130B
magscale 1 2
timestamp 1667049787
<< obsli1 >>
rect 121104 82159 188816 257681
<< obsm1 >>
rect 14 2592 583082 703044
<< metal2 >>
rect 1278 703520 1390 704960
rect 5142 703520 5254 704960
rect 9006 703520 9118 704960
rect 12870 703520 12982 704960
rect 16090 703520 16202 704960
rect 19954 703520 20066 704960
rect 23818 703520 23930 704960
rect 27682 703520 27794 704960
rect 31546 703520 31658 704960
rect 35410 703520 35522 704960
rect 39274 703520 39386 704960
rect 43138 703520 43250 704960
rect 47002 703520 47114 704960
rect 50866 703520 50978 704960
rect 54730 703520 54842 704960
rect 58594 703520 58706 704960
rect 62458 703520 62570 704960
rect 66322 703520 66434 704960
rect 70186 703520 70298 704960
rect 73406 703520 73518 704960
rect 77270 703520 77382 704960
rect 81134 703520 81246 704960
rect 84998 703520 85110 704960
rect 88862 703520 88974 704960
rect 92726 703520 92838 704960
rect 96590 703520 96702 704960
rect 100454 703520 100566 704960
rect 104318 703520 104430 704960
rect 108182 703520 108294 704960
rect 112046 703520 112158 704960
rect 115910 703520 116022 704960
rect 119774 703520 119886 704960
rect 123638 703520 123750 704960
rect 127502 703520 127614 704960
rect 130722 703520 130834 704960
rect 134586 703520 134698 704960
rect 138450 703520 138562 704960
rect 142314 703520 142426 704960
rect 146178 703520 146290 704960
rect 150042 703520 150154 704960
rect 153906 703520 154018 704960
rect 157770 703520 157882 704960
rect 161634 703520 161746 704960
rect 165498 703520 165610 704960
rect 169362 703520 169474 704960
rect 173226 703520 173338 704960
rect 177090 703520 177202 704960
rect 180954 703520 181066 704960
rect 184818 703520 184930 704960
rect 188038 703520 188150 704960
rect 191902 703520 192014 704960
rect 195766 703520 195878 704960
rect 199630 703520 199742 704960
rect 203494 703520 203606 704960
rect 207358 703520 207470 704960
rect 211222 703520 211334 704960
rect 215086 703520 215198 704960
rect 218950 703520 219062 704960
rect 222814 703520 222926 704960
rect 226678 703520 226790 704960
rect 230542 703520 230654 704960
rect 234406 703520 234518 704960
rect 238270 703520 238382 704960
rect 242134 703520 242246 704960
rect 245354 703520 245466 704960
rect 249218 703520 249330 704960
rect 253082 703520 253194 704960
rect 256946 703520 257058 704960
rect 260810 703520 260922 704960
rect 264674 703520 264786 704960
rect 268538 703520 268650 704960
rect 272402 703520 272514 704960
rect 276266 703520 276378 704960
rect 280130 703520 280242 704960
rect 283994 703520 284106 704960
rect 287858 703520 287970 704960
rect 291722 703520 291834 704960
rect 295586 703520 295698 704960
rect 299450 703520 299562 704960
rect 302670 703520 302782 704960
rect 306534 703520 306646 704960
rect 310398 703520 310510 704960
rect 314262 703520 314374 704960
rect 318126 703520 318238 704960
rect 321990 703520 322102 704960
rect 325854 703520 325966 704960
rect 329718 703520 329830 704960
rect 333582 703520 333694 704960
rect 337446 703520 337558 704960
rect 341310 703520 341422 704960
rect 345174 703520 345286 704960
rect 349038 703520 349150 704960
rect 352902 703520 353014 704960
rect 356122 703520 356234 704960
rect 359986 703520 360098 704960
rect 363850 703520 363962 704960
rect 367714 703520 367826 704960
rect 371578 703520 371690 704960
rect 375442 703520 375554 704960
rect 379306 703520 379418 704960
rect 383170 703520 383282 704960
rect 387034 703520 387146 704960
rect 390898 703520 391010 704960
rect 394762 703520 394874 704960
rect 398626 703520 398738 704960
rect 402490 703520 402602 704960
rect 406354 703520 406466 704960
rect 410218 703520 410330 704960
rect 413438 703520 413550 704960
rect 417302 703520 417414 704960
rect 421166 703520 421278 704960
rect 425030 703520 425142 704960
rect 428894 703520 429006 704960
rect 432758 703520 432870 704960
rect 436622 703520 436734 704960
rect 440486 703520 440598 704960
rect 444350 703520 444462 704960
rect 448214 703520 448326 704960
rect 452078 703520 452190 704960
rect 455942 703520 456054 704960
rect 459806 703520 459918 704960
rect 463670 703520 463782 704960
rect 467534 703520 467646 704960
rect 470754 703520 470866 704960
rect 474618 703520 474730 704960
rect 478482 703520 478594 704960
rect 482346 703520 482458 704960
rect 486210 703520 486322 704960
rect 490074 703520 490186 704960
rect 493938 703520 494050 704960
rect 497802 703520 497914 704960
rect 501666 703520 501778 704960
rect 505530 703520 505642 704960
rect 509394 703520 509506 704960
rect 513258 703520 513370 704960
rect 517122 703520 517234 704960
rect 520986 703520 521098 704960
rect 524850 703520 524962 704960
rect 528070 703520 528182 704960
rect 531934 703520 532046 704960
rect 535798 703520 535910 704960
rect 539662 703520 539774 704960
rect 543526 703520 543638 704960
rect 547390 703520 547502 704960
rect 551254 703520 551366 704960
rect 555118 703520 555230 704960
rect 558982 703520 559094 704960
rect 562846 703520 562958 704960
rect 566710 703520 566822 704960
rect 570574 703520 570686 704960
rect 574438 703520 574550 704960
rect 578302 703520 578414 704960
rect 582166 703520 582278 704960
rect -10 -960 102 480
rect 3210 -960 3322 480
rect 7074 -960 7186 480
rect 10938 -960 11050 480
rect 14802 -960 14914 480
rect 18666 -960 18778 480
rect 22530 -960 22642 480
rect 26394 -960 26506 480
rect 30258 -960 30370 480
rect 34122 -960 34234 480
rect 37986 -960 38098 480
rect 41850 -960 41962 480
rect 45714 -960 45826 480
rect 49578 -960 49690 480
rect 53442 -960 53554 480
rect 56662 -960 56774 480
rect 60526 -960 60638 480
rect 64390 -960 64502 480
rect 68254 -960 68366 480
rect 72118 -960 72230 480
rect 75982 -960 76094 480
rect 79846 -960 79958 480
rect 83710 -960 83822 480
rect 87574 -960 87686 480
rect 91438 -960 91550 480
rect 95302 -960 95414 480
rect 99166 -960 99278 480
rect 103030 -960 103142 480
rect 106894 -960 107006 480
rect 110758 -960 110870 480
rect 113978 -960 114090 480
rect 117842 -960 117954 480
rect 121706 -960 121818 480
rect 125570 -960 125682 480
rect 129434 -960 129546 480
rect 133298 -960 133410 480
rect 137162 -960 137274 480
rect 141026 -960 141138 480
rect 144890 -960 145002 480
rect 148754 -960 148866 480
rect 152618 -960 152730 480
rect 156482 -960 156594 480
rect 160346 -960 160458 480
rect 164210 -960 164322 480
rect 168074 -960 168186 480
rect 171294 -960 171406 480
rect 175158 -960 175270 480
rect 179022 -960 179134 480
rect 182886 -960 182998 480
rect 186750 -960 186862 480
rect 190614 -960 190726 480
rect 194478 -960 194590 480
rect 198342 -960 198454 480
rect 202206 -960 202318 480
rect 206070 -960 206182 480
rect 209934 -960 210046 480
rect 213798 -960 213910 480
rect 217662 -960 217774 480
rect 221526 -960 221638 480
rect 225390 -960 225502 480
rect 228610 -960 228722 480
rect 232474 -960 232586 480
rect 236338 -960 236450 480
rect 240202 -960 240314 480
rect 244066 -960 244178 480
rect 247930 -960 248042 480
rect 251794 -960 251906 480
rect 255658 -960 255770 480
rect 259522 -960 259634 480
rect 263386 -960 263498 480
rect 267250 -960 267362 480
rect 271114 -960 271226 480
rect 274978 -960 275090 480
rect 278842 -960 278954 480
rect 282706 -960 282818 480
rect 285926 -960 286038 480
rect 289790 -960 289902 480
rect 293654 -960 293766 480
rect 297518 -960 297630 480
rect 301382 -960 301494 480
rect 305246 -960 305358 480
rect 309110 -960 309222 480
rect 312974 -960 313086 480
rect 316838 -960 316950 480
rect 320702 -960 320814 480
rect 324566 -960 324678 480
rect 328430 -960 328542 480
rect 332294 -960 332406 480
rect 336158 -960 336270 480
rect 340022 -960 340134 480
rect 343242 -960 343354 480
rect 347106 -960 347218 480
rect 350970 -960 351082 480
rect 354834 -960 354946 480
rect 358698 -960 358810 480
rect 362562 -960 362674 480
rect 366426 -960 366538 480
rect 370290 -960 370402 480
rect 374154 -960 374266 480
rect 378018 -960 378130 480
rect 381882 -960 381994 480
rect 385746 -960 385858 480
rect 389610 -960 389722 480
rect 393474 -960 393586 480
rect 397338 -960 397450 480
rect 400558 -960 400670 480
rect 404422 -960 404534 480
rect 408286 -960 408398 480
rect 412150 -960 412262 480
rect 416014 -960 416126 480
rect 419878 -960 419990 480
rect 423742 -960 423854 480
rect 427606 -960 427718 480
rect 431470 -960 431582 480
rect 435334 -960 435446 480
rect 439198 -960 439310 480
rect 443062 -960 443174 480
rect 446926 -960 447038 480
rect 450790 -960 450902 480
rect 454654 -960 454766 480
rect 457874 -960 457986 480
rect 461738 -960 461850 480
rect 465602 -960 465714 480
rect 469466 -960 469578 480
rect 473330 -960 473442 480
rect 477194 -960 477306 480
rect 481058 -960 481170 480
rect 484922 -960 485034 480
rect 488786 -960 488898 480
rect 492650 -960 492762 480
rect 496514 -960 496626 480
rect 500378 -960 500490 480
rect 504242 -960 504354 480
rect 508106 -960 508218 480
rect 511326 -960 511438 480
rect 515190 -960 515302 480
rect 519054 -960 519166 480
rect 522918 -960 523030 480
rect 526782 -960 526894 480
rect 530646 -960 530758 480
rect 534510 -960 534622 480
rect 538374 -960 538486 480
rect 542238 -960 542350 480
rect 546102 -960 546214 480
rect 549966 -960 550078 480
rect 553830 -960 553942 480
rect 557694 -960 557806 480
rect 561558 -960 561670 480
rect 565422 -960 565534 480
rect 568642 -960 568754 480
rect 572506 -960 572618 480
rect 576370 -960 576482 480
rect 580234 -960 580346 480
<< obsm2 >>
rect 20 703464 1222 703610
rect 1446 703464 5086 703610
rect 5310 703464 8950 703610
rect 9174 703464 12814 703610
rect 13038 703464 16034 703610
rect 16258 703464 19898 703610
rect 20122 703464 23762 703610
rect 23986 703464 27626 703610
rect 27850 703464 31490 703610
rect 31714 703464 35354 703610
rect 35578 703464 39218 703610
rect 39442 703464 43082 703610
rect 43306 703464 46946 703610
rect 47170 703464 50810 703610
rect 51034 703464 54674 703610
rect 54898 703464 58538 703610
rect 58762 703464 62402 703610
rect 62626 703464 66266 703610
rect 66490 703464 70130 703610
rect 70354 703464 73350 703610
rect 73574 703464 77214 703610
rect 77438 703464 81078 703610
rect 81302 703464 84942 703610
rect 85166 703464 88806 703610
rect 89030 703464 92670 703610
rect 92894 703464 96534 703610
rect 96758 703464 100398 703610
rect 100622 703464 104262 703610
rect 104486 703464 108126 703610
rect 108350 703464 111990 703610
rect 112214 703464 115854 703610
rect 116078 703464 119718 703610
rect 119942 703464 123582 703610
rect 123806 703464 127446 703610
rect 127670 703464 130666 703610
rect 130890 703464 134530 703610
rect 134754 703464 138394 703610
rect 138618 703464 142258 703610
rect 142482 703464 146122 703610
rect 146346 703464 149986 703610
rect 150210 703464 153850 703610
rect 154074 703464 157714 703610
rect 157938 703464 161578 703610
rect 161802 703464 165442 703610
rect 165666 703464 169306 703610
rect 169530 703464 173170 703610
rect 173394 703464 177034 703610
rect 177258 703464 180898 703610
rect 181122 703464 184762 703610
rect 184986 703464 187982 703610
rect 188206 703464 191846 703610
rect 192070 703464 195710 703610
rect 195934 703464 199574 703610
rect 199798 703464 203438 703610
rect 203662 703464 207302 703610
rect 207526 703464 211166 703610
rect 211390 703464 215030 703610
rect 215254 703464 218894 703610
rect 219118 703464 222758 703610
rect 222982 703464 226622 703610
rect 226846 703464 230486 703610
rect 230710 703464 234350 703610
rect 234574 703464 238214 703610
rect 238438 703464 242078 703610
rect 242302 703464 245298 703610
rect 245522 703464 249162 703610
rect 249386 703464 253026 703610
rect 253250 703464 256890 703610
rect 257114 703464 260754 703610
rect 260978 703464 264618 703610
rect 264842 703464 268482 703610
rect 268706 703464 272346 703610
rect 272570 703464 276210 703610
rect 276434 703464 280074 703610
rect 280298 703464 283938 703610
rect 284162 703464 287802 703610
rect 288026 703464 291666 703610
rect 291890 703464 295530 703610
rect 295754 703464 299394 703610
rect 299618 703464 302614 703610
rect 302838 703464 306478 703610
rect 306702 703464 310342 703610
rect 310566 703464 314206 703610
rect 314430 703464 318070 703610
rect 318294 703464 321934 703610
rect 322158 703464 325798 703610
rect 326022 703464 329662 703610
rect 329886 703464 333526 703610
rect 333750 703464 337390 703610
rect 337614 703464 341254 703610
rect 341478 703464 345118 703610
rect 345342 703464 348982 703610
rect 349206 703464 352846 703610
rect 353070 703464 356066 703610
rect 356290 703464 359930 703610
rect 360154 703464 363794 703610
rect 364018 703464 367658 703610
rect 367882 703464 371522 703610
rect 371746 703464 375386 703610
rect 375610 703464 379250 703610
rect 379474 703464 383114 703610
rect 383338 703464 386978 703610
rect 387202 703464 390842 703610
rect 391066 703464 394706 703610
rect 394930 703464 398570 703610
rect 398794 703464 402434 703610
rect 402658 703464 406298 703610
rect 406522 703464 410162 703610
rect 410386 703464 413382 703610
rect 413606 703464 417246 703610
rect 417470 703464 421110 703610
rect 421334 703464 424974 703610
rect 425198 703464 428838 703610
rect 429062 703464 432702 703610
rect 432926 703464 436566 703610
rect 436790 703464 440430 703610
rect 440654 703464 444294 703610
rect 444518 703464 448158 703610
rect 448382 703464 452022 703610
rect 452246 703464 455886 703610
rect 456110 703464 459750 703610
rect 459974 703464 463614 703610
rect 463838 703464 467478 703610
rect 467702 703464 470698 703610
rect 470922 703464 474562 703610
rect 474786 703464 478426 703610
rect 478650 703464 482290 703610
rect 482514 703464 486154 703610
rect 486378 703464 490018 703610
rect 490242 703464 493882 703610
rect 494106 703464 497746 703610
rect 497970 703464 501610 703610
rect 501834 703464 505474 703610
rect 505698 703464 509338 703610
rect 509562 703464 513202 703610
rect 513426 703464 517066 703610
rect 517290 703464 520930 703610
rect 521154 703464 524794 703610
rect 525018 703464 528014 703610
rect 528238 703464 531878 703610
rect 532102 703464 535742 703610
rect 535966 703464 539606 703610
rect 539830 703464 543470 703610
rect 543694 703464 547334 703610
rect 547558 703464 551198 703610
rect 551422 703464 555062 703610
rect 555286 703464 558926 703610
rect 559150 703464 562790 703610
rect 563014 703464 566654 703610
rect 566878 703464 570518 703610
rect 570742 703464 574382 703610
rect 574606 703464 578246 703610
rect 578470 703464 582110 703610
rect 582334 703464 583078 703610
rect 20 536 583078 703464
rect 158 31 3154 536
rect 3378 31 7018 536
rect 7242 31 10882 536
rect 11106 31 14746 536
rect 14970 31 18610 536
rect 18834 31 22474 536
rect 22698 31 26338 536
rect 26562 31 30202 536
rect 30426 31 34066 536
rect 34290 31 37930 536
rect 38154 31 41794 536
rect 42018 31 45658 536
rect 45882 31 49522 536
rect 49746 31 53386 536
rect 53610 31 56606 536
rect 56830 31 60470 536
rect 60694 31 64334 536
rect 64558 31 68198 536
rect 68422 31 72062 536
rect 72286 31 75926 536
rect 76150 31 79790 536
rect 80014 31 83654 536
rect 83878 31 87518 536
rect 87742 31 91382 536
rect 91606 31 95246 536
rect 95470 31 99110 536
rect 99334 31 102974 536
rect 103198 31 106838 536
rect 107062 31 110702 536
rect 110926 31 113922 536
rect 114146 31 117786 536
rect 118010 31 121650 536
rect 121874 31 125514 536
rect 125738 31 129378 536
rect 129602 31 133242 536
rect 133466 31 137106 536
rect 137330 31 140970 536
rect 141194 31 144834 536
rect 145058 31 148698 536
rect 148922 31 152562 536
rect 152786 31 156426 536
rect 156650 31 160290 536
rect 160514 31 164154 536
rect 164378 31 168018 536
rect 168242 31 171238 536
rect 171462 31 175102 536
rect 175326 31 178966 536
rect 179190 31 182830 536
rect 183054 31 186694 536
rect 186918 31 190558 536
rect 190782 31 194422 536
rect 194646 31 198286 536
rect 198510 31 202150 536
rect 202374 31 206014 536
rect 206238 31 209878 536
rect 210102 31 213742 536
rect 213966 31 217606 536
rect 217830 31 221470 536
rect 221694 31 225334 536
rect 225558 31 228554 536
rect 228778 31 232418 536
rect 232642 31 236282 536
rect 236506 31 240146 536
rect 240370 31 244010 536
rect 244234 31 247874 536
rect 248098 31 251738 536
rect 251962 31 255602 536
rect 255826 31 259466 536
rect 259690 31 263330 536
rect 263554 31 267194 536
rect 267418 31 271058 536
rect 271282 31 274922 536
rect 275146 31 278786 536
rect 279010 31 282650 536
rect 282874 31 285870 536
rect 286094 31 289734 536
rect 289958 31 293598 536
rect 293822 31 297462 536
rect 297686 31 301326 536
rect 301550 31 305190 536
rect 305414 31 309054 536
rect 309278 31 312918 536
rect 313142 31 316782 536
rect 317006 31 320646 536
rect 320870 31 324510 536
rect 324734 31 328374 536
rect 328598 31 332238 536
rect 332462 31 336102 536
rect 336326 31 339966 536
rect 340190 31 343186 536
rect 343410 31 347050 536
rect 347274 31 350914 536
rect 351138 31 354778 536
rect 355002 31 358642 536
rect 358866 31 362506 536
rect 362730 31 366370 536
rect 366594 31 370234 536
rect 370458 31 374098 536
rect 374322 31 377962 536
rect 378186 31 381826 536
rect 382050 31 385690 536
rect 385914 31 389554 536
rect 389778 31 393418 536
rect 393642 31 397282 536
rect 397506 31 400502 536
rect 400726 31 404366 536
rect 404590 31 408230 536
rect 408454 31 412094 536
rect 412318 31 415958 536
rect 416182 31 419822 536
rect 420046 31 423686 536
rect 423910 31 427550 536
rect 427774 31 431414 536
rect 431638 31 435278 536
rect 435502 31 439142 536
rect 439366 31 443006 536
rect 443230 31 446870 536
rect 447094 31 450734 536
rect 450958 31 454598 536
rect 454822 31 457818 536
rect 458042 31 461682 536
rect 461906 31 465546 536
rect 465770 31 469410 536
rect 469634 31 473274 536
rect 473498 31 477138 536
rect 477362 31 481002 536
rect 481226 31 484866 536
rect 485090 31 488730 536
rect 488954 31 492594 536
rect 492818 31 496458 536
rect 496682 31 500322 536
rect 500546 31 504186 536
rect 504410 31 508050 536
rect 508274 31 511270 536
rect 511494 31 515134 536
rect 515358 31 518998 536
rect 519222 31 522862 536
rect 523086 31 526726 536
rect 526950 31 530590 536
rect 530814 31 534454 536
rect 534678 31 538318 536
rect 538542 31 542182 536
rect 542406 31 546046 536
rect 546270 31 549910 536
rect 550134 31 553774 536
rect 553998 31 557638 536
rect 557862 31 561502 536
rect 561726 31 565366 536
rect 565590 31 568586 536
rect 568810 31 572450 536
rect 572674 31 576314 536
rect 576538 31 580178 536
rect 580402 31 583078 536
<< metal3 >>
rect 583520 702388 584960 702628
rect -960 701708 480 701948
rect 583520 698308 584960 698548
rect -960 697628 480 697868
rect 583520 694228 584960 694468
rect -960 693548 480 693788
rect 583520 690148 584960 690388
rect -960 689468 480 689708
rect 583520 686068 584960 686308
rect -960 685388 480 685628
rect 583520 681988 584960 682228
rect -960 681308 480 681548
rect 583520 677908 584960 678148
rect -960 677228 480 677468
rect 583520 673828 584960 674068
rect -960 673148 480 673388
rect 583520 669748 584960 669988
rect -960 669068 480 669308
rect 583520 665668 584960 665908
rect -960 664988 480 665228
rect 583520 661588 584960 661828
rect -960 660908 480 661148
rect -960 657508 480 657748
rect 583520 657508 584960 657748
rect -960 653428 480 653668
rect 583520 653428 584960 653668
rect -960 649348 480 649588
rect 583520 649348 584960 649588
rect -960 645268 480 645508
rect 583520 645268 584960 645508
rect 583520 641868 584960 642108
rect -960 641188 480 641428
rect 583520 637788 584960 638028
rect -960 637108 480 637348
rect 583520 633708 584960 633948
rect -960 633028 480 633268
rect 583520 629628 584960 629868
rect -960 628948 480 629188
rect 583520 625548 584960 625788
rect -960 624868 480 625108
rect 583520 621468 584960 621708
rect -960 620788 480 621028
rect 583520 617388 584960 617628
rect -960 616708 480 616948
rect 583520 613308 584960 613548
rect -960 612628 480 612868
rect 583520 609228 584960 609468
rect -960 608548 480 608788
rect 583520 605148 584960 605388
rect -960 604468 480 604708
rect 583520 601068 584960 601308
rect -960 600388 480 600628
rect -960 596988 480 597228
rect 583520 596988 584960 597228
rect -960 592908 480 593148
rect 583520 592908 584960 593148
rect -960 588828 480 589068
rect 583520 588828 584960 589068
rect -960 584748 480 584988
rect 583520 584748 584960 584988
rect 583520 581348 584960 581588
rect -960 580668 480 580908
rect 583520 577268 584960 577508
rect -960 576588 480 576828
rect 583520 573188 584960 573428
rect -960 572508 480 572748
rect 583520 569108 584960 569348
rect -960 568428 480 568668
rect 583520 565028 584960 565268
rect -960 564348 480 564588
rect 583520 560948 584960 561188
rect -960 560268 480 560508
rect 583520 556868 584960 557108
rect -960 556188 480 556428
rect 583520 552788 584960 553028
rect -960 552108 480 552348
rect 583520 548708 584960 548948
rect -960 548028 480 548268
rect 583520 544628 584960 544868
rect -960 543948 480 544188
rect 583520 540548 584960 540788
rect -960 539868 480 540108
rect -960 536468 480 536708
rect 583520 536468 584960 536708
rect -960 532388 480 532628
rect 583520 532388 584960 532628
rect -960 528308 480 528548
rect 583520 528308 584960 528548
rect -960 524228 480 524468
rect 583520 524228 584960 524468
rect 583520 520828 584960 521068
rect -960 520148 480 520388
rect 583520 516748 584960 516988
rect -960 516068 480 516308
rect 583520 512668 584960 512908
rect -960 511988 480 512228
rect 583520 508588 584960 508828
rect -960 507908 480 508148
rect 583520 504508 584960 504748
rect -960 503828 480 504068
rect 583520 500428 584960 500668
rect -960 499748 480 499988
rect 583520 496348 584960 496588
rect -960 495668 480 495908
rect 583520 492268 584960 492508
rect -960 491588 480 491828
rect 583520 488188 584960 488428
rect -960 487508 480 487748
rect 583520 484108 584960 484348
rect -960 483428 480 483668
rect -960 480028 480 480268
rect 583520 480028 584960 480268
rect -960 475948 480 476188
rect 583520 475948 584960 476188
rect -960 471868 480 472108
rect 583520 471868 584960 472108
rect -960 467788 480 468028
rect 583520 467788 584960 468028
rect -960 463708 480 463948
rect 583520 463708 584960 463948
rect 583520 460308 584960 460548
rect -960 459628 480 459868
rect 583520 456228 584960 456468
rect -960 455548 480 455788
rect 583520 452148 584960 452388
rect -960 451468 480 451708
rect 583520 448068 584960 448308
rect -960 447388 480 447628
rect 583520 443988 584960 444228
rect -960 443308 480 443548
rect 583520 439908 584960 440148
rect -960 439228 480 439468
rect 583520 435828 584960 436068
rect -960 435148 480 435388
rect 583520 431748 584960 431988
rect -960 431068 480 431308
rect 583520 427668 584960 427908
rect -960 426988 480 427228
rect 583520 423588 584960 423828
rect -960 422908 480 423148
rect -960 419508 480 419748
rect 583520 419508 584960 419748
rect -960 415428 480 415668
rect 583520 415428 584960 415668
rect -960 411348 480 411588
rect 583520 411348 584960 411588
rect -960 407268 480 407508
rect 583520 407268 584960 407508
rect 583520 403868 584960 404108
rect -960 403188 480 403428
rect 583520 399788 584960 400028
rect -960 399108 480 399348
rect 583520 395708 584960 395948
rect -960 395028 480 395268
rect 583520 391628 584960 391868
rect -960 390948 480 391188
rect 583520 387548 584960 387788
rect -960 386868 480 387108
rect 583520 383468 584960 383708
rect -960 382788 480 383028
rect 583520 379388 584960 379628
rect -960 378708 480 378948
rect 583520 375308 584960 375548
rect -960 374628 480 374868
rect 583520 371228 584960 371468
rect -960 370548 480 370788
rect 583520 367148 584960 367388
rect -960 366468 480 366708
rect 583520 363068 584960 363308
rect -960 362388 480 362628
rect -960 358988 480 359228
rect 583520 358988 584960 359228
rect -960 354908 480 355148
rect 583520 354908 584960 355148
rect -960 350828 480 351068
rect 583520 350828 584960 351068
rect -960 346748 480 346988
rect 583520 346748 584960 346988
rect 583520 343348 584960 343588
rect -960 342668 480 342908
rect 583520 339268 584960 339508
rect -960 338588 480 338828
rect 583520 335188 584960 335428
rect -960 334508 480 334748
rect 583520 331108 584960 331348
rect -960 330428 480 330668
rect 583520 327028 584960 327268
rect -960 326348 480 326588
rect 583520 322948 584960 323188
rect -960 322268 480 322508
rect 583520 318868 584960 319108
rect -960 318188 480 318428
rect 583520 314788 584960 315028
rect -960 314108 480 314348
rect 583520 310708 584960 310948
rect -960 310028 480 310268
rect 583520 306628 584960 306868
rect -960 305948 480 306188
rect 583520 302548 584960 302788
rect -960 301868 480 302108
rect -960 298468 480 298708
rect 583520 298468 584960 298708
rect -960 294388 480 294628
rect 583520 294388 584960 294628
rect -960 290308 480 290548
rect 583520 290308 584960 290548
rect -960 286228 480 286468
rect 583520 286228 584960 286468
rect 583520 282828 584960 283068
rect -960 282148 480 282388
rect 583520 278748 584960 278988
rect -960 278068 480 278308
rect 583520 274668 584960 274908
rect -960 273988 480 274228
rect 583520 270588 584960 270828
rect -960 269908 480 270148
rect 583520 266508 584960 266748
rect -960 265828 480 266068
rect 583520 262428 584960 262668
rect -960 261748 480 261988
rect 583520 258348 584960 258588
rect -960 257668 480 257908
rect 583520 254268 584960 254508
rect -960 253588 480 253828
rect 583520 250188 584960 250428
rect -960 249508 480 249748
rect 583520 246108 584960 246348
rect -960 245428 480 245668
rect 583520 242028 584960 242268
rect -960 241348 480 241588
rect -960 237948 480 238188
rect 583520 237948 584960 238188
rect -960 233868 480 234108
rect 583520 233868 584960 234108
rect -960 229788 480 230028
rect 583520 229788 584960 230028
rect -960 225708 480 225948
rect 583520 225708 584960 225948
rect 583520 222308 584960 222548
rect -960 221628 480 221868
rect 583520 218228 584960 218468
rect -960 217548 480 217788
rect 583520 214148 584960 214388
rect -960 213468 480 213708
rect 583520 210068 584960 210308
rect -960 209388 480 209628
rect 583520 205988 584960 206228
rect -960 205308 480 205548
rect 583520 201908 584960 202148
rect -960 201228 480 201468
rect 583520 197828 584960 198068
rect -960 197148 480 197388
rect 583520 193748 584960 193988
rect -960 193068 480 193308
rect 583520 189668 584960 189908
rect -960 188988 480 189228
rect 583520 185588 584960 185828
rect -960 184908 480 185148
rect 583520 181508 584960 181748
rect -960 180828 480 181068
rect -960 177428 480 177668
rect 583520 177428 584960 177668
rect -960 173348 480 173588
rect 583520 173348 584960 173588
rect -960 169268 480 169508
rect 583520 169268 584960 169508
rect -960 165188 480 165428
rect 583520 165188 584960 165428
rect 583520 161788 584960 162028
rect -960 161108 480 161348
rect 583520 157708 584960 157948
rect -960 157028 480 157268
rect 583520 153628 584960 153868
rect -960 152948 480 153188
rect 583520 149548 584960 149788
rect -960 148868 480 149108
rect 583520 145468 584960 145708
rect -960 144788 480 145028
rect 583520 141388 584960 141628
rect -960 140708 480 140948
rect 583520 137308 584960 137548
rect -960 136628 480 136868
rect 583520 133228 584960 133468
rect -960 132548 480 132788
rect 583520 129148 584960 129388
rect -960 128468 480 128708
rect 583520 125068 584960 125308
rect -960 124388 480 124628
rect 583520 120988 584960 121228
rect -960 120308 480 120548
rect -960 116908 480 117148
rect 583520 116908 584960 117148
rect -960 112828 480 113068
rect 583520 112828 584960 113068
rect -960 108748 480 108988
rect 583520 108748 584960 108988
rect -960 104668 480 104908
rect 583520 104668 584960 104908
rect 583520 101268 584960 101508
rect -960 100588 480 100828
rect 583520 97188 584960 97428
rect -960 96508 480 96748
rect 583520 93108 584960 93348
rect -960 92428 480 92668
rect 583520 89028 584960 89268
rect -960 88348 480 88588
rect 583520 84948 584960 85188
rect -960 84268 480 84508
rect 583520 80868 584960 81108
rect -960 80188 480 80428
rect 583520 76788 584960 77028
rect -960 76108 480 76348
rect 583520 72708 584960 72948
rect -960 72028 480 72268
rect 583520 68628 584960 68868
rect -960 67948 480 68188
rect 583520 64548 584960 64788
rect -960 63868 480 64108
rect 583520 60468 584960 60708
rect -960 59788 480 60028
rect -960 56388 480 56628
rect 583520 56388 584960 56628
rect -960 52308 480 52548
rect 583520 52308 584960 52548
rect -960 48228 480 48468
rect 583520 48228 584960 48468
rect -960 44148 480 44388
rect 583520 44148 584960 44388
rect 583520 40748 584960 40988
rect -960 40068 480 40308
rect 583520 36668 584960 36908
rect -960 35988 480 36228
rect 583520 32588 584960 32828
rect -960 31908 480 32148
rect 583520 28508 584960 28748
rect -960 27828 480 28068
rect 583520 24428 584960 24668
rect -960 23748 480 23988
rect 583520 20348 584960 20588
rect -960 19668 480 19908
rect 583520 16268 584960 16508
rect -960 15588 480 15828
rect 583520 12188 584960 12428
rect -960 11508 480 11748
rect 583520 8108 584960 8348
rect -960 7428 480 7668
rect 583520 4028 584960 4268
rect -960 3348 480 3588
rect 583520 -52 584960 188
<< obsm3 >>
rect 246 702308 583440 702541
rect 246 702028 583586 702308
rect 560 701628 583586 702028
rect 246 698628 583586 701628
rect 246 698228 583440 698628
rect 246 697948 583586 698228
rect 560 697548 583586 697948
rect 246 694548 583586 697548
rect 246 694148 583440 694548
rect 246 693868 583586 694148
rect 560 693468 583586 693868
rect 246 690468 583586 693468
rect 246 690068 583440 690468
rect 246 689788 583586 690068
rect 560 689388 583586 689788
rect 246 686388 583586 689388
rect 246 685988 583440 686388
rect 246 685708 583586 685988
rect 560 685308 583586 685708
rect 246 682308 583586 685308
rect 246 681908 583440 682308
rect 246 681628 583586 681908
rect 560 681228 583586 681628
rect 246 678228 583586 681228
rect 246 677828 583440 678228
rect 246 677548 583586 677828
rect 560 677148 583586 677548
rect 246 674148 583586 677148
rect 246 673748 583440 674148
rect 246 673468 583586 673748
rect 560 673068 583586 673468
rect 246 670068 583586 673068
rect 246 669668 583440 670068
rect 246 669388 583586 669668
rect 560 668988 583586 669388
rect 246 665988 583586 668988
rect 246 665588 583440 665988
rect 246 665308 583586 665588
rect 560 664908 583586 665308
rect 246 661908 583586 664908
rect 246 661508 583440 661908
rect 246 661228 583586 661508
rect 560 660828 583586 661228
rect 246 657828 583586 660828
rect 560 657428 583440 657828
rect 246 653748 583586 657428
rect 560 653348 583440 653748
rect 246 649668 583586 653348
rect 560 649268 583440 649668
rect 246 645588 583586 649268
rect 560 645188 583440 645588
rect 246 642188 583586 645188
rect 246 641788 583440 642188
rect 246 641508 583586 641788
rect 560 641108 583586 641508
rect 246 638108 583586 641108
rect 246 637708 583440 638108
rect 246 637428 583586 637708
rect 560 637028 583586 637428
rect 246 634028 583586 637028
rect 246 633628 583440 634028
rect 246 633348 583586 633628
rect 560 632948 583586 633348
rect 246 629948 583586 632948
rect 246 629548 583440 629948
rect 246 629268 583586 629548
rect 560 628868 583586 629268
rect 246 625868 583586 628868
rect 246 625468 583440 625868
rect 246 625188 583586 625468
rect 560 624788 583586 625188
rect 246 621788 583586 624788
rect 246 621388 583440 621788
rect 246 621108 583586 621388
rect 560 620708 583586 621108
rect 246 617708 583586 620708
rect 246 617308 583440 617708
rect 246 617028 583586 617308
rect 560 616628 583586 617028
rect 246 613628 583586 616628
rect 246 613228 583440 613628
rect 246 612948 583586 613228
rect 560 612548 583586 612948
rect 246 609548 583586 612548
rect 246 609148 583440 609548
rect 246 608868 583586 609148
rect 560 608468 583586 608868
rect 246 605468 583586 608468
rect 246 605068 583440 605468
rect 246 604788 583586 605068
rect 560 604388 583586 604788
rect 246 601388 583586 604388
rect 246 600988 583440 601388
rect 246 600708 583586 600988
rect 560 600308 583586 600708
rect 246 597308 583586 600308
rect 560 596908 583440 597308
rect 246 593228 583586 596908
rect 560 592828 583440 593228
rect 246 589148 583586 592828
rect 560 588748 583440 589148
rect 246 585068 583586 588748
rect 560 584668 583440 585068
rect 246 581668 583586 584668
rect 246 581268 583440 581668
rect 246 580988 583586 581268
rect 560 580588 583586 580988
rect 246 577588 583586 580588
rect 246 577188 583440 577588
rect 246 576908 583586 577188
rect 560 576508 583586 576908
rect 246 573508 583586 576508
rect 246 573108 583440 573508
rect 246 572828 583586 573108
rect 560 572428 583586 572828
rect 246 569428 583586 572428
rect 246 569028 583440 569428
rect 246 568748 583586 569028
rect 560 568348 583586 568748
rect 246 565348 583586 568348
rect 246 564948 583440 565348
rect 246 564668 583586 564948
rect 560 564268 583586 564668
rect 246 561268 583586 564268
rect 246 560868 583440 561268
rect 246 560588 583586 560868
rect 560 560188 583586 560588
rect 246 557188 583586 560188
rect 246 556788 583440 557188
rect 246 556508 583586 556788
rect 560 556108 583586 556508
rect 246 553108 583586 556108
rect 246 552708 583440 553108
rect 246 552428 583586 552708
rect 560 552028 583586 552428
rect 246 549028 583586 552028
rect 246 548628 583440 549028
rect 246 548348 583586 548628
rect 560 547948 583586 548348
rect 246 544948 583586 547948
rect 246 544548 583440 544948
rect 246 544268 583586 544548
rect 560 543868 583586 544268
rect 246 540868 583586 543868
rect 246 540468 583440 540868
rect 246 540188 583586 540468
rect 560 539788 583586 540188
rect 246 536788 583586 539788
rect 560 536388 583440 536788
rect 246 532708 583586 536388
rect 560 532308 583440 532708
rect 246 528628 583586 532308
rect 560 528228 583440 528628
rect 246 524548 583586 528228
rect 560 524148 583440 524548
rect 246 521148 583586 524148
rect 246 520748 583440 521148
rect 246 520468 583586 520748
rect 560 520068 583586 520468
rect 246 517068 583586 520068
rect 246 516668 583440 517068
rect 246 516388 583586 516668
rect 560 515988 583586 516388
rect 246 512988 583586 515988
rect 246 512588 583440 512988
rect 246 512308 583586 512588
rect 560 511908 583586 512308
rect 246 508908 583586 511908
rect 246 508508 583440 508908
rect 246 508228 583586 508508
rect 560 507828 583586 508228
rect 246 504828 583586 507828
rect 246 504428 583440 504828
rect 246 504148 583586 504428
rect 560 503748 583586 504148
rect 246 500748 583586 503748
rect 246 500348 583440 500748
rect 246 500068 583586 500348
rect 560 499668 583586 500068
rect 246 496668 583586 499668
rect 246 496268 583440 496668
rect 246 495988 583586 496268
rect 560 495588 583586 495988
rect 246 492588 583586 495588
rect 246 492188 583440 492588
rect 246 491908 583586 492188
rect 560 491508 583586 491908
rect 246 488508 583586 491508
rect 246 488108 583440 488508
rect 246 487828 583586 488108
rect 560 487428 583586 487828
rect 246 484428 583586 487428
rect 246 484028 583440 484428
rect 246 483748 583586 484028
rect 560 483348 583586 483748
rect 246 480348 583586 483348
rect 560 479948 583440 480348
rect 246 476268 583586 479948
rect 560 475868 583440 476268
rect 246 472188 583586 475868
rect 560 471788 583440 472188
rect 246 468108 583586 471788
rect 560 467708 583440 468108
rect 246 464028 583586 467708
rect 560 463628 583440 464028
rect 246 460628 583586 463628
rect 246 460228 583440 460628
rect 246 459948 583586 460228
rect 560 459548 583586 459948
rect 246 456548 583586 459548
rect 246 456148 583440 456548
rect 246 455868 583586 456148
rect 560 455468 583586 455868
rect 246 452468 583586 455468
rect 246 452068 583440 452468
rect 246 451788 583586 452068
rect 560 451388 583586 451788
rect 246 448388 583586 451388
rect 246 447988 583440 448388
rect 246 447708 583586 447988
rect 560 447308 583586 447708
rect 246 444308 583586 447308
rect 246 443908 583440 444308
rect 246 443628 583586 443908
rect 560 443228 583586 443628
rect 246 440228 583586 443228
rect 246 439828 583440 440228
rect 246 439548 583586 439828
rect 560 439148 583586 439548
rect 246 436148 583586 439148
rect 246 435748 583440 436148
rect 246 435468 583586 435748
rect 560 435068 583586 435468
rect 246 432068 583586 435068
rect 246 431668 583440 432068
rect 246 431388 583586 431668
rect 560 430988 583586 431388
rect 246 427988 583586 430988
rect 246 427588 583440 427988
rect 246 427308 583586 427588
rect 560 426908 583586 427308
rect 246 423908 583586 426908
rect 246 423508 583440 423908
rect 246 423228 583586 423508
rect 560 422828 583586 423228
rect 246 419828 583586 422828
rect 560 419428 583440 419828
rect 246 415748 583586 419428
rect 560 415348 583440 415748
rect 246 411668 583586 415348
rect 560 411268 583440 411668
rect 246 407588 583586 411268
rect 560 407188 583440 407588
rect 246 404188 583586 407188
rect 246 403788 583440 404188
rect 246 403508 583586 403788
rect 560 403108 583586 403508
rect 246 400108 583586 403108
rect 246 399708 583440 400108
rect 246 399428 583586 399708
rect 560 399028 583586 399428
rect 246 396028 583586 399028
rect 246 395628 583440 396028
rect 246 395348 583586 395628
rect 560 394948 583586 395348
rect 246 391948 583586 394948
rect 246 391548 583440 391948
rect 246 391268 583586 391548
rect 560 390868 583586 391268
rect 246 387868 583586 390868
rect 246 387468 583440 387868
rect 246 387188 583586 387468
rect 560 386788 583586 387188
rect 246 383788 583586 386788
rect 246 383388 583440 383788
rect 246 383108 583586 383388
rect 560 382708 583586 383108
rect 246 379708 583586 382708
rect 246 379308 583440 379708
rect 246 379028 583586 379308
rect 560 378628 583586 379028
rect 246 375628 583586 378628
rect 246 375228 583440 375628
rect 246 374948 583586 375228
rect 560 374548 583586 374948
rect 246 371548 583586 374548
rect 246 371148 583440 371548
rect 246 370868 583586 371148
rect 560 370468 583586 370868
rect 246 367468 583586 370468
rect 246 367068 583440 367468
rect 246 366788 583586 367068
rect 560 366388 583586 366788
rect 246 363388 583586 366388
rect 246 362988 583440 363388
rect 246 362708 583586 362988
rect 560 362308 583586 362708
rect 246 359308 583586 362308
rect 560 358908 583440 359308
rect 246 355228 583586 358908
rect 560 354828 583440 355228
rect 246 351148 583586 354828
rect 560 350748 583440 351148
rect 246 347068 583586 350748
rect 560 346668 583440 347068
rect 246 343668 583586 346668
rect 246 343268 583440 343668
rect 246 342988 583586 343268
rect 560 342588 583586 342988
rect 246 339588 583586 342588
rect 246 339188 583440 339588
rect 246 338908 583586 339188
rect 560 338508 583586 338908
rect 246 335508 583586 338508
rect 246 335108 583440 335508
rect 246 334828 583586 335108
rect 560 334428 583586 334828
rect 246 331428 583586 334428
rect 246 331028 583440 331428
rect 246 330748 583586 331028
rect 560 330348 583586 330748
rect 246 327348 583586 330348
rect 246 326948 583440 327348
rect 246 326668 583586 326948
rect 560 326268 583586 326668
rect 246 323268 583586 326268
rect 246 322868 583440 323268
rect 246 322588 583586 322868
rect 560 322188 583586 322588
rect 246 319188 583586 322188
rect 246 318788 583440 319188
rect 246 318508 583586 318788
rect 560 318108 583586 318508
rect 246 315108 583586 318108
rect 246 314708 583440 315108
rect 246 314428 583586 314708
rect 560 314028 583586 314428
rect 246 311028 583586 314028
rect 246 310628 583440 311028
rect 246 310348 583586 310628
rect 560 309948 583586 310348
rect 246 306948 583586 309948
rect 246 306548 583440 306948
rect 246 306268 583586 306548
rect 560 305868 583586 306268
rect 246 302868 583586 305868
rect 246 302468 583440 302868
rect 246 302188 583586 302468
rect 560 301788 583586 302188
rect 246 298788 583586 301788
rect 560 298388 583440 298788
rect 246 294708 583586 298388
rect 560 294308 583440 294708
rect 246 290628 583586 294308
rect 560 290228 583440 290628
rect 246 286548 583586 290228
rect 560 286148 583440 286548
rect 246 283148 583586 286148
rect 246 282748 583440 283148
rect 246 282468 583586 282748
rect 560 282068 583586 282468
rect 246 279068 583586 282068
rect 246 278668 583440 279068
rect 246 278388 583586 278668
rect 560 277988 583586 278388
rect 246 274988 583586 277988
rect 246 274588 583440 274988
rect 246 274308 583586 274588
rect 560 273908 583586 274308
rect 246 270908 583586 273908
rect 246 270508 583440 270908
rect 246 270228 583586 270508
rect 560 269828 583586 270228
rect 246 266828 583586 269828
rect 246 266428 583440 266828
rect 246 266148 583586 266428
rect 560 265748 583586 266148
rect 246 262748 583586 265748
rect 246 262348 583440 262748
rect 246 262068 583586 262348
rect 560 261668 583586 262068
rect 246 258668 583586 261668
rect 246 258268 583440 258668
rect 246 257988 583586 258268
rect 560 257588 583586 257988
rect 246 254588 583586 257588
rect 246 254188 583440 254588
rect 246 253908 583586 254188
rect 560 253508 583586 253908
rect 246 250508 583586 253508
rect 246 250108 583440 250508
rect 246 249828 583586 250108
rect 560 249428 583586 249828
rect 246 246428 583586 249428
rect 246 246028 583440 246428
rect 246 245748 583586 246028
rect 560 245348 583586 245748
rect 246 242348 583586 245348
rect 246 241948 583440 242348
rect 246 241668 583586 241948
rect 560 241268 583586 241668
rect 246 238268 583586 241268
rect 560 237868 583440 238268
rect 246 234188 583586 237868
rect 560 233788 583440 234188
rect 246 230108 583586 233788
rect 560 229708 583440 230108
rect 246 226028 583586 229708
rect 560 225628 583440 226028
rect 246 222628 583586 225628
rect 246 222228 583440 222628
rect 246 221948 583586 222228
rect 560 221548 583586 221948
rect 246 218548 583586 221548
rect 246 218148 583440 218548
rect 246 217868 583586 218148
rect 560 217468 583586 217868
rect 246 214468 583586 217468
rect 246 214068 583440 214468
rect 246 213788 583586 214068
rect 560 213388 583586 213788
rect 246 210388 583586 213388
rect 246 209988 583440 210388
rect 246 209708 583586 209988
rect 560 209308 583586 209708
rect 246 206308 583586 209308
rect 246 205908 583440 206308
rect 246 205628 583586 205908
rect 560 205228 583586 205628
rect 246 202228 583586 205228
rect 246 201828 583440 202228
rect 246 201548 583586 201828
rect 560 201148 583586 201548
rect 246 198148 583586 201148
rect 246 197748 583440 198148
rect 246 197468 583586 197748
rect 560 197068 583586 197468
rect 246 194068 583586 197068
rect 246 193668 583440 194068
rect 246 193388 583586 193668
rect 560 192988 583586 193388
rect 246 189988 583586 192988
rect 246 189588 583440 189988
rect 246 189308 583586 189588
rect 560 188908 583586 189308
rect 246 185908 583586 188908
rect 246 185508 583440 185908
rect 246 185228 583586 185508
rect 560 184828 583586 185228
rect 246 181828 583586 184828
rect 246 181428 583440 181828
rect 246 181148 583586 181428
rect 560 180748 583586 181148
rect 246 177748 583586 180748
rect 560 177348 583440 177748
rect 246 173668 583586 177348
rect 560 173268 583440 173668
rect 246 169588 583586 173268
rect 560 169188 583440 169588
rect 246 165508 583586 169188
rect 560 165108 583440 165508
rect 246 162108 583586 165108
rect 246 161708 583440 162108
rect 246 161428 583586 161708
rect 560 161028 583586 161428
rect 246 158028 583586 161028
rect 246 157628 583440 158028
rect 246 157348 583586 157628
rect 560 156948 583586 157348
rect 246 153948 583586 156948
rect 246 153548 583440 153948
rect 246 153268 583586 153548
rect 560 152868 583586 153268
rect 246 149868 583586 152868
rect 246 149468 583440 149868
rect 246 149188 583586 149468
rect 560 148788 583586 149188
rect 246 145788 583586 148788
rect 246 145388 583440 145788
rect 246 145108 583586 145388
rect 560 144708 583586 145108
rect 246 141708 583586 144708
rect 246 141308 583440 141708
rect 246 141028 583586 141308
rect 560 140628 583586 141028
rect 246 137628 583586 140628
rect 246 137228 583440 137628
rect 246 136948 583586 137228
rect 560 136548 583586 136948
rect 246 133548 583586 136548
rect 246 133148 583440 133548
rect 246 132868 583586 133148
rect 560 132468 583586 132868
rect 246 129468 583586 132468
rect 246 129068 583440 129468
rect 246 128788 583586 129068
rect 560 128388 583586 128788
rect 246 125388 583586 128388
rect 246 124988 583440 125388
rect 246 124708 583586 124988
rect 560 124308 583586 124708
rect 246 121308 583586 124308
rect 246 120908 583440 121308
rect 246 120628 583586 120908
rect 560 120228 583586 120628
rect 246 117228 583586 120228
rect 560 116828 583440 117228
rect 246 113148 583586 116828
rect 560 112748 583440 113148
rect 246 109068 583586 112748
rect 560 108668 583440 109068
rect 246 104988 583586 108668
rect 560 104588 583440 104988
rect 246 101588 583586 104588
rect 246 101188 583440 101588
rect 246 100908 583586 101188
rect 560 100508 583586 100908
rect 246 97508 583586 100508
rect 246 97108 583440 97508
rect 246 96828 583586 97108
rect 560 96428 583586 96828
rect 246 93428 583586 96428
rect 246 93028 583440 93428
rect 246 92748 583586 93028
rect 560 92348 583586 92748
rect 246 89348 583586 92348
rect 246 88948 583440 89348
rect 246 88668 583586 88948
rect 560 88268 583586 88668
rect 246 85268 583586 88268
rect 246 84868 583440 85268
rect 246 84588 583586 84868
rect 560 84188 583586 84588
rect 246 81188 583586 84188
rect 246 80788 583440 81188
rect 246 80508 583586 80788
rect 560 80108 583586 80508
rect 246 77108 583586 80108
rect 246 76708 583440 77108
rect 246 76428 583586 76708
rect 560 76028 583586 76428
rect 246 73028 583586 76028
rect 246 72628 583440 73028
rect 246 72348 583586 72628
rect 560 71948 583586 72348
rect 246 68948 583586 71948
rect 246 68548 583440 68948
rect 246 68268 583586 68548
rect 560 67868 583586 68268
rect 246 64868 583586 67868
rect 246 64468 583440 64868
rect 246 64188 583586 64468
rect 560 63788 583586 64188
rect 246 60788 583586 63788
rect 246 60388 583440 60788
rect 246 60108 583586 60388
rect 560 59708 583586 60108
rect 246 56708 583586 59708
rect 560 56308 583440 56708
rect 246 52628 583586 56308
rect 560 52228 583440 52628
rect 246 48548 583586 52228
rect 560 48148 583440 48548
rect 246 44468 583586 48148
rect 560 44068 583440 44468
rect 246 41068 583586 44068
rect 246 40668 583440 41068
rect 246 40388 583586 40668
rect 560 39988 583586 40388
rect 246 36988 583586 39988
rect 246 36588 583440 36988
rect 246 36308 583586 36588
rect 560 35908 583586 36308
rect 246 32908 583586 35908
rect 246 32508 583440 32908
rect 246 32228 583586 32508
rect 560 31828 583586 32228
rect 246 28828 583586 31828
rect 246 28428 583440 28828
rect 246 28148 583586 28428
rect 560 27748 583586 28148
rect 246 24748 583586 27748
rect 246 24348 583440 24748
rect 246 24068 583586 24348
rect 560 23668 583586 24068
rect 246 20668 583586 23668
rect 246 20268 583440 20668
rect 246 19988 583586 20268
rect 560 19588 583586 19988
rect 246 16588 583586 19588
rect 246 16188 583440 16588
rect 246 15908 583586 16188
rect 560 15508 583586 15908
rect 246 12508 583586 15508
rect 246 12108 583440 12508
rect 246 11828 583586 12108
rect 560 11428 583586 11828
rect 246 8428 583586 11428
rect 246 8028 583440 8428
rect 246 7748 583586 8028
rect 560 7348 583586 7748
rect 246 4348 583586 7348
rect 246 3948 583440 4348
rect 246 3668 583586 3948
rect 560 3268 583586 3668
rect 246 268 583586 3268
rect 246 35 583440 268
<< metal4 >>
rect -8726 -7654 -8106 711590
rect -7766 -6694 -7146 710630
rect -6806 -5734 -6186 709670
rect -5846 -4774 -5226 708710
rect -4886 -3814 -4266 707750
rect -3926 -2854 -3306 706790
rect -2966 -1894 -2346 705830
rect -2006 -934 -1386 704870
rect 1794 -7654 2414 711590
rect 6294 -7654 6914 711590
rect 10794 -7654 11414 711590
rect 15294 -7654 15914 711590
rect 19794 -7654 20414 711590
rect 24294 -7654 24914 711590
rect 28794 -7654 29414 711590
rect 33294 -7654 33914 711590
rect 37794 -7654 38414 711590
rect 42294 -7654 42914 711590
rect 46794 -7654 47414 711590
rect 51294 -7654 51914 711590
rect 55794 -7654 56414 711590
rect 60294 -7654 60914 711590
rect 64794 -7654 65414 711590
rect 69294 -7654 69914 711590
rect 73794 -7654 74414 711590
rect 78294 -7654 78914 711590
rect 82794 -7654 83414 711590
rect 87294 -7654 87914 711590
rect 91794 -7654 92414 711590
rect 96294 -7654 96914 711590
rect 100794 -7654 101414 711590
rect 105294 -7654 105914 711590
rect 109794 -7654 110414 711590
rect 114294 -7654 114914 711590
rect 118794 262000 119414 711590
rect 123294 262000 123914 711590
rect 127794 262000 128414 711590
rect 132294 262000 132914 711590
rect 136794 262000 137414 711590
rect 141294 262000 141914 711590
rect 145794 262000 146414 711590
rect 150294 262000 150914 711590
rect 154794 262000 155414 711590
rect 159294 262000 159914 711590
rect 163794 262000 164414 711590
rect 168294 262000 168914 711590
rect 172794 262000 173414 711590
rect 177294 262000 177914 711590
rect 181794 262000 182414 711590
rect 186294 262000 186914 711590
rect 190794 262000 191414 711590
rect 118794 142000 119414 198000
rect 123294 142000 123914 198000
rect 141294 142000 141914 198000
rect 145794 142000 146414 198000
rect 150294 142000 150914 198000
rect 154794 142000 155414 198000
rect 159294 142000 159914 198000
rect 177294 142000 177914 198000
rect 181794 142000 182414 198000
rect 186294 142000 186914 198000
rect 190794 142000 191414 198000
rect 118794 -7654 119414 78000
rect 123294 -7654 123914 78000
rect 127794 -7654 128414 78000
rect 132294 -7654 132914 78000
rect 136794 -7654 137414 78000
rect 141294 -7654 141914 78000
rect 145794 -7654 146414 78000
rect 150294 -7654 150914 78000
rect 154794 -7654 155414 78000
rect 159294 -7654 159914 78000
rect 163794 -7654 164414 78000
rect 168294 -7654 168914 78000
rect 172794 -7654 173414 78000
rect 177294 -7654 177914 78000
rect 181794 -7654 182414 78000
rect 186294 -7654 186914 78000
rect 190794 -7654 191414 78000
rect 195294 -7654 195914 711590
rect 199794 -7654 200414 711590
rect 204294 -7654 204914 711590
rect 208794 -7654 209414 711590
rect 213294 -7654 213914 711590
rect 217794 -7654 218414 711590
rect 222294 -7654 222914 711590
rect 226794 -7654 227414 711590
rect 231294 -7654 231914 711590
rect 235794 -7654 236414 711590
rect 240294 -7654 240914 711590
rect 244794 -7654 245414 711590
rect 249294 -7654 249914 711590
rect 253794 -7654 254414 711590
rect 258294 -7654 258914 711590
rect 262794 -7654 263414 711590
rect 267294 -7654 267914 711590
rect 271794 -7654 272414 711590
rect 276294 -7654 276914 711590
rect 280794 -7654 281414 711590
rect 285294 -7654 285914 711590
rect 289794 -7654 290414 711590
rect 294294 -7654 294914 711590
rect 298794 -7654 299414 711590
rect 303294 -7654 303914 711590
rect 307794 -7654 308414 711590
rect 312294 -7654 312914 711590
rect 316794 -7654 317414 711590
rect 321294 -7654 321914 711590
rect 325794 -7654 326414 711590
rect 330294 -7654 330914 711590
rect 334794 -7654 335414 711590
rect 339294 -7654 339914 711590
rect 343794 -7654 344414 711590
rect 348294 -7654 348914 711590
rect 352794 -7654 353414 711590
rect 357294 -7654 357914 711590
rect 361794 -7654 362414 711590
rect 366294 -7654 366914 711590
rect 370794 -7654 371414 711590
rect 375294 -7654 375914 711590
rect 379794 -7654 380414 711590
rect 384294 -7654 384914 711590
rect 388794 -7654 389414 711590
rect 393294 -7654 393914 711590
rect 397794 -7654 398414 711590
rect 402294 -7654 402914 711590
rect 406794 -7654 407414 711590
rect 411294 -7654 411914 711590
rect 415794 -7654 416414 711590
rect 420294 -7654 420914 711590
rect 424794 -7654 425414 711590
rect 429294 -7654 429914 711590
rect 433794 -7654 434414 711590
rect 438294 -7654 438914 711590
rect 442794 -7654 443414 711590
rect 447294 -7654 447914 711590
rect 451794 -7654 452414 711590
rect 456294 -7654 456914 711590
rect 460794 -7654 461414 711590
rect 465294 -7654 465914 711590
rect 469794 -7654 470414 711590
rect 474294 -7654 474914 711590
rect 478794 -7654 479414 711590
rect 483294 -7654 483914 711590
rect 487794 -7654 488414 711590
rect 492294 -7654 492914 711590
rect 496794 -7654 497414 711590
rect 501294 -7654 501914 711590
rect 505794 -7654 506414 711590
rect 510294 -7654 510914 711590
rect 514794 -7654 515414 711590
rect 519294 -7654 519914 711590
rect 523794 -7654 524414 711590
rect 528294 -7654 528914 711590
rect 532794 -7654 533414 711590
rect 537294 -7654 537914 711590
rect 541794 -7654 542414 711590
rect 546294 -7654 546914 711590
rect 550794 -7654 551414 711590
rect 555294 -7654 555914 711590
rect 559794 -7654 560414 711590
rect 564294 -7654 564914 711590
rect 568794 -7654 569414 711590
rect 573294 -7654 573914 711590
rect 577794 -7654 578414 711590
rect 582294 -7654 582914 711590
rect 585310 -934 585930 704870
rect 586270 -1894 586890 705830
rect 587230 -2854 587850 706790
rect 588190 -3814 588810 707750
rect 589150 -4774 589770 708710
rect 590110 -5734 590730 709670
rect 591070 -6694 591690 710630
rect 592030 -7654 592650 711590
<< obsm4 >>
rect 99051 62051 100714 269789
rect 101494 62051 105214 269789
rect 105994 62051 109714 269789
rect 110494 62051 114214 269789
rect 114994 261920 118714 269789
rect 119494 261920 123214 269789
rect 123994 261920 127714 269789
rect 128494 261920 132214 269789
rect 132994 261920 136714 269789
rect 137494 261920 141214 269789
rect 141994 261920 145714 269789
rect 146494 261920 150214 269789
rect 150994 261920 154714 269789
rect 155494 261920 159214 269789
rect 159994 261920 163714 269789
rect 164494 261920 168214 269789
rect 168994 261920 172714 269789
rect 173494 261920 177214 269789
rect 177994 261920 181714 269789
rect 182494 261920 186214 269789
rect 186994 261920 190714 269789
rect 191494 261920 195214 269789
rect 114994 198080 195214 261920
rect 114994 141920 118714 198080
rect 119494 141920 123214 198080
rect 123994 141920 141214 198080
rect 141994 141920 145714 198080
rect 146494 141920 150214 198080
rect 150994 141920 154714 198080
rect 155494 141920 159214 198080
rect 159994 141920 177214 198080
rect 177994 141920 181714 198080
rect 182494 141920 186214 198080
rect 186994 141920 190714 198080
rect 191494 141920 195214 198080
rect 114994 78080 195214 141920
rect 114994 62051 118714 78080
rect 119494 62051 123214 78080
rect 123994 62051 127714 78080
rect 128494 62051 132214 78080
rect 132994 62051 136714 78080
rect 137494 62051 141214 78080
rect 141994 62051 145714 78080
rect 146494 62051 150214 78080
rect 150994 62051 154714 78080
rect 155494 62051 159214 78080
rect 159994 62051 163714 78080
rect 164494 62051 168214 78080
rect 168994 62051 172714 78080
rect 173494 62051 177214 78080
rect 177994 62051 181714 78080
rect 182494 62051 186214 78080
rect 186994 62051 190714 78080
rect 191494 62051 195214 78080
rect 195994 62051 199714 269789
rect 200494 62051 204214 269789
rect 204994 62051 208714 269789
rect 209494 62051 213214 269789
rect 213994 62051 214117 269789
<< metal5 >>
rect -8726 710970 592650 711590
rect -7766 710010 591690 710630
rect -6806 709050 590730 709670
rect -5846 708090 589770 708710
rect -4886 707130 588810 707750
rect -3926 706170 587850 706790
rect -2966 705210 586890 705830
rect -2006 704250 585930 704870
rect -8726 700366 592650 700986
rect -8726 695866 592650 696486
rect -8726 691366 592650 691986
rect -8726 686866 592650 687486
rect -8726 682366 592650 682986
rect -8726 677866 592650 678486
rect -8726 673366 592650 673986
rect -8726 668866 592650 669486
rect -8726 664366 592650 664986
rect -8726 659866 592650 660486
rect -8726 655366 592650 655986
rect -8726 650866 592650 651486
rect -8726 646366 592650 646986
rect -8726 641866 592650 642486
rect -8726 637366 592650 637986
rect -8726 632866 592650 633486
rect -8726 628366 592650 628986
rect -8726 623866 592650 624486
rect -8726 619366 592650 619986
rect -8726 614866 592650 615486
rect -8726 610366 592650 610986
rect -8726 605866 592650 606486
rect -8726 601366 592650 601986
rect -8726 596866 592650 597486
rect -8726 592366 592650 592986
rect -8726 587866 592650 588486
rect -8726 583366 592650 583986
rect -8726 578866 592650 579486
rect -8726 574366 592650 574986
rect -8726 569866 592650 570486
rect -8726 565366 592650 565986
rect -8726 560866 592650 561486
rect -8726 556366 592650 556986
rect -8726 551866 592650 552486
rect -8726 547366 592650 547986
rect -8726 542866 592650 543486
rect -8726 538366 592650 538986
rect -8726 533866 592650 534486
rect -8726 529366 592650 529986
rect -8726 524866 592650 525486
rect -8726 520366 592650 520986
rect -8726 515866 592650 516486
rect -8726 511366 592650 511986
rect -8726 506866 592650 507486
rect -8726 502366 592650 502986
rect -8726 497866 592650 498486
rect -8726 493366 592650 493986
rect -8726 488866 592650 489486
rect -8726 484366 592650 484986
rect -8726 479866 592650 480486
rect -8726 475366 592650 475986
rect -8726 470866 592650 471486
rect -8726 466366 592650 466986
rect -8726 461866 592650 462486
rect -8726 457366 592650 457986
rect -8726 452866 592650 453486
rect -8726 448366 592650 448986
rect -8726 443866 592650 444486
rect -8726 439366 592650 439986
rect -8726 434866 592650 435486
rect -8726 430366 592650 430986
rect -8726 425866 592650 426486
rect -8726 421366 592650 421986
rect -8726 416866 592650 417486
rect -8726 412366 592650 412986
rect -8726 407866 592650 408486
rect -8726 403366 592650 403986
rect -8726 398866 592650 399486
rect -8726 394366 592650 394986
rect -8726 389866 592650 390486
rect -8726 385366 592650 385986
rect -8726 380866 592650 381486
rect -8726 376366 592650 376986
rect -8726 371866 592650 372486
rect -8726 367366 592650 367986
rect -8726 362866 592650 363486
rect -8726 358366 592650 358986
rect -8726 353866 592650 354486
rect -8726 349366 592650 349986
rect -8726 344866 592650 345486
rect -8726 340366 592650 340986
rect -8726 335866 592650 336486
rect -8726 331366 592650 331986
rect -8726 326866 592650 327486
rect -8726 322366 592650 322986
rect -8726 317866 592650 318486
rect -8726 313366 592650 313986
rect -8726 308866 592650 309486
rect -8726 304366 592650 304986
rect -8726 299866 592650 300486
rect -8726 295366 592650 295986
rect -8726 290866 592650 291486
rect -8726 286366 592650 286986
rect -8726 281866 592650 282486
rect -8726 277366 592650 277986
rect -8726 272866 592650 273486
rect -8726 268366 592650 268986
rect -8726 263866 592650 264486
rect -8726 259366 592650 259986
rect -8726 254866 592650 255486
rect -8726 250366 592650 250986
rect -8726 245866 592650 246486
rect -8726 241366 592650 241986
rect -8726 236866 592650 237486
rect -8726 232366 592650 232986
rect -8726 227866 592650 228486
rect -8726 223366 592650 223986
rect -8726 218866 592650 219486
rect -8726 214366 592650 214986
rect -8726 209866 592650 210486
rect -8726 205366 592650 205986
rect -8726 200866 592650 201486
rect -8726 196366 592650 196986
rect -8726 191866 592650 192486
rect -8726 187366 592650 187986
rect -8726 182866 592650 183486
rect -8726 178366 592650 178986
rect -8726 173866 592650 174486
rect -8726 169366 592650 169986
rect -8726 164866 592650 165486
rect -8726 160366 592650 160986
rect -8726 155866 592650 156486
rect -8726 151366 592650 151986
rect -8726 146866 592650 147486
rect -8726 142366 592650 142986
rect -8726 137866 592650 138486
rect -8726 133366 592650 133986
rect -8726 128866 592650 129486
rect -8726 124366 592650 124986
rect -8726 119866 592650 120486
rect -8726 115366 592650 115986
rect -8726 110866 592650 111486
rect -8726 106366 592650 106986
rect -8726 101866 592650 102486
rect -8726 97366 592650 97986
rect -8726 92866 592650 93486
rect -8726 88366 592650 88986
rect -8726 83866 592650 84486
rect -8726 79366 592650 79986
rect -8726 74866 592650 75486
rect -8726 70366 592650 70986
rect -8726 65866 592650 66486
rect -8726 61366 592650 61986
rect -8726 56866 592650 57486
rect -8726 52366 592650 52986
rect -8726 47866 592650 48486
rect -8726 43366 592650 43986
rect -8726 38866 592650 39486
rect -8726 34366 592650 34986
rect -8726 29866 592650 30486
rect -8726 25366 592650 25986
rect -8726 20866 592650 21486
rect -8726 16366 592650 16986
rect -8726 11866 592650 12486
rect -8726 7366 592650 7986
rect -8726 2866 592650 3486
rect -2006 -934 585930 -314
rect -2966 -1894 586890 -1274
rect -3926 -2854 587850 -2234
rect -4886 -3814 588810 -3194
rect -5846 -4774 589770 -4154
rect -6806 -5734 590730 -5114
rect -7766 -6694 591690 -6074
rect -8726 -7654 592650 -7034
<< labels >>
rlabel metal2 s 87574 -960 87686 480 8 gpio_analog[0]
port 1 nsew signal bidirectional
rlabel metal2 s 156482 -960 156594 480 8 gpio_analog[10]
port 2 nsew signal bidirectional
rlabel metal3 s 583520 56388 584960 56628 6 gpio_analog[11]
port 3 nsew signal bidirectional
rlabel metal2 s 100454 703520 100566 704960 6 gpio_analog[12]
port 4 nsew signal bidirectional
rlabel metal3 s -960 326348 480 326588 4 gpio_analog[13]
port 5 nsew signal bidirectional
rlabel metal2 s 345174 703520 345286 704960 6 gpio_analog[14]
port 6 nsew signal bidirectional
rlabel metal3 s 583520 222308 584960 222548 6 gpio_analog[15]
port 7 nsew signal bidirectional
rlabel metal3 s -960 637108 480 637348 4 gpio_analog[16]
port 8 nsew signal bidirectional
rlabel metal3 s -960 128468 480 128708 4 gpio_analog[17]
port 9 nsew signal bidirectional
rlabel metal3 s 583520 80868 584960 81108 6 gpio_analog[1]
port 10 nsew signal bidirectional
rlabel metal2 s 259522 -960 259634 480 8 gpio_analog[2]
port 11 nsew signal bidirectional
rlabel metal3 s -960 435148 480 435388 4 gpio_analog[3]
port 12 nsew signal bidirectional
rlabel metal3 s 583520 673828 584960 674068 6 gpio_analog[4]
port 13 nsew signal bidirectional
rlabel metal3 s -960 205308 480 205548 4 gpio_analog[5]
port 14 nsew signal bidirectional
rlabel metal3 s -960 399108 480 399348 4 gpio_analog[6]
port 15 nsew signal bidirectional
rlabel metal2 s 75982 -960 76094 480 8 gpio_analog[7]
port 16 nsew signal bidirectional
rlabel metal2 s 546102 -960 546214 480 8 gpio_analog[8]
port 17 nsew signal bidirectional
rlabel metal2 s 412150 -960 412262 480 8 gpio_analog[9]
port 18 nsew signal bidirectional
rlabel metal2 s 240202 -960 240314 480 8 gpio_noesd[0]
port 19 nsew signal bidirectional
rlabel metal3 s -960 536468 480 536708 4 gpio_noesd[10]
port 20 nsew signal bidirectional
rlabel metal3 s -960 447388 480 447628 4 gpio_noesd[11]
port 21 nsew signal bidirectional
rlabel metal2 s 173226 703520 173338 704960 6 gpio_noesd[12]
port 22 nsew signal bidirectional
rlabel metal2 s 390898 703520 391010 704960 6 gpio_noesd[13]
port 23 nsew signal bidirectional
rlabel metal3 s -960 382788 480 383028 4 gpio_noesd[14]
port 24 nsew signal bidirectional
rlabel metal3 s -960 59788 480 60028 4 gpio_noesd[15]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 28508 584960 28748 6 gpio_noesd[16]
port 26 nsew signal bidirectional
rlabel metal2 s 211222 703520 211334 704960 6 gpio_noesd[17]
port 27 nsew signal bidirectional
rlabel metal2 s 121706 -960 121818 480 8 gpio_noesd[1]
port 28 nsew signal bidirectional
rlabel metal2 s 328430 -960 328542 480 8 gpio_noesd[2]
port 29 nsew signal bidirectional
rlabel metal3 s 583520 641868 584960 642108 6 gpio_noesd[3]
port 30 nsew signal bidirectional
rlabel metal2 s 191902 703520 192014 704960 6 gpio_noesd[4]
port 31 nsew signal bidirectional
rlabel metal3 s 583520 64548 584960 64788 6 gpio_noesd[5]
port 32 nsew signal bidirectional
rlabel metal3 s 583520 601068 584960 601308 6 gpio_noesd[6]
port 33 nsew signal bidirectional
rlabel metal3 s 583520 492268 584960 492508 6 gpio_noesd[7]
port 34 nsew signal bidirectional
rlabel metal3 s -960 88348 480 88588 4 gpio_noesd[8]
port 35 nsew signal bidirectional
rlabel metal3 s -960 132548 480 132788 4 gpio_noesd[9]
port 36 nsew signal bidirectional
rlabel metal3 s -960 245428 480 245668 4 io_analog[0]
port 37 nsew signal bidirectional
rlabel metal2 s 56662 -960 56774 480 8 io_analog[10]
port 38 nsew signal bidirectional
rlabel metal3 s 583520 60468 584960 60708 6 io_analog[1]
port 39 nsew signal bidirectional
rlabel metal3 s 583520 552788 584960 553028 6 io_analog[2]
port 40 nsew signal bidirectional
rlabel metal2 s 228610 -960 228722 480 8 io_analog[3]
port 41 nsew signal bidirectional
rlabel metal2 s 113978 -960 114090 480 8 io_analog[4]
port 42 nsew signal bidirectional
rlabel metal2 s 88862 703520 88974 704960 6 io_analog[5]
port 43 nsew signal bidirectional
rlabel metal2 s 450790 -960 450902 480 8 io_analog[6]
port 44 nsew signal bidirectional
rlabel metal3 s -960 233868 480 234108 4 io_analog[7]
port 45 nsew signal bidirectional
rlabel metal2 s 209934 -960 210046 480 8 io_analog[8]
port 46 nsew signal bidirectional
rlabel metal3 s -960 334508 480 334748 4 io_analog[9]
port 47 nsew signal bidirectional
rlabel metal2 s 22530 -960 22642 480 8 io_clamp_high[0]
port 48 nsew signal bidirectional
rlabel metal3 s 583520 581348 584960 581588 6 io_clamp_high[1]
port 49 nsew signal bidirectional
rlabel metal3 s 583520 363068 584960 363308 6 io_clamp_high[2]
port 50 nsew signal bidirectional
rlabel metal3 s -960 124388 480 124628 4 io_clamp_low[0]
port 51 nsew signal bidirectional
rlabel metal2 s 285926 -960 286038 480 8 io_clamp_low[1]
port 52 nsew signal bidirectional
rlabel metal3 s -960 649348 480 649588 4 io_clamp_low[2]
port 53 nsew signal bidirectional
rlabel metal2 s 37986 -960 38098 480 8 io_in[0]
port 54 nsew signal input
rlabel metal3 s 583520 504508 584960 504748 6 io_in[10]
port 55 nsew signal input
rlabel metal2 s 493938 703520 494050 704960 6 io_in[11]
port 56 nsew signal input
rlabel metal2 s 402490 703520 402602 704960 6 io_in[12]
port 57 nsew signal input
rlabel metal2 s 99166 -960 99278 480 8 io_in[13]
port 58 nsew signal input
rlabel metal2 s 416014 -960 416126 480 8 io_in[14]
port 59 nsew signal input
rlabel metal3 s -960 76108 480 76348 4 io_in[15]
port 60 nsew signal input
rlabel metal2 s 519054 -960 519166 480 8 io_in[16]
port 61 nsew signal input
rlabel metal3 s 583520 237948 584960 238188 6 io_in[17]
port 62 nsew signal input
rlabel metal3 s 583520 72708 584960 72948 6 io_in[18]
port 63 nsew signal input
rlabel metal3 s -960 564348 480 564588 4 io_in[19]
port 64 nsew signal input
rlabel metal2 s 492650 -960 492762 480 8 io_in[1]
port 65 nsew signal input
rlabel metal2 s 534510 -960 534622 480 8 io_in[20]
port 66 nsew signal input
rlabel metal2 s 336158 -960 336270 480 8 io_in[21]
port 67 nsew signal input
rlabel metal3 s 583520 133228 584960 133468 6 io_in[22]
port 68 nsew signal input
rlabel metal2 s 264674 703520 264786 704960 6 io_in[23]
port 69 nsew signal input
rlabel metal3 s 583520 399788 584960 400028 6 io_in[24]
port 70 nsew signal input
rlabel metal2 s 580234 -960 580346 480 8 io_in[25]
port 71 nsew signal input
rlabel metal2 s 535798 703520 535910 704960 6 io_in[26]
port 72 nsew signal input
rlabel metal3 s 583520 452148 584960 452388 6 io_in[2]
port 73 nsew signal input
rlabel metal3 s -960 314108 480 314348 4 io_in[3]
port 74 nsew signal input
rlabel metal2 s 427606 -960 427718 480 8 io_in[4]
port 75 nsew signal input
rlabel metal2 s 130722 703520 130834 704960 6 io_in[5]
port 76 nsew signal input
rlabel metal3 s 583520 548708 584960 548948 6 io_in[6]
port 77 nsew signal input
rlabel metal3 s -960 56388 480 56628 4 io_in[7]
port 78 nsew signal input
rlabel metal2 s 83710 -960 83822 480 8 io_in[8]
port 79 nsew signal input
rlabel metal2 s 230542 703520 230654 704960 6 io_in[9]
port 80 nsew signal input
rlabel metal2 s 164210 -960 164322 480 8 io_in_3v3[0]
port 81 nsew signal input
rlabel metal2 s 45714 -960 45826 480 8 io_in_3v3[10]
port 82 nsew signal input
rlabel metal2 s 337446 703520 337558 704960 6 io_in_3v3[11]
port 83 nsew signal input
rlabel metal2 s 531934 703520 532046 704960 6 io_in_3v3[12]
port 84 nsew signal input
rlabel metal2 s 10938 -960 11050 480 8 io_in_3v3[13]
port 85 nsew signal input
rlabel metal3 s -960 641188 480 641428 4 io_in_3v3[14]
port 86 nsew signal input
rlabel metal3 s 583520 205988 584960 206228 6 io_in_3v3[15]
port 87 nsew signal input
rlabel metal3 s 583520 157708 584960 157948 6 io_in_3v3[16]
port 88 nsew signal input
rlabel metal3 s -960 657508 480 657748 4 io_in_3v3[17]
port 89 nsew signal input
rlabel metal3 s -960 366468 480 366708 4 io_in_3v3[18]
port 90 nsew signal input
rlabel metal3 s -960 633028 480 633268 4 io_in_3v3[19]
port 91 nsew signal input
rlabel metal3 s 583520 52308 584960 52548 6 io_in_3v3[1]
port 92 nsew signal input
rlabel metal2 s 73406 703520 73518 704960 6 io_in_3v3[20]
port 93 nsew signal input
rlabel metal3 s -960 592908 480 593148 4 io_in_3v3[21]
port 94 nsew signal input
rlabel metal3 s -960 697628 480 697868 4 io_in_3v3[22]
port 95 nsew signal input
rlabel metal3 s -960 677228 480 677468 4 io_in_3v3[23]
port 96 nsew signal input
rlabel metal2 s 293654 -960 293766 480 8 io_in_3v3[24]
port 97 nsew signal input
rlabel metal3 s 583520 335188 584960 335428 6 io_in_3v3[25]
port 98 nsew signal input
rlabel metal3 s -960 395028 480 395268 4 io_in_3v3[26]
port 99 nsew signal input
rlabel metal2 s 1278 703520 1390 704960 6 io_in_3v3[2]
port 100 nsew signal input
rlabel metal3 s 583520 653428 584960 653668 6 io_in_3v3[3]
port 101 nsew signal input
rlabel metal2 s 566710 703520 566822 704960 6 io_in_3v3[4]
port 102 nsew signal input
rlabel metal2 s 312974 -960 313086 480 8 io_in_3v3[5]
port 103 nsew signal input
rlabel metal2 s 446926 -960 447038 480 8 io_in_3v3[6]
port 104 nsew signal input
rlabel metal2 s 198342 -960 198454 480 8 io_in_3v3[7]
port 105 nsew signal input
rlabel metal2 s 295586 703520 295698 704960 6 io_in_3v3[8]
port 106 nsew signal input
rlabel metal2 s 553830 -960 553942 480 8 io_in_3v3[9]
port 107 nsew signal input
rlabel metal3 s -960 475948 480 476188 4 io_oeb[0]
port 108 nsew signal output
rlabel metal2 s 474618 703520 474730 704960 6 io_oeb[10]
port 109 nsew signal output
rlabel metal2 s 218950 703520 219062 704960 6 io_oeb[11]
port 110 nsew signal output
rlabel metal2 s 366426 -960 366538 480 8 io_oeb[12]
port 111 nsew signal output
rlabel metal2 s 515190 -960 515302 480 8 io_oeb[13]
port 112 nsew signal output
rlabel metal3 s 583520 350828 584960 351068 6 io_oeb[14]
port 113 nsew signal output
rlabel metal3 s -960 487508 480 487748 4 io_oeb[15]
port 114 nsew signal output
rlabel metal3 s -960 528308 480 528548 4 io_oeb[16]
port 115 nsew signal output
rlabel metal3 s 583520 592908 584960 593148 6 io_oeb[17]
port 116 nsew signal output
rlabel metal2 s 129434 -960 129546 480 8 io_oeb[18]
port 117 nsew signal output
rlabel metal3 s 583520 649348 584960 649588 6 io_oeb[19]
port 118 nsew signal output
rlabel metal2 s 501666 703520 501778 704960 6 io_oeb[1]
port 119 nsew signal output
rlabel metal2 s 524850 703520 524962 704960 6 io_oeb[20]
port 120 nsew signal output
rlabel metal2 s 478482 703520 478594 704960 6 io_oeb[21]
port 121 nsew signal output
rlabel metal2 s 60526 -960 60638 480 8 io_oeb[22]
port 122 nsew signal output
rlabel metal3 s 583520 169268 584960 169508 6 io_oeb[23]
port 123 nsew signal output
rlabel metal2 s 349038 703520 349150 704960 6 io_oeb[24]
port 124 nsew signal output
rlabel metal3 s 583520 484108 584960 484348 6 io_oeb[25]
port 125 nsew signal output
rlabel metal3 s 583520 375308 584960 375548 6 io_oeb[26]
port 126 nsew signal output
rlabel metal3 s -960 608548 480 608788 4 io_oeb[2]
port 127 nsew signal output
rlabel metal3 s -960 624868 480 625108 4 io_oeb[3]
port 128 nsew signal output
rlabel metal3 s -960 467788 480 468028 4 io_oeb[4]
port 129 nsew signal output
rlabel metal3 s 583520 560948 584960 561188 6 io_oeb[5]
port 130 nsew signal output
rlabel metal2 s 39274 703520 39386 704960 6 io_oeb[6]
port 131 nsew signal output
rlabel metal3 s -960 520148 480 520388 4 io_oeb[7]
port 132 nsew signal output
rlabel metal2 s 299450 703520 299562 704960 6 io_oeb[8]
port 133 nsew signal output
rlabel metal3 s 583520 294388 584960 294628 6 io_oeb[9]
port 134 nsew signal output
rlabel metal2 s 520986 703520 521098 704960 6 io_out[0]
port 135 nsew signal output
rlabel metal3 s -960 177428 480 177668 4 io_out[10]
port 136 nsew signal output
rlabel metal3 s 583520 665668 584960 665908 6 io_out[11]
port 137 nsew signal output
rlabel metal3 s -960 298468 480 298708 4 io_out[12]
port 138 nsew signal output
rlabel metal3 s 583520 415428 584960 415668 6 io_out[13]
port 139 nsew signal output
rlabel metal2 s 268538 703520 268650 704960 6 io_out[14]
port 140 nsew signal output
rlabel metal3 s -960 346748 480 346988 4 io_out[15]
port 141 nsew signal output
rlabel metal2 s 58594 703520 58706 704960 6 io_out[16]
port 142 nsew signal output
rlabel metal2 s 195766 703520 195878 704960 6 io_out[17]
port 143 nsew signal output
rlabel metal2 s 23818 703520 23930 704960 6 io_out[18]
port 144 nsew signal output
rlabel metal3 s 583520 266508 584960 266748 6 io_out[19]
port 145 nsew signal output
rlabel metal3 s 583520 407268 584960 407508 6 io_out[1]
port 146 nsew signal output
rlabel metal2 s 70186 703520 70298 704960 6 io_out[20]
port 147 nsew signal output
rlabel metal2 s 271114 -960 271226 480 8 io_out[21]
port 148 nsew signal output
rlabel metal3 s -960 184908 480 185148 4 io_out[22]
port 149 nsew signal output
rlabel metal3 s 583520 354908 584960 355148 6 io_out[23]
port 150 nsew signal output
rlabel metal3 s -960 685388 480 685628 4 io_out[24]
port 151 nsew signal output
rlabel metal3 s -960 269908 480 270148 4 io_out[25]
port 152 nsew signal output
rlabel metal2 s 221526 -960 221638 480 8 io_out[26]
port 153 nsew signal output
rlabel metal2 s 179022 -960 179134 480 8 io_out[2]
port 154 nsew signal output
rlabel metal2 s 276266 703520 276378 704960 6 io_out[3]
port 155 nsew signal output
rlabel metal2 s 470754 703520 470866 704960 6 io_out[4]
port 156 nsew signal output
rlabel metal3 s -960 483428 480 483668 4 io_out[5]
port 157 nsew signal output
rlabel metal3 s 583520 165188 584960 165428 6 io_out[6]
port 158 nsew signal output
rlabel metal3 s -960 653428 480 653668 4 io_out[7]
port 159 nsew signal output
rlabel metal3 s 583520 120988 584960 121228 6 io_out[8]
port 160 nsew signal output
rlabel metal3 s 583520 250188 584960 250428 6 io_out[9]
port 161 nsew signal output
rlabel metal2 s 157770 703520 157882 704960 6 la_data_in[0]
port 162 nsew signal input
rlabel metal3 s 583520 625548 584960 625788 6 la_data_in[100]
port 163 nsew signal input
rlabel metal3 s 583520 214148 584960 214388 6 la_data_in[101]
port 164 nsew signal input
rlabel metal2 s 387034 703520 387146 704960 6 la_data_in[102]
port 165 nsew signal input
rlabel metal3 s 583520 20348 584960 20588 6 la_data_in[103]
port 166 nsew signal input
rlabel metal3 s -960 370548 480 370788 4 la_data_in[104]
port 167 nsew signal input
rlabel metal2 s 222814 703520 222926 704960 6 la_data_in[105]
port 168 nsew signal input
rlabel metal2 s 134586 703520 134698 704960 6 la_data_in[106]
port 169 nsew signal input
rlabel metal3 s -960 415428 480 415668 4 la_data_in[107]
port 170 nsew signal input
rlabel metal3 s 583520 584748 584960 584988 6 la_data_in[108]
port 171 nsew signal input
rlabel metal3 s -960 161108 480 161348 4 la_data_in[109]
port 172 nsew signal input
rlabel metal3 s 583520 379388 584960 379628 6 la_data_in[10]
port 173 nsew signal input
rlabel metal3 s -960 286228 480 286468 4 la_data_in[110]
port 174 nsew signal input
rlabel metal3 s 583520 270588 584960 270828 6 la_data_in[111]
port 175 nsew signal input
rlabel metal3 s -960 374628 480 374868 4 la_data_in[112]
port 176 nsew signal input
rlabel metal3 s -960 673148 480 673388 4 la_data_in[113]
port 177 nsew signal input
rlabel metal3 s -960 516068 480 516308 4 la_data_in[114]
port 178 nsew signal input
rlabel metal2 s 325854 703520 325966 704960 6 la_data_in[115]
port 179 nsew signal input
rlabel metal2 s 526782 -960 526894 480 8 la_data_in[116]
port 180 nsew signal input
rlabel metal3 s -960 338588 480 338828 4 la_data_in[117]
port 181 nsew signal input
rlabel metal3 s 583520 520828 584960 521068 6 la_data_in[118]
port 182 nsew signal input
rlabel metal3 s 583520 210068 584960 210308 6 la_data_in[119]
port 183 nsew signal input
rlabel metal2 s 96590 703520 96702 704960 6 la_data_in[11]
port 184 nsew signal input
rlabel metal3 s -960 305948 480 306188 4 la_data_in[120]
port 185 nsew signal input
rlabel metal2 s 160346 -960 160458 480 8 la_data_in[121]
port 186 nsew signal input
rlabel metal2 s 137162 -960 137274 480 8 la_data_in[122]
port 187 nsew signal input
rlabel metal3 s -960 426988 480 427228 4 la_data_in[123]
port 188 nsew signal input
rlabel metal2 s 413438 703520 413550 704960 6 la_data_in[124]
port 189 nsew signal input
rlabel metal2 s 484922 -960 485034 480 8 la_data_in[125]
port 190 nsew signal input
rlabel metal3 s -960 419508 480 419748 4 la_data_in[126]
port 191 nsew signal input
rlabel metal2 s 558982 703520 559094 704960 6 la_data_in[127]
port 192 nsew signal input
rlabel metal3 s 583520 185588 584960 185828 6 la_data_in[12]
port 193 nsew signal input
rlabel metal3 s 583520 339268 584960 339508 6 la_data_in[13]
port 194 nsew signal input
rlabel metal3 s -960 539868 480 540108 4 la_data_in[14]
port 195 nsew signal input
rlabel metal3 s -960 548028 480 548268 4 la_data_in[15]
port 196 nsew signal input
rlabel metal3 s -960 67948 480 68188 4 la_data_in[16]
port 197 nsew signal input
rlabel metal3 s -960 157028 480 157268 4 la_data_in[17]
port 198 nsew signal input
rlabel metal3 s -960 451468 480 451708 4 la_data_in[18]
port 199 nsew signal input
rlabel metal2 s 448214 703520 448326 704960 6 la_data_in[19]
port 200 nsew signal input
rlabel metal2 s 301382 -960 301494 480 8 la_data_in[1]
port 201 nsew signal input
rlabel metal3 s -960 310028 480 310268 4 la_data_in[20]
port 202 nsew signal input
rlabel metal2 s 27682 703520 27794 704960 6 la_data_in[21]
port 203 nsew signal input
rlabel metal2 s 180954 703520 181066 704960 6 la_data_in[22]
port 204 nsew signal input
rlabel metal3 s -960 439228 480 439468 4 la_data_in[23]
port 205 nsew signal input
rlabel metal3 s 583520 423588 584960 423828 6 la_data_in[24]
port 206 nsew signal input
rlabel metal2 s 432758 703520 432870 704960 6 la_data_in[25]
port 207 nsew signal input
rlabel metal2 s 504242 -960 504354 480 8 la_data_in[26]
port 208 nsew signal input
rlabel metal2 s 289790 -960 289902 480 8 la_data_in[27]
port 209 nsew signal input
rlabel metal3 s -960 463708 480 463948 4 la_data_in[28]
port 210 nsew signal input
rlabel metal3 s -960 342668 480 342908 4 la_data_in[29]
port 211 nsew signal input
rlabel metal2 s 439198 -960 439310 480 8 la_data_in[2]
port 212 nsew signal input
rlabel metal3 s -960 491588 480 491828 4 la_data_in[30]
port 213 nsew signal input
rlabel metal3 s 583520 605148 584960 605388 6 la_data_in[31]
port 214 nsew signal input
rlabel metal2 s 302670 703520 302782 704960 6 la_data_in[32]
port 215 nsew signal input
rlabel metal3 s 583520 588828 584960 589068 6 la_data_in[33]
port 216 nsew signal input
rlabel metal3 s -960 7428 480 7668 4 la_data_in[34]
port 217 nsew signal input
rlabel metal3 s -960 664988 480 665228 4 la_data_in[35]
port 218 nsew signal input
rlabel metal2 s 551254 703520 551366 704960 6 la_data_in[36]
port 219 nsew signal input
rlabel metal2 s 543526 703520 543638 704960 6 la_data_in[37]
port 220 nsew signal input
rlabel metal2 s 329718 703520 329830 704960 6 la_data_in[38]
port 221 nsew signal input
rlabel metal2 s 148754 -960 148866 480 8 la_data_in[39]
port 222 nsew signal input
rlabel metal3 s 583520 395708 584960 395948 6 la_data_in[3]
port 223 nsew signal input
rlabel metal2 s 138450 703520 138562 704960 6 la_data_in[40]
port 224 nsew signal input
rlabel metal3 s -960 620788 480 621028 4 la_data_in[41]
port 225 nsew signal input
rlabel metal3 s -960 144788 480 145028 4 la_data_in[42]
port 226 nsew signal input
rlabel metal3 s 583520 318868 584960 319108 6 la_data_in[43]
port 227 nsew signal input
rlabel metal3 s -960 459628 480 459868 4 la_data_in[44]
port 228 nsew signal input
rlabel metal2 s 81134 703520 81246 704960 6 la_data_in[45]
port 229 nsew signal input
rlabel metal2 s 123638 703520 123750 704960 6 la_data_in[46]
port 230 nsew signal input
rlabel metal3 s -960 580668 480 580908 4 la_data_in[47]
port 231 nsew signal input
rlabel metal3 s 583520 419508 584960 419748 6 la_data_in[48]
port 232 nsew signal input
rlabel metal3 s 583520 32588 584960 32828 6 la_data_in[49]
port 233 nsew signal input
rlabel metal2 s 431470 -960 431582 480 8 la_data_in[4]
port 234 nsew signal input
rlabel metal2 s 488786 -960 488898 480 8 la_data_in[50]
port 235 nsew signal input
rlabel metal3 s 583520 500428 584960 500668 6 la_data_in[51]
port 236 nsew signal input
rlabel metal3 s -960 552108 480 552348 4 la_data_in[52]
port 237 nsew signal input
rlabel metal2 s 255658 -960 255770 480 8 la_data_in[53]
port 238 nsew signal input
rlabel metal2 s 3210 -960 3322 480 8 la_data_in[54]
port 239 nsew signal input
rlabel metal3 s 583520 322948 584960 323188 6 la_data_in[55]
port 240 nsew signal input
rlabel metal3 s -960 507908 480 508148 4 la_data_in[56]
port 241 nsew signal input
rlabel metal3 s 583520 411348 584960 411588 6 la_data_in[57]
port 242 nsew signal input
rlabel metal2 s 394762 703520 394874 704960 6 la_data_in[58]
port 243 nsew signal input
rlabel metal3 s -960 104668 480 104908 4 la_data_in[59]
port 244 nsew signal input
rlabel metal3 s -960 612628 480 612868 4 la_data_in[5]
port 245 nsew signal input
rlabel metal2 s 542238 -960 542350 480 8 la_data_in[60]
port 246 nsew signal input
rlabel metal2 s 568642 -960 568754 480 8 la_data_in[61]
port 247 nsew signal input
rlabel metal3 s 583520 48228 584960 48468 6 la_data_in[62]
port 248 nsew signal input
rlabel metal3 s -960 188988 480 189228 4 la_data_in[63]
port 249 nsew signal input
rlabel metal3 s 583520 173348 584960 173588 6 la_data_in[64]
port 250 nsew signal input
rlabel metal3 s 583520 577268 584960 577508 6 la_data_in[65]
port 251 nsew signal input
rlabel metal3 s 583520 331108 584960 331348 6 la_data_in[66]
port 252 nsew signal input
rlabel metal2 s 79846 -960 79958 480 8 la_data_in[67]
port 253 nsew signal input
rlabel metal3 s 583520 565028 584960 565268 6 la_data_in[68]
port 254 nsew signal input
rlabel metal3 s 583520 677908 584960 678148 6 la_data_in[69]
port 255 nsew signal input
rlabel metal3 s 583520 298468 584960 298708 6 la_data_in[6]
port 256 nsew signal input
rlabel metal3 s -960 499748 480 499988 4 la_data_in[70]
port 257 nsew signal input
rlabel metal3 s -960 165188 480 165428 4 la_data_in[71]
port 258 nsew signal input
rlabel metal2 s 62458 703520 62570 704960 6 la_data_in[72]
port 259 nsew signal input
rlabel metal3 s -960 100588 480 100828 4 la_data_in[73]
port 260 nsew signal input
rlabel metal3 s 583520 327028 584960 327268 6 la_data_in[74]
port 261 nsew signal input
rlabel metal2 s 127502 703520 127614 704960 6 la_data_in[75]
port 262 nsew signal input
rlabel metal3 s 583520 149548 584960 149788 6 la_data_in[76]
port 263 nsew signal input
rlabel metal2 s 165498 703520 165610 704960 6 la_data_in[77]
port 264 nsew signal input
rlabel metal2 s 238270 703520 238382 704960 6 la_data_in[78]
port 265 nsew signal input
rlabel metal3 s 583520 536468 584960 536708 6 la_data_in[79]
port 266 nsew signal input
rlabel metal2 s 343242 -960 343354 480 8 la_data_in[7]
port 267 nsew signal input
rlabel metal3 s -960 330428 480 330668 4 la_data_in[80]
port 268 nsew signal input
rlabel metal2 s 505530 703520 505642 704960 6 la_data_in[81]
port 269 nsew signal input
rlabel metal2 s 150042 703520 150154 704960 6 la_data_in[82]
port 270 nsew signal input
rlabel metal3 s 583520 661588 584960 661828 6 la_data_in[83]
port 271 nsew signal input
rlabel metal3 s -960 681308 480 681548 4 la_data_in[84]
port 272 nsew signal input
rlabel metal3 s 583520 367148 584960 367388 6 la_data_in[85]
port 273 nsew signal input
rlabel metal3 s 583520 448068 584960 448308 6 la_data_in[86]
port 274 nsew signal input
rlabel metal2 s 95302 -960 95414 480 8 la_data_in[87]
port 275 nsew signal input
rlabel metal3 s 583520 488188 584960 488428 6 la_data_in[88]
port 276 nsew signal input
rlabel metal2 s 251794 -960 251906 480 8 la_data_in[89]
port 277 nsew signal input
rlabel metal2 s 274978 -960 275090 480 8 la_data_in[8]
port 278 nsew signal input
rlabel metal3 s -960 604468 480 604708 4 la_data_in[90]
port 279 nsew signal input
rlabel metal3 s -960 532388 480 532628 4 la_data_in[91]
port 280 nsew signal input
rlabel metal3 s 583520 12188 584960 12428 6 la_data_in[92]
port 281 nsew signal input
rlabel metal3 s -960 197148 480 197388 4 la_data_in[93]
port 282 nsew signal input
rlabel metal3 s 583520 314788 584960 315028 6 la_data_in[94]
port 283 nsew signal input
rlabel metal3 s -960 96508 480 96748 4 la_data_in[95]
port 284 nsew signal input
rlabel metal3 s -960 511988 480 512228 4 la_data_in[96]
port 285 nsew signal input
rlabel metal3 s -960 568428 480 568668 4 la_data_in[97]
port 286 nsew signal input
rlabel metal2 s 282706 -960 282818 480 8 la_data_in[98]
port 287 nsew signal input
rlabel metal3 s 583520 573188 584960 573428 6 la_data_in[99]
port 288 nsew signal input
rlabel metal2 s 119774 703520 119886 704960 6 la_data_in[9]
port 289 nsew signal input
rlabel metal3 s -960 503828 480 504068 4 la_data_out[0]
port 290 nsew signal output
rlabel metal2 s 253082 703520 253194 704960 6 la_data_out[100]
port 291 nsew signal output
rlabel metal2 s 232474 -960 232586 480 8 la_data_out[101]
port 292 nsew signal output
rlabel metal2 s 169362 703520 169474 704960 6 la_data_out[102]
port 293 nsew signal output
rlabel metal3 s 583520 254268 584960 254508 6 la_data_out[103]
port 294 nsew signal output
rlabel metal2 s 161634 703520 161746 704960 6 la_data_out[104]
port 295 nsew signal output
rlabel metal3 s 583520 189668 584960 189908 6 la_data_out[105]
port 296 nsew signal output
rlabel metal2 s 152618 -960 152730 480 8 la_data_out[106]
port 297 nsew signal output
rlabel metal3 s 583520 387548 584960 387788 6 la_data_out[107]
port 298 nsew signal output
rlabel metal3 s 583520 512668 584960 512908 6 la_data_out[108]
port 299 nsew signal output
rlabel metal2 s 509394 703520 509506 704960 6 la_data_out[109]
port 300 nsew signal output
rlabel metal3 s -960 386868 480 387108 4 la_data_out[10]
port 301 nsew signal output
rlabel metal3 s -960 213468 480 213708 4 la_data_out[110]
port 302 nsew signal output
rlabel metal3 s -960 282148 480 282388 4 la_data_out[111]
port 303 nsew signal output
rlabel metal3 s -960 701708 480 701948 4 la_data_out[112]
port 304 nsew signal output
rlabel metal2 s 202206 -960 202318 480 8 la_data_out[113]
port 305 nsew signal output
rlabel metal2 s 570574 703520 570686 704960 6 la_data_out[114]
port 306 nsew signal output
rlabel metal2 s 375442 703520 375554 704960 6 la_data_out[115]
port 307 nsew signal output
rlabel metal2 s 408286 -960 408398 480 8 la_data_out[116]
port 308 nsew signal output
rlabel metal3 s 583520 645268 584960 645508 6 la_data_out[117]
port 309 nsew signal output
rlabel metal3 s 583520 391628 584960 391868 6 la_data_out[118]
port 310 nsew signal output
rlabel metal3 s 583520 24428 584960 24668 6 la_data_out[119]
port 311 nsew signal output
rlabel metal2 s 452078 703520 452190 704960 6 la_data_out[11]
port 312 nsew signal output
rlabel metal2 s 18666 -960 18778 480 8 la_data_out[120]
port 313 nsew signal output
rlabel metal2 s 184818 703520 184930 704960 6 la_data_out[121]
port 314 nsew signal output
rlabel metal2 s 379306 703520 379418 704960 6 la_data_out[122]
port 315 nsew signal output
rlabel metal3 s -960 229788 480 230028 4 la_data_out[123]
port 316 nsew signal output
rlabel metal3 s 583520 137308 584960 137548 6 la_data_out[124]
port 317 nsew signal output
rlabel metal3 s 583520 480028 584960 480268 6 la_data_out[125]
port 318 nsew signal output
rlabel metal3 s -960 31908 480 32148 4 la_data_out[126]
port 319 nsew signal output
rlabel metal3 s -960 354908 480 355148 4 la_data_out[127]
port 320 nsew signal output
rlabel metal2 s 225390 -960 225502 480 8 la_data_out[12]
port 321 nsew signal output
rlabel metal3 s 583520 40748 584960 40988 6 la_data_out[13]
port 322 nsew signal output
rlabel metal3 s -960 362388 480 362628 4 la_data_out[14]
port 323 nsew signal output
rlabel metal3 s -960 455548 480 455788 4 la_data_out[15]
port 324 nsew signal output
rlabel metal2 s 341310 703520 341422 704960 6 la_data_out[16]
port 325 nsew signal output
rlabel metal3 s 583520 431748 584960 431988 6 la_data_out[17]
port 326 nsew signal output
rlabel metal2 s 110758 -960 110870 480 8 la_data_out[18]
port 327 nsew signal output
rlabel metal2 s 188038 703520 188150 704960 6 la_data_out[19]
port 328 nsew signal output
rlabel metal3 s 583520 93108 584960 93348 6 la_data_out[1]
port 329 nsew signal output
rlabel metal3 s -960 27828 480 28068 4 la_data_out[20]
port 330 nsew signal output
rlabel metal3 s 583520 225708 584960 225948 6 la_data_out[21]
port 331 nsew signal output
rlabel metal3 s 583520 698308 584960 698548 6 la_data_out[22]
port 332 nsew signal output
rlabel metal3 s 583520 229788 584960 230028 6 la_data_out[23]
port 333 nsew signal output
rlabel metal3 s -960 689468 480 689708 4 la_data_out[24]
port 334 nsew signal output
rlabel metal2 s 469466 -960 469578 480 8 la_data_out[25]
port 335 nsew signal output
rlabel metal3 s 583520 467788 584960 468028 6 la_data_out[26]
port 336 nsew signal output
rlabel metal3 s -960 92428 480 92668 4 la_data_out[27]
port 337 nsew signal output
rlabel metal2 s 309110 -960 309222 480 8 la_data_out[28]
port 338 nsew signal output
rlabel metal2 s 305246 -960 305358 480 8 la_data_out[29]
port 339 nsew signal output
rlabel metal2 s 477194 -960 477306 480 8 la_data_out[2]
port 340 nsew signal output
rlabel metal2 s 272402 703520 272514 704960 6 la_data_out[30]
port 341 nsew signal output
rlabel metal3 s -960 237948 480 238188 4 la_data_out[31]
port 342 nsew signal output
rlabel metal3 s -960 217548 480 217788 4 la_data_out[32]
port 343 nsew signal output
rlabel metal3 s 583520 201908 584960 202148 6 la_data_out[33]
port 344 nsew signal output
rlabel metal2 s 316838 -960 316950 480 8 la_data_out[34]
port 345 nsew signal output
rlabel metal3 s -960 322268 480 322508 4 la_data_out[35]
port 346 nsew signal output
rlabel metal2 s 528070 703520 528182 704960 6 la_data_out[36]
port 347 nsew signal output
rlabel metal3 s 583520 8108 584960 8348 6 la_data_out[37]
port 348 nsew signal output
rlabel metal3 s 583520 68628 584960 68868 6 la_data_out[38]
port 349 nsew signal output
rlabel metal3 s 583520 129148 584960 129388 6 la_data_out[39]
port 350 nsew signal output
rlabel metal3 s -960 80188 480 80428 4 la_data_out[3]
port 351 nsew signal output
rlabel metal3 s 583520 346748 584960 346988 6 la_data_out[40]
port 352 nsew signal output
rlabel metal2 s 371578 703520 371690 704960 6 la_data_out[41]
port 353 nsew signal output
rlabel metal2 s 245354 703520 245466 704960 6 la_data_out[42]
port 354 nsew signal output
rlabel metal3 s -960 693548 480 693788 4 la_data_out[43]
port 355 nsew signal output
rlabel metal2 s 465602 -960 465714 480 8 la_data_out[44]
port 356 nsew signal output
rlabel metal2 s 378018 -960 378130 480 8 la_data_out[45]
port 357 nsew signal output
rlabel metal2 s 84998 703520 85110 704960 6 la_data_out[46]
port 358 nsew signal output
rlabel metal3 s -960 628948 480 629188 4 la_data_out[47]
port 359 nsew signal output
rlabel metal2 s 561558 -960 561670 480 8 la_data_out[48]
port 360 nsew signal output
rlabel metal2 s 146178 703520 146290 704960 6 la_data_out[49]
port 361 nsew signal output
rlabel metal2 s 486210 703520 486322 704960 6 la_data_out[4]
port 362 nsew signal output
rlabel metal3 s -960 431068 480 431308 4 la_data_out[50]
port 363 nsew signal output
rlabel metal2 s 370290 -960 370402 480 8 la_data_out[51]
port 364 nsew signal output
rlabel metal3 s -960 84268 480 84508 4 la_data_out[52]
port 365 nsew signal output
rlabel metal2 s 440486 703520 440598 704960 6 la_data_out[53]
port 366 nsew signal output
rlabel metal2 s 397338 -960 397450 480 8 la_data_out[54]
port 367 nsew signal output
rlabel metal3 s -960 201228 480 201468 4 la_data_out[55]
port 368 nsew signal output
rlabel metal2 s 280130 703520 280242 704960 6 la_data_out[56]
port 369 nsew signal output
rlabel metal2 s 47002 703520 47114 704960 6 la_data_out[57]
port 370 nsew signal output
rlabel metal3 s 583520 125068 584960 125308 6 la_data_out[58]
port 371 nsew signal output
rlabel metal3 s 583520 427668 584960 427908 6 la_data_out[59]
port 372 nsew signal output
rlabel metal2 s 354834 -960 354946 480 8 la_data_out[5]
port 373 nsew signal output
rlabel metal3 s -960 645268 480 645508 4 la_data_out[60]
port 374 nsew signal output
rlabel metal3 s -960 411348 480 411588 4 la_data_out[61]
port 375 nsew signal output
rlabel metal2 s 362562 -960 362674 480 8 la_data_out[62]
port 376 nsew signal output
rlabel metal2 s 436622 703520 436734 704960 6 la_data_out[63]
port 377 nsew signal output
rlabel metal3 s -960 273988 480 274228 4 la_data_out[64]
port 378 nsew signal output
rlabel metal2 s 522918 -960 523030 480 8 la_data_out[65]
port 379 nsew signal output
rlabel metal3 s 583520 -52 584960 188 6 la_data_out[66]
port 380 nsew signal output
rlabel metal3 s -960 148868 480 149108 4 la_data_out[67]
port 381 nsew signal output
rlabel metal3 s -960 63868 480 64108 4 la_data_out[68]
port 382 nsew signal output
rlabel metal3 s 583520 181508 584960 181748 6 la_data_out[69]
port 383 nsew signal output
rlabel metal2 s 320702 -960 320814 480 8 la_data_out[6]
port 384 nsew signal output
rlabel metal2 s 473330 -960 473442 480 8 la_data_out[70]
port 385 nsew signal output
rlabel metal3 s -960 48228 480 48468 4 la_data_out[71]
port 386 nsew signal output
rlabel metal2 s 444350 703520 444462 704960 6 la_data_out[72]
port 387 nsew signal output
rlabel metal2 s 358698 -960 358810 480 8 la_data_out[73]
port 388 nsew signal output
rlabel metal2 s 5142 703520 5254 704960 6 la_data_out[74]
port 389 nsew signal output
rlabel metal2 s 400558 -960 400670 480 8 la_data_out[75]
port 390 nsew signal output
rlabel metal3 s -960 669068 480 669308 4 la_data_out[76]
port 391 nsew signal output
rlabel metal3 s 583520 475948 584960 476188 6 la_data_out[77]
port 392 nsew signal output
rlabel metal2 s 332294 -960 332406 480 8 la_data_out[78]
port 393 nsew signal output
rlabel metal3 s 583520 153628 584960 153868 6 la_data_out[79]
port 394 nsew signal output
rlabel metal3 s 583520 44148 584960 44388 6 la_data_out[7]
port 395 nsew signal output
rlabel metal3 s 583520 233868 584960 234108 6 la_data_out[80]
port 396 nsew signal output
rlabel metal3 s -960 572508 480 572748 4 la_data_out[81]
port 397 nsew signal output
rlabel metal2 s 247930 -960 248042 480 8 la_data_out[82]
port 398 nsew signal output
rlabel metal3 s -960 560268 480 560508 4 la_data_out[83]
port 399 nsew signal output
rlabel metal2 s 461738 -960 461850 480 8 la_data_out[84]
port 400 nsew signal output
rlabel metal2 s 517122 703520 517234 704960 6 la_data_out[85]
port 401 nsew signal output
rlabel metal2 s 115910 703520 116022 704960 6 la_data_out[86]
port 402 nsew signal output
rlabel metal2 s 578302 703520 578414 704960 6 la_data_out[87]
port 403 nsew signal output
rlabel metal3 s -960 112828 480 113068 4 la_data_out[88]
port 404 nsew signal output
rlabel metal3 s 583520 76788 584960 77028 6 la_data_out[89]
port 405 nsew signal output
rlabel metal3 s 583520 439908 584960 440148 6 la_data_out[8]
port 406 nsew signal output
rlabel metal2 s 226678 703520 226790 704960 6 la_data_out[90]
port 407 nsew signal output
rlabel metal2 s 423742 -960 423854 480 8 la_data_out[91]
port 408 nsew signal output
rlabel metal2 s 171294 -960 171406 480 8 la_data_out[92]
port 409 nsew signal output
rlabel metal2 s 417302 703520 417414 704960 6 la_data_out[93]
port 410 nsew signal output
rlabel metal2 s 496514 -960 496626 480 8 la_data_out[94]
port 411 nsew signal output
rlabel metal3 s -960 278068 480 278308 4 la_data_out[95]
port 412 nsew signal output
rlabel metal2 s 9006 703520 9118 704960 6 la_data_out[96]
port 413 nsew signal output
rlabel metal2 s 190614 -960 190726 480 8 la_data_out[97]
port 414 nsew signal output
rlabel metal2 s 555118 703520 555230 704960 6 la_data_out[98]
port 415 nsew signal output
rlabel metal2 s 511326 -960 511438 480 8 la_data_out[99]
port 416 nsew signal output
rlabel metal3 s 583520 286228 584960 286468 6 la_data_out[9]
port 417 nsew signal output
rlabel metal2 s 425030 703520 425142 704960 6 la_oenb[0]
port 418 nsew signal input
rlabel metal3 s -960 209388 480 209628 4 la_oenb[100]
port 419 nsew signal input
rlabel metal3 s -960 480028 480 480268 4 la_oenb[101]
port 420 nsew signal input
rlabel metal2 s 297518 -960 297630 480 8 la_oenb[102]
port 421 nsew signal input
rlabel metal2 s 350970 -960 351082 480 8 la_oenb[103]
port 422 nsew signal input
rlabel metal2 s 43138 703520 43250 704960 6 la_oenb[104]
port 423 nsew signal input
rlabel metal3 s 583520 161788 584960 162028 6 la_oenb[105]
port 424 nsew signal input
rlabel metal2 s 421166 703520 421278 704960 6 la_oenb[106]
port 425 nsew signal input
rlabel metal2 s 168074 -960 168186 480 8 la_oenb[107]
port 426 nsew signal input
rlabel metal3 s 583520 471868 584960 472108 6 la_oenb[108]
port 427 nsew signal input
rlabel metal2 s 177090 703520 177202 704960 6 la_oenb[109]
port 428 nsew signal input
rlabel metal2 s 513258 703520 513370 704960 6 la_oenb[10]
port 429 nsew signal input
rlabel metal2 s 142314 703520 142426 704960 6 la_oenb[110]
port 430 nsew signal input
rlabel metal2 s 35410 703520 35522 704960 6 la_oenb[111]
port 431 nsew signal input
rlabel metal3 s -960 120308 480 120548 4 la_oenb[112]
port 432 nsew signal input
rlabel metal2 s 263386 -960 263498 480 8 la_oenb[113]
port 433 nsew signal input
rlabel metal3 s 583520 596988 584960 597228 6 la_oenb[114]
port 434 nsew signal input
rlabel metal2 s 481058 -960 481170 480 8 la_oenb[115]
port 435 nsew signal input
rlabel metal3 s 583520 435828 584960 436068 6 la_oenb[116]
port 436 nsew signal input
rlabel metal2 s 125570 -960 125682 480 8 la_oenb[117]
port 437 nsew signal input
rlabel metal2 s 260810 703520 260922 704960 6 la_oenb[118]
port 438 nsew signal input
rlabel metal3 s -960 44148 480 44388 4 la_oenb[119]
port 439 nsew signal input
rlabel metal2 s 340022 -960 340134 480 8 la_oenb[11]
port 440 nsew signal input
rlabel metal2 s 562846 703520 562958 704960 6 la_oenb[120]
port 441 nsew signal input
rlabel metal3 s -960 378708 480 378948 4 la_oenb[121]
port 442 nsew signal input
rlabel metal3 s 583520 112828 584960 113068 6 la_oenb[122]
port 443 nsew signal input
rlabel metal2 s 12870 703520 12982 704960 6 la_oenb[123]
port 444 nsew signal input
rlabel metal2 s 50866 703520 50978 704960 6 la_oenb[124]
port 445 nsew signal input
rlabel metal2 s 236338 -960 236450 480 8 la_oenb[125]
port 446 nsew signal input
rlabel metal2 s 287858 703520 287970 704960 6 la_oenb[126]
port 447 nsew signal input
rlabel metal3 s 583520 637788 584960 638028 6 la_oenb[127]
port 448 nsew signal input
rlabel metal3 s 583520 302548 584960 302788 6 la_oenb[12]
port 449 nsew signal input
rlabel metal3 s -960 318188 480 318428 4 la_oenb[13]
port 450 nsew signal input
rlabel metal3 s -960 193068 480 193308 4 la_oenb[14]
port 451 nsew signal input
rlabel metal3 s 583520 246108 584960 246348 6 la_oenb[15]
port 452 nsew signal input
rlabel metal3 s -960 40068 480 40308 4 la_oenb[16]
port 453 nsew signal input
rlabel metal2 s 283994 703520 284106 704960 6 la_oenb[17]
port 454 nsew signal input
rlabel metal3 s -960 152948 480 153188 4 la_oenb[18]
port 455 nsew signal input
rlabel metal3 s -960 72028 480 72268 4 la_oenb[19]
port 456 nsew signal input
rlabel metal2 s 186750 -960 186862 480 8 la_oenb[1]
port 457 nsew signal input
rlabel metal3 s 583520 193748 584960 193988 6 la_oenb[20]
port 458 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 la_oenb[21]
port 459 nsew signal input
rlabel metal2 s 194478 -960 194590 480 8 la_oenb[22]
port 460 nsew signal input
rlabel metal3 s 583520 177428 584960 177668 6 la_oenb[23]
port 461 nsew signal input
rlabel metal2 s 582166 703520 582278 704960 6 la_oenb[24]
port 462 nsew signal input
rlabel metal3 s 583520 358988 584960 359228 6 la_oenb[25]
port 463 nsew signal input
rlabel metal2 s 68254 -960 68366 480 8 la_oenb[26]
port 464 nsew signal input
rlabel metal3 s 583520 306628 584960 306868 6 la_oenb[27]
port 465 nsew signal input
rlabel metal3 s -960 15588 480 15828 4 la_oenb[28]
port 466 nsew signal input
rlabel metal2 s 459806 703520 459918 704960 6 la_oenb[29]
port 467 nsew signal input
rlabel metal2 s 419878 -960 419990 480 8 la_oenb[2]
port 468 nsew signal input
rlabel metal3 s 583520 443988 584960 444228 6 la_oenb[30]
port 469 nsew signal input
rlabel metal2 s 539662 703520 539774 704960 6 la_oenb[31]
port 470 nsew signal input
rlabel metal3 s -960 23748 480 23988 4 la_oenb[32]
port 471 nsew signal input
rlabel metal2 s 306534 703520 306646 704960 6 la_oenb[33]
port 472 nsew signal input
rlabel metal2 s 547390 703520 547502 704960 6 la_oenb[34]
port 473 nsew signal input
rlabel metal2 s 77270 703520 77382 704960 6 la_oenb[35]
port 474 nsew signal input
rlabel metal3 s -960 301868 480 302108 4 la_oenb[36]
port 475 nsew signal input
rlabel metal3 s 583520 116908 584960 117148 6 la_oenb[37]
port 476 nsew signal input
rlabel metal3 s -960 290308 480 290548 4 la_oenb[38]
port 477 nsew signal input
rlabel metal3 s 583520 463708 584960 463948 6 la_oenb[39]
port 478 nsew signal input
rlabel metal2 s 215086 703520 215198 704960 6 la_oenb[3]
port 479 nsew signal input
rlabel metal2 s 500378 -960 500490 480 8 la_oenb[40]
port 480 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 la_oenb[41]
port 481 nsew signal input
rlabel metal3 s 583520 532388 584960 532628 6 la_oenb[42]
port 482 nsew signal input
rlabel metal2 s 490074 703520 490186 704960 6 la_oenb[43]
port 483 nsew signal input
rlabel metal3 s 583520 681988 584960 682228 6 la_oenb[44]
port 484 nsew signal input
rlabel metal3 s 583520 16268 584960 16508 6 la_oenb[45]
port 485 nsew signal input
rlabel metal3 s -960 11508 480 11748 4 la_oenb[46]
port 486 nsew signal input
rlabel metal2 s 576370 -960 576482 480 8 la_oenb[47]
port 487 nsew signal input
rlabel metal3 s 583520 108748 584960 108988 6 la_oenb[48]
port 488 nsew signal input
rlabel metal2 s 117842 -960 117954 480 8 la_oenb[49]
port 489 nsew signal input
rlabel metal2 s 175158 -960 175270 480 8 la_oenb[4]
port 490 nsew signal input
rlabel metal3 s 583520 36668 584960 36908 6 la_oenb[50]
port 491 nsew signal input
rlabel metal3 s 583520 274668 584960 274908 6 la_oenb[51]
port 492 nsew signal input
rlabel metal3 s 583520 621468 584960 621708 6 la_oenb[52]
port 493 nsew signal input
rlabel metal2 s 234406 703520 234518 704960 6 la_oenb[53]
port 494 nsew signal input
rlabel metal2 s 203494 703520 203606 704960 6 la_oenb[54]
port 495 nsew signal input
rlabel metal2 s 104318 703520 104430 704960 6 la_oenb[55]
port 496 nsew signal input
rlabel metal2 s 217662 -960 217774 480 8 la_oenb[56]
port 497 nsew signal input
rlabel metal3 s 583520 690148 584960 690388 6 la_oenb[57]
port 498 nsew signal input
rlabel metal3 s -960 180828 480 181068 4 la_oenb[58]
port 499 nsew signal input
rlabel metal2 s 66322 703520 66434 704960 6 la_oenb[59]
port 500 nsew signal input
rlabel metal3 s -960 52308 480 52548 4 la_oenb[5]
port 501 nsew signal input
rlabel metal3 s 583520 609228 584960 609468 6 la_oenb[60]
port 502 nsew signal input
rlabel metal2 s 356122 703520 356234 704960 6 la_oenb[61]
port 503 nsew signal input
rlabel metal2 s 314262 703520 314374 704960 6 la_oenb[62]
port 504 nsew signal input
rlabel metal2 s 428894 703520 429006 704960 6 la_oenb[63]
port 505 nsew signal input
rlabel metal2 s 463670 703520 463782 704960 6 la_oenb[64]
port 506 nsew signal input
rlabel metal2 s 467534 703520 467646 704960 6 la_oenb[65]
port 507 nsew signal input
rlabel metal3 s -960 241348 480 241588 4 la_oenb[66]
port 508 nsew signal input
rlabel metal2 s 249218 703520 249330 704960 6 la_oenb[67]
port 509 nsew signal input
rlabel metal3 s -960 225708 480 225948 4 la_oenb[68]
port 510 nsew signal input
rlabel metal2 s 7074 -960 7186 480 8 la_oenb[69]
port 511 nsew signal input
rlabel metal2 s 572506 -960 572618 480 8 la_oenb[6]
port 512 nsew signal input
rlabel metal3 s -960 253588 480 253828 4 la_oenb[70]
port 513 nsew signal input
rlabel metal3 s 583520 197828 584960 198068 6 la_oenb[71]
port 514 nsew signal input
rlabel metal3 s -960 443308 480 443548 4 la_oenb[72]
port 515 nsew signal input
rlabel metal3 s 583520 262428 584960 262668 6 la_oenb[73]
port 516 nsew signal input
rlabel metal3 s -960 584748 480 584988 4 la_oenb[74]
port 517 nsew signal input
rlabel metal2 s 30258 -960 30370 480 8 la_oenb[75]
port 518 nsew signal input
rlabel metal3 s -960 261748 480 261988 4 la_oenb[76]
port 519 nsew signal input
rlabel metal3 s -960 173348 480 173588 4 la_oenb[77]
port 520 nsew signal input
rlabel metal2 s 242134 703520 242246 704960 6 la_oenb[78]
port 521 nsew signal input
rlabel metal3 s 583520 4028 584960 4268 6 la_oenb[79]
port 522 nsew signal input
rlabel metal2 s 278842 -960 278954 480 8 la_oenb[7]
port 523 nsew signal input
rlabel metal3 s -960 495668 480 495908 4 la_oenb[80]
port 524 nsew signal input
rlabel metal3 s 583520 528308 584960 528548 6 la_oenb[81]
port 525 nsew signal input
rlabel metal3 s 583520 669748 584960 669988 6 la_oenb[82]
port 526 nsew signal input
rlabel metal2 s 565422 -960 565534 480 8 la_oenb[83]
port 527 nsew signal input
rlabel metal3 s -960 588828 480 589068 4 la_oenb[84]
port 528 nsew signal input
rlabel metal3 s 583520 141388 584960 141628 6 la_oenb[85]
port 529 nsew signal input
rlabel metal3 s 583520 633708 584960 633948 6 la_oenb[86]
port 530 nsew signal input
rlabel metal2 s 153906 703520 154018 704960 6 la_oenb[87]
port 531 nsew signal input
rlabel metal3 s 583520 540548 584960 540788 6 la_oenb[88]
port 532 nsew signal input
rlabel metal2 s 549966 -960 550078 480 8 la_oenb[89]
port 533 nsew signal input
rlabel metal2 s 310398 703520 310510 704960 6 la_oenb[8]
port 534 nsew signal input
rlabel metal3 s 583520 218228 584960 218468 6 la_oenb[90]
port 535 nsew signal input
rlabel metal2 s 108182 703520 108294 704960 6 la_oenb[91]
port 536 nsew signal input
rlabel metal3 s 583520 84948 584960 85188 6 la_oenb[92]
port 537 nsew signal input
rlabel metal3 s -960 422908 480 423148 4 la_oenb[93]
port 538 nsew signal input
rlabel metal2 s 91438 -960 91550 480 8 la_oenb[94]
port 539 nsew signal input
rlabel metal3 s 583520 516748 584960 516988 6 la_oenb[95]
port 540 nsew signal input
rlabel metal2 s 404422 -960 404534 480 8 la_oenb[96]
port 541 nsew signal input
rlabel metal3 s -960 221628 480 221868 4 la_oenb[97]
port 542 nsew signal input
rlabel metal2 s 182886 -960 182998 480 8 la_oenb[98]
port 543 nsew signal input
rlabel metal3 s -960 294388 480 294628 4 la_oenb[99]
port 544 nsew signal input
rlabel metal3 s -960 616708 480 616948 4 la_oenb[9]
port 545 nsew signal input
rlabel metal2 s 318126 703520 318238 704960 6 user_clock2
port 546 nsew signal input
rlabel metal3 s 583520 702388 584960 702628 6 user_irq[0]
port 547 nsew signal output
rlabel metal3 s -960 596988 480 597228 4 user_irq[1]
port 548 nsew signal output
rlabel metal3 s -960 660908 480 661148 4 user_irq[2]
port 549 nsew signal output
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 550 nsew power bidirectional
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 550 nsew power bidirectional
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 550 nsew power bidirectional
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 550 nsew power bidirectional
rlabel metal4 s 1794 -7654 2414 711590 6 vccd1
port 550 nsew power bidirectional
rlabel metal4 s 37794 -7654 38414 711590 6 vccd1
port 550 nsew power bidirectional
rlabel metal4 s 73794 -7654 74414 711590 6 vccd1
port 550 nsew power bidirectional
rlabel metal4 s 109794 -7654 110414 711590 6 vccd1
port 550 nsew power bidirectional
rlabel metal4 s 145794 -7654 146414 78000 6 vccd1
port 550 nsew power bidirectional
rlabel metal4 s 145794 142000 146414 198000 6 vccd1
port 550 nsew power bidirectional
rlabel metal4 s 145794 262000 146414 711590 6 vccd1
port 550 nsew power bidirectional
rlabel metal4 s 181794 -7654 182414 78000 6 vccd1
port 550 nsew power bidirectional
rlabel metal4 s 181794 142000 182414 198000 6 vccd1
port 550 nsew power bidirectional
rlabel metal4 s 181794 262000 182414 711590 6 vccd1
port 550 nsew power bidirectional
rlabel metal4 s 217794 -7654 218414 711590 6 vccd1
port 550 nsew power bidirectional
rlabel metal4 s 253794 -7654 254414 711590 6 vccd1
port 550 nsew power bidirectional
rlabel metal4 s 289794 -7654 290414 711590 6 vccd1
port 550 nsew power bidirectional
rlabel metal4 s 325794 -7654 326414 711590 6 vccd1
port 550 nsew power bidirectional
rlabel metal4 s 361794 -7654 362414 711590 6 vccd1
port 550 nsew power bidirectional
rlabel metal4 s 397794 -7654 398414 711590 6 vccd1
port 550 nsew power bidirectional
rlabel metal4 s 433794 -7654 434414 711590 6 vccd1
port 550 nsew power bidirectional
rlabel metal4 s 469794 -7654 470414 711590 6 vccd1
port 550 nsew power bidirectional
rlabel metal4 s 505794 -7654 506414 711590 6 vccd1
port 550 nsew power bidirectional
rlabel metal4 s 541794 -7654 542414 711590 6 vccd1
port 550 nsew power bidirectional
rlabel metal4 s 577794 -7654 578414 711590 6 vccd1
port 550 nsew power bidirectional
rlabel metal5 s -8726 2866 592650 3486 6 vccd1
port 550 nsew power bidirectional
rlabel metal5 s -8726 38866 592650 39486 6 vccd1
port 550 nsew power bidirectional
rlabel metal5 s -8726 74866 592650 75486 6 vccd1
port 550 nsew power bidirectional
rlabel metal5 s -8726 110866 592650 111486 6 vccd1
port 550 nsew power bidirectional
rlabel metal5 s -8726 146866 592650 147486 6 vccd1
port 550 nsew power bidirectional
rlabel metal5 s -8726 182866 592650 183486 6 vccd1
port 550 nsew power bidirectional
rlabel metal5 s -8726 218866 592650 219486 6 vccd1
port 550 nsew power bidirectional
rlabel metal5 s -8726 254866 592650 255486 6 vccd1
port 550 nsew power bidirectional
rlabel metal5 s -8726 290866 592650 291486 6 vccd1
port 550 nsew power bidirectional
rlabel metal5 s -8726 326866 592650 327486 6 vccd1
port 550 nsew power bidirectional
rlabel metal5 s -8726 362866 592650 363486 6 vccd1
port 550 nsew power bidirectional
rlabel metal5 s -8726 398866 592650 399486 6 vccd1
port 550 nsew power bidirectional
rlabel metal5 s -8726 434866 592650 435486 6 vccd1
port 550 nsew power bidirectional
rlabel metal5 s -8726 470866 592650 471486 6 vccd1
port 550 nsew power bidirectional
rlabel metal5 s -8726 506866 592650 507486 6 vccd1
port 550 nsew power bidirectional
rlabel metal5 s -8726 542866 592650 543486 6 vccd1
port 550 nsew power bidirectional
rlabel metal5 s -8726 578866 592650 579486 6 vccd1
port 550 nsew power bidirectional
rlabel metal5 s -8726 614866 592650 615486 6 vccd1
port 550 nsew power bidirectional
rlabel metal5 s -8726 650866 592650 651486 6 vccd1
port 550 nsew power bidirectional
rlabel metal5 s -8726 686866 592650 687486 6 vccd1
port 550 nsew power bidirectional
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 551 nsew power bidirectional
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 551 nsew power bidirectional
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 551 nsew power bidirectional
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 551 nsew power bidirectional
rlabel metal4 s 10794 -7654 11414 711590 6 vccd2
port 551 nsew power bidirectional
rlabel metal4 s 46794 -7654 47414 711590 6 vccd2
port 551 nsew power bidirectional
rlabel metal4 s 82794 -7654 83414 711590 6 vccd2
port 551 nsew power bidirectional
rlabel metal4 s 118794 -7654 119414 78000 6 vccd2
port 551 nsew power bidirectional
rlabel metal4 s 118794 142000 119414 198000 6 vccd2
port 551 nsew power bidirectional
rlabel metal4 s 118794 262000 119414 711590 6 vccd2
port 551 nsew power bidirectional
rlabel metal4 s 154794 -7654 155414 78000 6 vccd2
port 551 nsew power bidirectional
rlabel metal4 s 154794 142000 155414 198000 6 vccd2
port 551 nsew power bidirectional
rlabel metal4 s 154794 262000 155414 711590 6 vccd2
port 551 nsew power bidirectional
rlabel metal4 s 190794 -7654 191414 78000 6 vccd2
port 551 nsew power bidirectional
rlabel metal4 s 190794 142000 191414 198000 6 vccd2
port 551 nsew power bidirectional
rlabel metal4 s 190794 262000 191414 711590 6 vccd2
port 551 nsew power bidirectional
rlabel metal4 s 226794 -7654 227414 711590 6 vccd2
port 551 nsew power bidirectional
rlabel metal4 s 262794 -7654 263414 711590 6 vccd2
port 551 nsew power bidirectional
rlabel metal4 s 298794 -7654 299414 711590 6 vccd2
port 551 nsew power bidirectional
rlabel metal4 s 334794 -7654 335414 711590 6 vccd2
port 551 nsew power bidirectional
rlabel metal4 s 370794 -7654 371414 711590 6 vccd2
port 551 nsew power bidirectional
rlabel metal4 s 406794 -7654 407414 711590 6 vccd2
port 551 nsew power bidirectional
rlabel metal4 s 442794 -7654 443414 711590 6 vccd2
port 551 nsew power bidirectional
rlabel metal4 s 478794 -7654 479414 711590 6 vccd2
port 551 nsew power bidirectional
rlabel metal4 s 514794 -7654 515414 711590 6 vccd2
port 551 nsew power bidirectional
rlabel metal4 s 550794 -7654 551414 711590 6 vccd2
port 551 nsew power bidirectional
rlabel metal5 s -8726 11866 592650 12486 6 vccd2
port 551 nsew power bidirectional
rlabel metal5 s -8726 47866 592650 48486 6 vccd2
port 551 nsew power bidirectional
rlabel metal5 s -8726 83866 592650 84486 6 vccd2
port 551 nsew power bidirectional
rlabel metal5 s -8726 119866 592650 120486 6 vccd2
port 551 nsew power bidirectional
rlabel metal5 s -8726 155866 592650 156486 6 vccd2
port 551 nsew power bidirectional
rlabel metal5 s -8726 191866 592650 192486 6 vccd2
port 551 nsew power bidirectional
rlabel metal5 s -8726 227866 592650 228486 6 vccd2
port 551 nsew power bidirectional
rlabel metal5 s -8726 263866 592650 264486 6 vccd2
port 551 nsew power bidirectional
rlabel metal5 s -8726 299866 592650 300486 6 vccd2
port 551 nsew power bidirectional
rlabel metal5 s -8726 335866 592650 336486 6 vccd2
port 551 nsew power bidirectional
rlabel metal5 s -8726 371866 592650 372486 6 vccd2
port 551 nsew power bidirectional
rlabel metal5 s -8726 407866 592650 408486 6 vccd2
port 551 nsew power bidirectional
rlabel metal5 s -8726 443866 592650 444486 6 vccd2
port 551 nsew power bidirectional
rlabel metal5 s -8726 479866 592650 480486 6 vccd2
port 551 nsew power bidirectional
rlabel metal5 s -8726 515866 592650 516486 6 vccd2
port 551 nsew power bidirectional
rlabel metal5 s -8726 551866 592650 552486 6 vccd2
port 551 nsew power bidirectional
rlabel metal5 s -8726 587866 592650 588486 6 vccd2
port 551 nsew power bidirectional
rlabel metal5 s -8726 623866 592650 624486 6 vccd2
port 551 nsew power bidirectional
rlabel metal5 s -8726 659866 592650 660486 6 vccd2
port 551 nsew power bidirectional
rlabel metal5 s -8726 695866 592650 696486 6 vccd2
port 551 nsew power bidirectional
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 552 nsew power bidirectional
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 552 nsew power bidirectional
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 552 nsew power bidirectional
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 552 nsew power bidirectional
rlabel metal4 s 19794 -7654 20414 711590 6 vdda1
port 552 nsew power bidirectional
rlabel metal4 s 55794 -7654 56414 711590 6 vdda1
port 552 nsew power bidirectional
rlabel metal4 s 91794 -7654 92414 711590 6 vdda1
port 552 nsew power bidirectional
rlabel metal4 s 127794 -7654 128414 78000 6 vdda1
port 552 nsew power bidirectional
rlabel metal4 s 127794 262000 128414 711590 6 vdda1
port 552 nsew power bidirectional
rlabel metal4 s 163794 -7654 164414 78000 6 vdda1
port 552 nsew power bidirectional
rlabel metal4 s 163794 262000 164414 711590 6 vdda1
port 552 nsew power bidirectional
rlabel metal4 s 199794 -7654 200414 711590 6 vdda1
port 552 nsew power bidirectional
rlabel metal4 s 235794 -7654 236414 711590 6 vdda1
port 552 nsew power bidirectional
rlabel metal4 s 271794 -7654 272414 711590 6 vdda1
port 552 nsew power bidirectional
rlabel metal4 s 307794 -7654 308414 711590 6 vdda1
port 552 nsew power bidirectional
rlabel metal4 s 343794 -7654 344414 711590 6 vdda1
port 552 nsew power bidirectional
rlabel metal4 s 379794 -7654 380414 711590 6 vdda1
port 552 nsew power bidirectional
rlabel metal4 s 415794 -7654 416414 711590 6 vdda1
port 552 nsew power bidirectional
rlabel metal4 s 451794 -7654 452414 711590 6 vdda1
port 552 nsew power bidirectional
rlabel metal4 s 487794 -7654 488414 711590 6 vdda1
port 552 nsew power bidirectional
rlabel metal4 s 523794 -7654 524414 711590 6 vdda1
port 552 nsew power bidirectional
rlabel metal4 s 559794 -7654 560414 711590 6 vdda1
port 552 nsew power bidirectional
rlabel metal5 s -8726 20866 592650 21486 6 vdda1
port 552 nsew power bidirectional
rlabel metal5 s -8726 56866 592650 57486 6 vdda1
port 552 nsew power bidirectional
rlabel metal5 s -8726 92866 592650 93486 6 vdda1
port 552 nsew power bidirectional
rlabel metal5 s -8726 128866 592650 129486 6 vdda1
port 552 nsew power bidirectional
rlabel metal5 s -8726 164866 592650 165486 6 vdda1
port 552 nsew power bidirectional
rlabel metal5 s -8726 200866 592650 201486 6 vdda1
port 552 nsew power bidirectional
rlabel metal5 s -8726 236866 592650 237486 6 vdda1
port 552 nsew power bidirectional
rlabel metal5 s -8726 272866 592650 273486 6 vdda1
port 552 nsew power bidirectional
rlabel metal5 s -8726 308866 592650 309486 6 vdda1
port 552 nsew power bidirectional
rlabel metal5 s -8726 344866 592650 345486 6 vdda1
port 552 nsew power bidirectional
rlabel metal5 s -8726 380866 592650 381486 6 vdda1
port 552 nsew power bidirectional
rlabel metal5 s -8726 416866 592650 417486 6 vdda1
port 552 nsew power bidirectional
rlabel metal5 s -8726 452866 592650 453486 6 vdda1
port 552 nsew power bidirectional
rlabel metal5 s -8726 488866 592650 489486 6 vdda1
port 552 nsew power bidirectional
rlabel metal5 s -8726 524866 592650 525486 6 vdda1
port 552 nsew power bidirectional
rlabel metal5 s -8726 560866 592650 561486 6 vdda1
port 552 nsew power bidirectional
rlabel metal5 s -8726 596866 592650 597486 6 vdda1
port 552 nsew power bidirectional
rlabel metal5 s -8726 632866 592650 633486 6 vdda1
port 552 nsew power bidirectional
rlabel metal5 s -8726 668866 592650 669486 6 vdda1
port 552 nsew power bidirectional
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 553 nsew power bidirectional
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 553 nsew power bidirectional
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 553 nsew power bidirectional
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 553 nsew power bidirectional
rlabel metal4 s 28794 -7654 29414 711590 6 vdda2
port 553 nsew power bidirectional
rlabel metal4 s 64794 -7654 65414 711590 6 vdda2
port 553 nsew power bidirectional
rlabel metal4 s 100794 -7654 101414 711590 6 vdda2
port 553 nsew power bidirectional
rlabel metal4 s 136794 -7654 137414 78000 6 vdda2
port 553 nsew power bidirectional
rlabel metal4 s 136794 262000 137414 711590 6 vdda2
port 553 nsew power bidirectional
rlabel metal4 s 172794 -7654 173414 78000 6 vdda2
port 553 nsew power bidirectional
rlabel metal4 s 172794 262000 173414 711590 6 vdda2
port 553 nsew power bidirectional
rlabel metal4 s 208794 -7654 209414 711590 6 vdda2
port 553 nsew power bidirectional
rlabel metal4 s 244794 -7654 245414 711590 6 vdda2
port 553 nsew power bidirectional
rlabel metal4 s 280794 -7654 281414 711590 6 vdda2
port 553 nsew power bidirectional
rlabel metal4 s 316794 -7654 317414 711590 6 vdda2
port 553 nsew power bidirectional
rlabel metal4 s 352794 -7654 353414 711590 6 vdda2
port 553 nsew power bidirectional
rlabel metal4 s 388794 -7654 389414 711590 6 vdda2
port 553 nsew power bidirectional
rlabel metal4 s 424794 -7654 425414 711590 6 vdda2
port 553 nsew power bidirectional
rlabel metal4 s 460794 -7654 461414 711590 6 vdda2
port 553 nsew power bidirectional
rlabel metal4 s 496794 -7654 497414 711590 6 vdda2
port 553 nsew power bidirectional
rlabel metal4 s 532794 -7654 533414 711590 6 vdda2
port 553 nsew power bidirectional
rlabel metal4 s 568794 -7654 569414 711590 6 vdda2
port 553 nsew power bidirectional
rlabel metal5 s -8726 29866 592650 30486 6 vdda2
port 553 nsew power bidirectional
rlabel metal5 s -8726 65866 592650 66486 6 vdda2
port 553 nsew power bidirectional
rlabel metal5 s -8726 101866 592650 102486 6 vdda2
port 553 nsew power bidirectional
rlabel metal5 s -8726 137866 592650 138486 6 vdda2
port 553 nsew power bidirectional
rlabel metal5 s -8726 173866 592650 174486 6 vdda2
port 553 nsew power bidirectional
rlabel metal5 s -8726 209866 592650 210486 6 vdda2
port 553 nsew power bidirectional
rlabel metal5 s -8726 245866 592650 246486 6 vdda2
port 553 nsew power bidirectional
rlabel metal5 s -8726 281866 592650 282486 6 vdda2
port 553 nsew power bidirectional
rlabel metal5 s -8726 317866 592650 318486 6 vdda2
port 553 nsew power bidirectional
rlabel metal5 s -8726 353866 592650 354486 6 vdda2
port 553 nsew power bidirectional
rlabel metal5 s -8726 389866 592650 390486 6 vdda2
port 553 nsew power bidirectional
rlabel metal5 s -8726 425866 592650 426486 6 vdda2
port 553 nsew power bidirectional
rlabel metal5 s -8726 461866 592650 462486 6 vdda2
port 553 nsew power bidirectional
rlabel metal5 s -8726 497866 592650 498486 6 vdda2
port 553 nsew power bidirectional
rlabel metal5 s -8726 533866 592650 534486 6 vdda2
port 553 nsew power bidirectional
rlabel metal5 s -8726 569866 592650 570486 6 vdda2
port 553 nsew power bidirectional
rlabel metal5 s -8726 605866 592650 606486 6 vdda2
port 553 nsew power bidirectional
rlabel metal5 s -8726 641866 592650 642486 6 vdda2
port 553 nsew power bidirectional
rlabel metal5 s -8726 677866 592650 678486 6 vdda2
port 553 nsew power bidirectional
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 554 nsew ground bidirectional
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 554 nsew ground bidirectional
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 554 nsew ground bidirectional
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 554 nsew ground bidirectional
rlabel metal4 s 24294 -7654 24914 711590 6 vssa1
port 554 nsew ground bidirectional
rlabel metal4 s 60294 -7654 60914 711590 6 vssa1
port 554 nsew ground bidirectional
rlabel metal4 s 96294 -7654 96914 711590 6 vssa1
port 554 nsew ground bidirectional
rlabel metal4 s 132294 -7654 132914 78000 6 vssa1
port 554 nsew ground bidirectional
rlabel metal4 s 132294 262000 132914 711590 6 vssa1
port 554 nsew ground bidirectional
rlabel metal4 s 168294 -7654 168914 78000 6 vssa1
port 554 nsew ground bidirectional
rlabel metal4 s 168294 262000 168914 711590 6 vssa1
port 554 nsew ground bidirectional
rlabel metal4 s 204294 -7654 204914 711590 6 vssa1
port 554 nsew ground bidirectional
rlabel metal4 s 240294 -7654 240914 711590 6 vssa1
port 554 nsew ground bidirectional
rlabel metal4 s 276294 -7654 276914 711590 6 vssa1
port 554 nsew ground bidirectional
rlabel metal4 s 312294 -7654 312914 711590 6 vssa1
port 554 nsew ground bidirectional
rlabel metal4 s 348294 -7654 348914 711590 6 vssa1
port 554 nsew ground bidirectional
rlabel metal4 s 384294 -7654 384914 711590 6 vssa1
port 554 nsew ground bidirectional
rlabel metal4 s 420294 -7654 420914 711590 6 vssa1
port 554 nsew ground bidirectional
rlabel metal4 s 456294 -7654 456914 711590 6 vssa1
port 554 nsew ground bidirectional
rlabel metal4 s 492294 -7654 492914 711590 6 vssa1
port 554 nsew ground bidirectional
rlabel metal4 s 528294 -7654 528914 711590 6 vssa1
port 554 nsew ground bidirectional
rlabel metal4 s 564294 -7654 564914 711590 6 vssa1
port 554 nsew ground bidirectional
rlabel metal5 s -8726 25366 592650 25986 6 vssa1
port 554 nsew ground bidirectional
rlabel metal5 s -8726 61366 592650 61986 6 vssa1
port 554 nsew ground bidirectional
rlabel metal5 s -8726 97366 592650 97986 6 vssa1
port 554 nsew ground bidirectional
rlabel metal5 s -8726 133366 592650 133986 6 vssa1
port 554 nsew ground bidirectional
rlabel metal5 s -8726 169366 592650 169986 6 vssa1
port 554 nsew ground bidirectional
rlabel metal5 s -8726 205366 592650 205986 6 vssa1
port 554 nsew ground bidirectional
rlabel metal5 s -8726 241366 592650 241986 6 vssa1
port 554 nsew ground bidirectional
rlabel metal5 s -8726 277366 592650 277986 6 vssa1
port 554 nsew ground bidirectional
rlabel metal5 s -8726 313366 592650 313986 6 vssa1
port 554 nsew ground bidirectional
rlabel metal5 s -8726 349366 592650 349986 6 vssa1
port 554 nsew ground bidirectional
rlabel metal5 s -8726 385366 592650 385986 6 vssa1
port 554 nsew ground bidirectional
rlabel metal5 s -8726 421366 592650 421986 6 vssa1
port 554 nsew ground bidirectional
rlabel metal5 s -8726 457366 592650 457986 6 vssa1
port 554 nsew ground bidirectional
rlabel metal5 s -8726 493366 592650 493986 6 vssa1
port 554 nsew ground bidirectional
rlabel metal5 s -8726 529366 592650 529986 6 vssa1
port 554 nsew ground bidirectional
rlabel metal5 s -8726 565366 592650 565986 6 vssa1
port 554 nsew ground bidirectional
rlabel metal5 s -8726 601366 592650 601986 6 vssa1
port 554 nsew ground bidirectional
rlabel metal5 s -8726 637366 592650 637986 6 vssa1
port 554 nsew ground bidirectional
rlabel metal5 s -8726 673366 592650 673986 6 vssa1
port 554 nsew ground bidirectional
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 555 nsew ground bidirectional
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 555 nsew ground bidirectional
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 555 nsew ground bidirectional
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 555 nsew ground bidirectional
rlabel metal4 s 33294 -7654 33914 711590 6 vssa2
port 555 nsew ground bidirectional
rlabel metal4 s 69294 -7654 69914 711590 6 vssa2
port 555 nsew ground bidirectional
rlabel metal4 s 105294 -7654 105914 711590 6 vssa2
port 555 nsew ground bidirectional
rlabel metal4 s 141294 -7654 141914 78000 6 vssa2
port 555 nsew ground bidirectional
rlabel metal4 s 141294 142000 141914 198000 6 vssa2
port 555 nsew ground bidirectional
rlabel metal4 s 141294 262000 141914 711590 6 vssa2
port 555 nsew ground bidirectional
rlabel metal4 s 177294 -7654 177914 78000 6 vssa2
port 555 nsew ground bidirectional
rlabel metal4 s 177294 142000 177914 198000 6 vssa2
port 555 nsew ground bidirectional
rlabel metal4 s 177294 262000 177914 711590 6 vssa2
port 555 nsew ground bidirectional
rlabel metal4 s 213294 -7654 213914 711590 6 vssa2
port 555 nsew ground bidirectional
rlabel metal4 s 249294 -7654 249914 711590 6 vssa2
port 555 nsew ground bidirectional
rlabel metal4 s 285294 -7654 285914 711590 6 vssa2
port 555 nsew ground bidirectional
rlabel metal4 s 321294 -7654 321914 711590 6 vssa2
port 555 nsew ground bidirectional
rlabel metal4 s 357294 -7654 357914 711590 6 vssa2
port 555 nsew ground bidirectional
rlabel metal4 s 393294 -7654 393914 711590 6 vssa2
port 555 nsew ground bidirectional
rlabel metal4 s 429294 -7654 429914 711590 6 vssa2
port 555 nsew ground bidirectional
rlabel metal4 s 465294 -7654 465914 711590 6 vssa2
port 555 nsew ground bidirectional
rlabel metal4 s 501294 -7654 501914 711590 6 vssa2
port 555 nsew ground bidirectional
rlabel metal4 s 537294 -7654 537914 711590 6 vssa2
port 555 nsew ground bidirectional
rlabel metal4 s 573294 -7654 573914 711590 6 vssa2
port 555 nsew ground bidirectional
rlabel metal5 s -8726 34366 592650 34986 6 vssa2
port 555 nsew ground bidirectional
rlabel metal5 s -8726 70366 592650 70986 6 vssa2
port 555 nsew ground bidirectional
rlabel metal5 s -8726 106366 592650 106986 6 vssa2
port 555 nsew ground bidirectional
rlabel metal5 s -8726 142366 592650 142986 6 vssa2
port 555 nsew ground bidirectional
rlabel metal5 s -8726 178366 592650 178986 6 vssa2
port 555 nsew ground bidirectional
rlabel metal5 s -8726 214366 592650 214986 6 vssa2
port 555 nsew ground bidirectional
rlabel metal5 s -8726 250366 592650 250986 6 vssa2
port 555 nsew ground bidirectional
rlabel metal5 s -8726 286366 592650 286986 6 vssa2
port 555 nsew ground bidirectional
rlabel metal5 s -8726 322366 592650 322986 6 vssa2
port 555 nsew ground bidirectional
rlabel metal5 s -8726 358366 592650 358986 6 vssa2
port 555 nsew ground bidirectional
rlabel metal5 s -8726 394366 592650 394986 6 vssa2
port 555 nsew ground bidirectional
rlabel metal5 s -8726 430366 592650 430986 6 vssa2
port 555 nsew ground bidirectional
rlabel metal5 s -8726 466366 592650 466986 6 vssa2
port 555 nsew ground bidirectional
rlabel metal5 s -8726 502366 592650 502986 6 vssa2
port 555 nsew ground bidirectional
rlabel metal5 s -8726 538366 592650 538986 6 vssa2
port 555 nsew ground bidirectional
rlabel metal5 s -8726 574366 592650 574986 6 vssa2
port 555 nsew ground bidirectional
rlabel metal5 s -8726 610366 592650 610986 6 vssa2
port 555 nsew ground bidirectional
rlabel metal5 s -8726 646366 592650 646986 6 vssa2
port 555 nsew ground bidirectional
rlabel metal5 s -8726 682366 592650 682986 6 vssa2
port 555 nsew ground bidirectional
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 556 nsew ground bidirectional
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 556 nsew ground bidirectional
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 556 nsew ground bidirectional
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 556 nsew ground bidirectional
rlabel metal4 s 6294 -7654 6914 711590 6 vssd1
port 556 nsew ground bidirectional
rlabel metal4 s 42294 -7654 42914 711590 6 vssd1
port 556 nsew ground bidirectional
rlabel metal4 s 78294 -7654 78914 711590 6 vssd1
port 556 nsew ground bidirectional
rlabel metal4 s 114294 -7654 114914 711590 6 vssd1
port 556 nsew ground bidirectional
rlabel metal4 s 150294 -7654 150914 78000 6 vssd1
port 556 nsew ground bidirectional
rlabel metal4 s 150294 142000 150914 198000 6 vssd1
port 556 nsew ground bidirectional
rlabel metal4 s 150294 262000 150914 711590 6 vssd1
port 556 nsew ground bidirectional
rlabel metal4 s 186294 -7654 186914 78000 6 vssd1
port 556 nsew ground bidirectional
rlabel metal4 s 186294 142000 186914 198000 6 vssd1
port 556 nsew ground bidirectional
rlabel metal4 s 186294 262000 186914 711590 6 vssd1
port 556 nsew ground bidirectional
rlabel metal4 s 222294 -7654 222914 711590 6 vssd1
port 556 nsew ground bidirectional
rlabel metal4 s 258294 -7654 258914 711590 6 vssd1
port 556 nsew ground bidirectional
rlabel metal4 s 294294 -7654 294914 711590 6 vssd1
port 556 nsew ground bidirectional
rlabel metal4 s 330294 -7654 330914 711590 6 vssd1
port 556 nsew ground bidirectional
rlabel metal4 s 366294 -7654 366914 711590 6 vssd1
port 556 nsew ground bidirectional
rlabel metal4 s 402294 -7654 402914 711590 6 vssd1
port 556 nsew ground bidirectional
rlabel metal4 s 438294 -7654 438914 711590 6 vssd1
port 556 nsew ground bidirectional
rlabel metal4 s 474294 -7654 474914 711590 6 vssd1
port 556 nsew ground bidirectional
rlabel metal4 s 510294 -7654 510914 711590 6 vssd1
port 556 nsew ground bidirectional
rlabel metal4 s 546294 -7654 546914 711590 6 vssd1
port 556 nsew ground bidirectional
rlabel metal4 s 582294 -7654 582914 711590 6 vssd1
port 556 nsew ground bidirectional
rlabel metal5 s -8726 7366 592650 7986 6 vssd1
port 556 nsew ground bidirectional
rlabel metal5 s -8726 43366 592650 43986 6 vssd1
port 556 nsew ground bidirectional
rlabel metal5 s -8726 79366 592650 79986 6 vssd1
port 556 nsew ground bidirectional
rlabel metal5 s -8726 115366 592650 115986 6 vssd1
port 556 nsew ground bidirectional
rlabel metal5 s -8726 151366 592650 151986 6 vssd1
port 556 nsew ground bidirectional
rlabel metal5 s -8726 187366 592650 187986 6 vssd1
port 556 nsew ground bidirectional
rlabel metal5 s -8726 223366 592650 223986 6 vssd1
port 556 nsew ground bidirectional
rlabel metal5 s -8726 259366 592650 259986 6 vssd1
port 556 nsew ground bidirectional
rlabel metal5 s -8726 295366 592650 295986 6 vssd1
port 556 nsew ground bidirectional
rlabel metal5 s -8726 331366 592650 331986 6 vssd1
port 556 nsew ground bidirectional
rlabel metal5 s -8726 367366 592650 367986 6 vssd1
port 556 nsew ground bidirectional
rlabel metal5 s -8726 403366 592650 403986 6 vssd1
port 556 nsew ground bidirectional
rlabel metal5 s -8726 439366 592650 439986 6 vssd1
port 556 nsew ground bidirectional
rlabel metal5 s -8726 475366 592650 475986 6 vssd1
port 556 nsew ground bidirectional
rlabel metal5 s -8726 511366 592650 511986 6 vssd1
port 556 nsew ground bidirectional
rlabel metal5 s -8726 547366 592650 547986 6 vssd1
port 556 nsew ground bidirectional
rlabel metal5 s -8726 583366 592650 583986 6 vssd1
port 556 nsew ground bidirectional
rlabel metal5 s -8726 619366 592650 619986 6 vssd1
port 556 nsew ground bidirectional
rlabel metal5 s -8726 655366 592650 655986 6 vssd1
port 556 nsew ground bidirectional
rlabel metal5 s -8726 691366 592650 691986 6 vssd1
port 556 nsew ground bidirectional
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 557 nsew ground bidirectional
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 557 nsew ground bidirectional
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 557 nsew ground bidirectional
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 557 nsew ground bidirectional
rlabel metal4 s 15294 -7654 15914 711590 6 vssd2
port 557 nsew ground bidirectional
rlabel metal4 s 51294 -7654 51914 711590 6 vssd2
port 557 nsew ground bidirectional
rlabel metal4 s 87294 -7654 87914 711590 6 vssd2
port 557 nsew ground bidirectional
rlabel metal4 s 123294 -7654 123914 78000 6 vssd2
port 557 nsew ground bidirectional
rlabel metal4 s 123294 142000 123914 198000 6 vssd2
port 557 nsew ground bidirectional
rlabel metal4 s 123294 262000 123914 711590 6 vssd2
port 557 nsew ground bidirectional
rlabel metal4 s 159294 -7654 159914 78000 6 vssd2
port 557 nsew ground bidirectional
rlabel metal4 s 159294 142000 159914 198000 6 vssd2
port 557 nsew ground bidirectional
rlabel metal4 s 159294 262000 159914 711590 6 vssd2
port 557 nsew ground bidirectional
rlabel metal4 s 195294 -7654 195914 711590 6 vssd2
port 557 nsew ground bidirectional
rlabel metal4 s 231294 -7654 231914 711590 6 vssd2
port 557 nsew ground bidirectional
rlabel metal4 s 267294 -7654 267914 711590 6 vssd2
port 557 nsew ground bidirectional
rlabel metal4 s 303294 -7654 303914 711590 6 vssd2
port 557 nsew ground bidirectional
rlabel metal4 s 339294 -7654 339914 711590 6 vssd2
port 557 nsew ground bidirectional
rlabel metal4 s 375294 -7654 375914 711590 6 vssd2
port 557 nsew ground bidirectional
rlabel metal4 s 411294 -7654 411914 711590 6 vssd2
port 557 nsew ground bidirectional
rlabel metal4 s 447294 -7654 447914 711590 6 vssd2
port 557 nsew ground bidirectional
rlabel metal4 s 483294 -7654 483914 711590 6 vssd2
port 557 nsew ground bidirectional
rlabel metal4 s 519294 -7654 519914 711590 6 vssd2
port 557 nsew ground bidirectional
rlabel metal4 s 555294 -7654 555914 711590 6 vssd2
port 557 nsew ground bidirectional
rlabel metal5 s -8726 16366 592650 16986 6 vssd2
port 557 nsew ground bidirectional
rlabel metal5 s -8726 52366 592650 52986 6 vssd2
port 557 nsew ground bidirectional
rlabel metal5 s -8726 88366 592650 88986 6 vssd2
port 557 nsew ground bidirectional
rlabel metal5 s -8726 124366 592650 124986 6 vssd2
port 557 nsew ground bidirectional
rlabel metal5 s -8726 160366 592650 160986 6 vssd2
port 557 nsew ground bidirectional
rlabel metal5 s -8726 196366 592650 196986 6 vssd2
port 557 nsew ground bidirectional
rlabel metal5 s -8726 232366 592650 232986 6 vssd2
port 557 nsew ground bidirectional
rlabel metal5 s -8726 268366 592650 268986 6 vssd2
port 557 nsew ground bidirectional
rlabel metal5 s -8726 304366 592650 304986 6 vssd2
port 557 nsew ground bidirectional
rlabel metal5 s -8726 340366 592650 340986 6 vssd2
port 557 nsew ground bidirectional
rlabel metal5 s -8726 376366 592650 376986 6 vssd2
port 557 nsew ground bidirectional
rlabel metal5 s -8726 412366 592650 412986 6 vssd2
port 557 nsew ground bidirectional
rlabel metal5 s -8726 448366 592650 448986 6 vssd2
port 557 nsew ground bidirectional
rlabel metal5 s -8726 484366 592650 484986 6 vssd2
port 557 nsew ground bidirectional
rlabel metal5 s -8726 520366 592650 520986 6 vssd2
port 557 nsew ground bidirectional
rlabel metal5 s -8726 556366 592650 556986 6 vssd2
port 557 nsew ground bidirectional
rlabel metal5 s -8726 592366 592650 592986 6 vssd2
port 557 nsew ground bidirectional
rlabel metal5 s -8726 628366 592650 628986 6 vssd2
port 557 nsew ground bidirectional
rlabel metal5 s -8726 664366 592650 664986 6 vssd2
port 557 nsew ground bidirectional
rlabel metal5 s -8726 700366 592650 700986 6 vssd2
port 557 nsew ground bidirectional
rlabel metal3 s 583520 258348 584960 258588 6 wb_clk_i
port 558 nsew signal input
rlabel metal3 s -960 350828 480 351068 4 wb_rst_i
port 559 nsew signal input
rlabel metal3 s 583520 383468 584960 383708 6 wbs_ack_o
port 560 nsew signal output
rlabel metal2 s 199630 703520 199742 704960 6 wbs_adr_i[0]
port 561 nsew signal input
rlabel metal2 s 54730 703520 54842 704960 6 wbs_adr_i[10]
port 562 nsew signal input
rlabel metal3 s -960 471868 480 472108 4 wbs_adr_i[11]
port 563 nsew signal input
rlabel metal2 s 64390 -960 64502 480 8 wbs_adr_i[12]
port 564 nsew signal input
rlabel metal2 s 389610 -960 389722 480 8 wbs_adr_i[13]
port 565 nsew signal input
rlabel metal3 s 583520 657508 584960 657748 6 wbs_adr_i[14]
port 566 nsew signal input
rlabel metal3 s 583520 613308 584960 613548 6 wbs_adr_i[15]
port 567 nsew signal input
rlabel metal2 s 443062 -960 443174 480 8 wbs_adr_i[16]
port 568 nsew signal input
rlabel metal3 s 583520 556868 584960 557108 6 wbs_adr_i[17]
port 569 nsew signal input
rlabel metal3 s 583520 343348 584960 343588 6 wbs_adr_i[18]
port 570 nsew signal input
rlabel metal3 s 583520 89028 584960 89268 6 wbs_adr_i[19]
port 571 nsew signal input
rlabel metal2 s 207358 703520 207470 704960 6 wbs_adr_i[1]
port 572 nsew signal input
rlabel metal2 s 406354 703520 406466 704960 6 wbs_adr_i[20]
port 573 nsew signal input
rlabel metal2 s 393474 -960 393586 480 8 wbs_adr_i[21]
port 574 nsew signal input
rlabel metal2 s 557694 -960 557806 480 8 wbs_adr_i[22]
port 575 nsew signal input
rlabel metal3 s 583520 278748 584960 278988 6 wbs_adr_i[23]
port 576 nsew signal input
rlabel metal3 s -960 556188 480 556428 4 wbs_adr_i[24]
port 577 nsew signal input
rlabel metal2 s 374154 -960 374266 480 8 wbs_adr_i[25]
port 578 nsew signal input
rlabel metal2 s 72118 -960 72230 480 8 wbs_adr_i[26]
port 579 nsew signal input
rlabel metal3 s -960 19668 480 19908 4 wbs_adr_i[27]
port 580 nsew signal input
rlabel metal3 s 583520 524228 584960 524468 6 wbs_adr_i[28]
port 581 nsew signal input
rlabel metal2 s 497802 703520 497914 704960 6 wbs_adr_i[29]
port 582 nsew signal input
rlabel metal2 s 267250 -960 267362 480 8 wbs_adr_i[2]
port 583 nsew signal input
rlabel metal2 s 333582 703520 333694 704960 6 wbs_adr_i[30]
port 584 nsew signal input
rlabel metal3 s 583520 403868 584960 404108 6 wbs_adr_i[31]
port 585 nsew signal input
rlabel metal2 s 530646 -960 530758 480 8 wbs_adr_i[3]
port 586 nsew signal input
rlabel metal2 s 321990 703520 322102 704960 6 wbs_adr_i[4]
port 587 nsew signal input
rlabel metal3 s -960 108748 480 108988 4 wbs_adr_i[5]
port 588 nsew signal input
rlabel metal2 s 213798 -960 213910 480 8 wbs_adr_i[6]
port 589 nsew signal input
rlabel metal2 s 34122 -960 34234 480 8 wbs_adr_i[7]
port 590 nsew signal input
rlabel metal3 s 583520 97188 584960 97428 6 wbs_adr_i[8]
port 591 nsew signal input
rlabel metal3 s 583520 290308 584960 290548 6 wbs_adr_i[9]
port 592 nsew signal input
rlabel metal2 s 31546 703520 31658 704960 6 wbs_cyc_i
port 593 nsew signal input
rlabel metal2 s 574438 703520 574550 704960 6 wbs_dat_i[0]
port 594 nsew signal input
rlabel metal3 s -960 358988 480 359228 4 wbs_dat_i[10]
port 595 nsew signal input
rlabel metal3 s -960 407268 480 407508 4 wbs_dat_i[11]
port 596 nsew signal input
rlabel metal3 s -960 390948 480 391188 4 wbs_dat_i[12]
port 597 nsew signal input
rlabel metal2 s 26394 -960 26506 480 8 wbs_dat_i[13]
port 598 nsew signal input
rlabel metal2 s 144890 -960 145002 480 8 wbs_dat_i[14]
port 599 nsew signal input
rlabel metal3 s 583520 456228 584960 456468 6 wbs_dat_i[15]
port 600 nsew signal input
rlabel metal2 s 385746 -960 385858 480 8 wbs_dat_i[16]
port 601 nsew signal input
rlabel metal2 s 291722 703520 291834 704960 6 wbs_dat_i[17]
port 602 nsew signal input
rlabel metal2 s 455942 703520 456054 704960 6 wbs_dat_i[18]
port 603 nsew signal input
rlabel metal3 s -960 576588 480 576828 4 wbs_dat_i[19]
port 604 nsew signal input
rlabel metal2 s 103030 -960 103142 480 8 wbs_dat_i[1]
port 605 nsew signal input
rlabel metal3 s 583520 508588 584960 508828 6 wbs_dat_i[20]
port 606 nsew signal input
rlabel metal2 s 482346 703520 482458 704960 6 wbs_dat_i[21]
port 607 nsew signal input
rlabel metal3 s -960 265828 480 266068 4 wbs_dat_i[22]
port 608 nsew signal input
rlabel metal3 s 583520 629628 584960 629868 6 wbs_dat_i[23]
port 609 nsew signal input
rlabel metal3 s 583520 310708 584960 310948 6 wbs_dat_i[24]
port 610 nsew signal input
rlabel metal2 s 457874 -960 457986 480 8 wbs_dat_i[25]
port 611 nsew signal input
rlabel metal2 s 410218 703520 410330 704960 6 wbs_dat_i[26]
port 612 nsew signal input
rlabel metal2 s 19954 703520 20066 704960 6 wbs_dat_i[27]
port 613 nsew signal input
rlabel metal2 s 206070 -960 206182 480 8 wbs_dat_i[28]
port 614 nsew signal input
rlabel metal3 s 583520 496348 584960 496588 6 wbs_dat_i[29]
port 615 nsew signal input
rlabel metal2 s 538374 -960 538486 480 8 wbs_dat_i[2]
port 616 nsew signal input
rlabel metal3 s 583520 282828 584960 283068 6 wbs_dat_i[30]
port 617 nsew signal input
rlabel metal3 s -960 249508 480 249748 4 wbs_dat_i[31]
port 618 nsew signal input
rlabel metal3 s 583520 101268 584960 101508 6 wbs_dat_i[3]
port 619 nsew signal input
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_i[4]
port 620 nsew signal input
rlabel metal2 s 324566 -960 324678 480 8 wbs_dat_i[5]
port 621 nsew signal input
rlabel metal3 s -960 3348 480 3588 4 wbs_dat_i[6]
port 622 nsew signal input
rlabel metal2 s 398626 703520 398738 704960 6 wbs_dat_i[7]
port 623 nsew signal input
rlabel metal3 s 583520 686068 584960 686308 6 wbs_dat_i[8]
port 624 nsew signal input
rlabel metal3 s 583520 104668 584960 104908 6 wbs_dat_i[9]
port 625 nsew signal input
rlabel metal2 s 53442 -960 53554 480 8 wbs_dat_o[0]
port 626 nsew signal output
rlabel metal3 s 583520 460308 584960 460548 6 wbs_dat_o[10]
port 627 nsew signal output
rlabel metal2 s 14802 -960 14914 480 8 wbs_dat_o[11]
port 628 nsew signal output
rlabel metal3 s 583520 694228 584960 694468 6 wbs_dat_o[12]
port 629 nsew signal output
rlabel metal2 s 383170 703520 383282 704960 6 wbs_dat_o[13]
port 630 nsew signal output
rlabel metal3 s 583520 145468 584960 145708 6 wbs_dat_o[14]
port 631 nsew signal output
rlabel metal2 s 363850 703520 363962 704960 6 wbs_dat_o[15]
port 632 nsew signal output
rlabel metal3 s -960 116908 480 117148 4 wbs_dat_o[16]
port 633 nsew signal output
rlabel metal3 s -960 136628 480 136868 4 wbs_dat_o[17]
port 634 nsew signal output
rlabel metal2 s 435334 -960 435446 480 8 wbs_dat_o[18]
port 635 nsew signal output
rlabel metal2 s -10 -960 102 480 8 wbs_dat_o[19]
port 636 nsew signal output
rlabel metal2 s 508106 -960 508218 480 8 wbs_dat_o[1]
port 637 nsew signal output
rlabel metal3 s -960 257668 480 257908 4 wbs_dat_o[20]
port 638 nsew signal output
rlabel metal3 s -960 524228 480 524468 4 wbs_dat_o[21]
port 639 nsew signal output
rlabel metal2 s 92726 703520 92838 704960 6 wbs_dat_o[22]
port 640 nsew signal output
rlabel metal3 s -960 169268 480 169508 4 wbs_dat_o[23]
port 641 nsew signal output
rlabel metal2 s 133298 -960 133410 480 8 wbs_dat_o[24]
port 642 nsew signal output
rlabel metal2 s 49578 -960 49690 480 8 wbs_dat_o[25]
port 643 nsew signal output
rlabel metal2 s 256946 703520 257058 704960 6 wbs_dat_o[26]
port 644 nsew signal output
rlabel metal2 s 112046 703520 112158 704960 6 wbs_dat_o[27]
port 645 nsew signal output
rlabel metal2 s 347106 -960 347218 480 8 wbs_dat_o[28]
port 646 nsew signal output
rlabel metal2 s 367714 703520 367826 704960 6 wbs_dat_o[29]
port 647 nsew signal output
rlabel metal3 s 583520 242028 584960 242268 6 wbs_dat_o[2]
port 648 nsew signal output
rlabel metal3 s -960 403188 480 403428 4 wbs_dat_o[30]
port 649 nsew signal output
rlabel metal3 s 583520 569108 584960 569348 6 wbs_dat_o[31]
port 650 nsew signal output
rlabel metal2 s 141026 -960 141138 480 8 wbs_dat_o[3]
port 651 nsew signal output
rlabel metal2 s 244066 -960 244178 480 8 wbs_dat_o[4]
port 652 nsew signal output
rlabel metal3 s -960 35988 480 36228 4 wbs_dat_o[5]
port 653 nsew signal output
rlabel metal3 s 583520 544628 584960 544868 6 wbs_dat_o[6]
port 654 nsew signal output
rlabel metal2 s 381882 -960 381994 480 8 wbs_dat_o[7]
port 655 nsew signal output
rlabel metal2 s 359986 703520 360098 704960 6 wbs_dat_o[8]
port 656 nsew signal output
rlabel metal2 s 352902 703520 353014 704960 6 wbs_dat_o[9]
port 657 nsew signal output
rlabel metal3 s -960 600388 480 600628 4 wbs_sel_i[0]
port 658 nsew signal input
rlabel metal2 s 16090 703520 16202 704960 6 wbs_sel_i[1]
port 659 nsew signal input
rlabel metal2 s 454654 -960 454766 480 8 wbs_sel_i[2]
port 660 nsew signal input
rlabel metal3 s -960 140708 480 140948 4 wbs_sel_i[3]
port 661 nsew signal input
rlabel metal3 s -960 543948 480 544188 4 wbs_stb_i
port 662 nsew signal input
rlabel metal3 s 583520 371228 584960 371468 6 wbs_we_i
port 663 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 7875646
string GDS_FILE /home/mxmont/Documents/Universidad/IC-UBB/MixPix/CARAVEL_WRAPPER/MixPix/openlane/user_project_wrapper/runs/22_10_29_10_11/results/signoff/user_analog_project_wrapper.magic.gds
string GDS_START 4284720
<< end >>

